-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Aug 18 2020 14:56:45

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    TX : out std_logic;
    GPIO11 : out std_logic;
    CLK : in std_logic;
    RX : in std_logic;
    GPIO9 : out std_logic;
    GPIO3 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49310\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46223\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVFTDI.RXbuffer_3C_net\ : std_logic;
signal \INVFTDI.RXbuffer_0C_net\ : std_logic;
signal \ctrlOut_8\ : std_logic;
signal \ALU.m289_nsZ0Z_1_cascade_\ : std_logic;
signal \ctrlOut_5\ : std_logic;
signal \ALU.N_223_0_cascade_\ : std_logic;
signal \ALU.a9_b_3_cascade_\ : std_logic;
signal \ALU.a7_b_5\ : std_logic;
signal \ALU.a9_b_3\ : std_logic;
signal \ALU.g0_0_a3_2_0_cascade_\ : std_logic;
signal \ALU.madd_315_0_cascade_\ : std_logic;
signal \ALU.a12_b_1\ : std_logic;
signal \ALU.madd_315_0\ : std_logic;
signal \ALU.a12_b_1_cascade_\ : std_logic;
signal \ALU.madd_264\ : std_logic;
signal \ALU.madd_141_0_cascade_\ : std_logic;
signal \ALU.N_1545_0\ : std_logic;
signal \ALU.madd_166_0\ : std_logic;
signal \ALU.madd_254_0_tz_cascade_\ : std_logic;
signal \ALU.madd_141\ : std_logic;
signal \ALU.madd_254_cascade_\ : std_logic;
signal \ALU.madd_254_0_tz\ : std_logic;
signal \ALU.m292_nsZ0Z_1\ : std_logic;
signal \ALU.N_90_0_cascade_\ : std_logic;
signal \ctrlOut_6\ : std_logic;
signal \ALU.N_217_0_cascade_\ : std_logic;
signal \ALU.un9_addsub_axb_10_cascade_\ : std_logic;
signal \ALU.a3_b_0_10_cascade_\ : std_logic;
signal \ALU.g0_2_cascade_\ : std_logic;
signal \ALU.N_1555_0\ : std_logic;
signal \ALU.N_1527_0\ : std_logic;
signal \ALU.madd_171_cascade_\ : std_logic;
signal \ALU.madd_161_0_cascade_\ : std_logic;
signal \ALU.madd_161\ : std_logic;
signal \ALU.madd_166\ : std_logic;
signal \ALU.madd_171\ : std_logic;
signal \ALU.madd_161_cascade_\ : std_logic;
signal \ALU.a8_b_3_cascade_\ : std_logic;
signal \ALU.a8_b_3\ : std_logic;
signal \ALU.g0_0_2\ : std_logic;
signal \ALU.g0_0_cascade_\ : std_logic;
signal \ALU.N_1527_1_0\ : std_logic;
signal \ALU.g2_0_1\ : std_logic;
signal \ALU.g1\ : std_logic;
signal \ALU.g0_1_0\ : std_logic;
signal \ALU.madd_124_0_cascade_\ : std_logic;
signal \ALU.madd_124_cascade_\ : std_logic;
signal \ALU.madd_144_cascade_\ : std_logic;
signal \ALU.madd_324_cascade_\ : std_logic;
signal \ALU.madd_N_9_cascade_\ : std_logic;
signal \ALU.madd_191_0\ : std_logic;
signal \ALU.madd_186\ : std_logic;
signal \ALU.madd_191_0_cascade_\ : std_logic;
signal \ALU.madd_324\ : std_logic;
signal \ALU.madd_326_cascade_\ : std_logic;
signal \ALU.madd_325\ : std_logic;
signal \clkdivZ0Z_0\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \clkdivZ0Z_1\ : std_logic;
signal clkdiv_cry_0 : std_logic;
signal \clkdivZ0Z_2\ : std_logic;
signal clkdiv_cry_1 : std_logic;
signal \clkdivZ0Z_3\ : std_logic;
signal clkdiv_cry_2 : std_logic;
signal \clkdivZ0Z_4\ : std_logic;
signal clkdiv_cry_3 : std_logic;
signal \clkdivZ0Z_5\ : std_logic;
signal clkdiv_cry_4 : std_logic;
signal \clkdivZ0Z_6\ : std_logic;
signal clkdiv_cry_5 : std_logic;
signal \clkdivZ0Z_7\ : std_logic;
signal clkdiv_cry_6 : std_logic;
signal clkdiv_cry_7 : std_logic;
signal \clkdivZ0Z_8\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \clkdivZ0Z_9\ : std_logic;
signal clkdiv_cry_8 : std_logic;
signal \clkdivZ0Z_10\ : std_logic;
signal clkdiv_cry_9 : std_logic;
signal \clkdivZ0Z_11\ : std_logic;
signal clkdiv_cry_10 : std_logic;
signal \clkdivZ0Z_12\ : std_logic;
signal clkdiv_cry_11 : std_logic;
signal \clkdivZ0Z_13\ : std_logic;
signal clkdiv_cry_12 : std_logic;
signal \clkdivZ0Z_14\ : std_logic;
signal clkdiv_cry_13 : std_logic;
signal \clkdivZ0Z_15\ : std_logic;
signal clkdiv_cry_14 : std_logic;
signal clkdiv_cry_15 : std_logic;
signal \clkdivZ0Z_16\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \clkdivZ0Z_17\ : std_logic;
signal clkdiv_cry_16 : std_logic;
signal \clkdivZ0Z_18\ : std_logic;
signal clkdiv_cry_17 : std_logic;
signal \clkdivZ0Z_19\ : std_logic;
signal clkdiv_cry_18 : std_logic;
signal \clkdivZ0Z_20\ : std_logic;
signal clkdiv_cry_19 : std_logic;
signal \clkdivZ0Z_21\ : std_logic;
signal clkdiv_cry_20 : std_logic;
signal \clkdivZ0Z_22\ : std_logic;
signal clkdiv_cry_21 : std_logic;
signal clkdiv_cry_22 : std_logic;
signal \GPIO3_c\ : std_logic;
signal \testWordZ0Z_13\ : std_logic;
signal \ALU.m304_nsZ0Z_1_cascade_\ : std_logic;
signal \ALU.i73_mux_1_cascade_\ : std_logic;
signal \RXbuffer_0\ : std_logic;
signal \RXbuffer_7\ : std_logic;
signal \RXbuffer_1\ : std_logic;
signal \RXbuffer_3\ : std_logic;
signal \N_661_0_cascade_\ : std_logic;
signal \ALU.un2_addsub_axb_8_cascade_\ : std_logic;
signal \ALU.N_275_0_cascade_\ : std_logic;
signal \ALU.g0_0_0_N_3L3\ : std_logic;
signal \ALU.g0_0_0_N_4L5_cascade_\ : std_logic;
signal \ALU.g0_0_0_N_3L3_0\ : std_logic;
signal \ALU.a5_b_9_cascade_\ : std_logic;
signal \ALU.operand2_8_cascade_\ : std_logic;
signal \ALU.a1_b_8\ : std_logic;
signal \ALU.a1_b_8_cascade_\ : std_logic;
signal \ALU.a4_b_8_cascade_\ : std_logic;
signal \ALU.madd_269\ : std_logic;
signal \ALU.madd_i1_mux_cascade_\ : std_logic;
signal \ALU.g0_14\ : std_logic;
signal \ALU.madd_i3_mux_cascade_\ : std_logic;
signal \ALU.madd_331_cascade_\ : std_logic;
signal \ALU.madd_328\ : std_logic;
signal \ALU.madd_340_0\ : std_logic;
signal \ALU.g0_1_cascade_\ : std_logic;
signal \ALU.g2\ : std_logic;
signal \ALU.N_1545_1\ : std_logic;
signal \ALU.g0_3_cascade_\ : std_logic;
signal \ALU.madd_350_0\ : std_logic;
signal \ALU.madd_350_0_cascade_\ : std_logic;
signal \ALU.madd_335\ : std_logic;
signal \ALU.madd_i1_mux_2\ : std_logic;
signal \ALU.madd_289\ : std_logic;
signal \ALU.madd_227\ : std_logic;
signal \ALU.madd_227_cascade_\ : std_logic;
signal \ALU.madd_165_0_0_cascade_\ : std_logic;
signal \ALU.madd_170_0_tz_cascade_\ : std_logic;
signal \ALU.madd_90\ : std_logic;
signal \ALU.madd_223_0_cascade_\ : std_logic;
signal \ALU.N_1533_0\ : std_logic;
signal \ALU.N_1559_0\ : std_logic;
signal \ALU.madd_165_0_tz\ : std_logic;
signal \ALU.madd_165_0\ : std_logic;
signal \ALU.a5_b_5\ : std_logic;
signal \ALU.a5_b_5_cascade_\ : std_logic;
signal \ALU.a4_b_6\ : std_logic;
signal \ALU.madd_175_cascade_\ : std_logic;
signal \ALU.madd_232\ : std_logic;
signal \ALU.madd_175\ : std_logic;
signal \ALU.madd_213_0\ : std_logic;
signal \ALU.a7_b_4_cascade_\ : std_logic;
signal \ALU.madd_208\ : std_logic;
signal \ALU.N_225_0_cascade_\ : std_logic;
signal \ALU.madd_290_0_cascade_\ : std_logic;
signal \ALU.madd_299_cascade_\ : std_logic;
signal \ALU.g0_11\ : std_logic;
signal \ALU.madd_299\ : std_logic;
signal \ALU.madd_223_0\ : std_logic;
signal \ALU.madd_228\ : std_logic;
signal \ALU.madd_170\ : std_logic;
signal \ALU.madd_265_0_cascade_\ : std_logic;
signal \ALU.madd_280\ : std_logic;
signal \ALU.madd_280_cascade_\ : std_logic;
signal \ALU.madd_285\ : std_logic;
signal \ALU.madd_326\ : std_logic;
signal \ALU.a4_b_7\ : std_logic;
signal \ALU.a4_b_7_cascade_\ : std_logic;
signal \ALU.madd_233_cascade_\ : std_logic;
signal \ALU.madd_237\ : std_logic;
signal \ALU.madd_242\ : std_logic;
signal \ALU.madd_247_cascade_\ : std_logic;
signal \ALU.madd_295_0\ : std_logic;
signal \ALU.madd_N_10\ : std_logic;
signal \ALU.madd_247\ : std_logic;
signal \ALU.madd_N_10_cascade_\ : std_logic;
signal \ALU.madd_N_5_0\ : std_logic;
signal \ALU.madd_190\ : std_logic;
signal \ALU.madd_238_0\ : std_logic;
signal \ALU.madd_233\ : std_logic;
signal \ALU.madd_327\ : std_logic;
signal \ALU.un2_addsub_axb_7_cascade_\ : std_logic;
signal \ALU.a0_b_8_cascade_\ : std_logic;
signal \ALU.madd_103\ : std_logic;
signal \ALU.madd_124\ : std_logic;
signal \ALU.madd_148\ : std_logic;
signal \ALU.madd_148_cascade_\ : std_logic;
signal \ALU.madd_247_0_tz_0\ : std_logic;
signal \ALU.madd_143\ : std_logic;
signal \ALU.madd_181\ : std_logic;
signal \ALU.madd_129\ : std_logic;
signal \ALU.a5_b_4\ : std_logic;
signal \ALU.a5_b_4_cascade_\ : std_logic;
signal \ALU.madd_133_cascade_\ : std_logic;
signal \ALU.madd_237_0_tz_0\ : std_logic;
signal \ALU.madd_133\ : std_logic;
signal \ALU.madd_138\ : std_logic;
signal \ALU.madd_128_0_0_0_cascade_\ : std_logic;
signal \ALU.madd_70\ : std_logic;
signal \ALU.madd_237_0_tz_0_1_cascade_\ : std_logic;
signal \ALU.g0_0_0\ : std_logic;
signal \ALU.N_1537_0_0_1\ : std_logic;
signal \ALU.i6_mux_cascade_\ : std_logic;
signal \N_51_0_cascade_\ : std_logic;
signal \testWordZ0Z_15\ : std_logic;
signal \N_662_0_cascade_\ : std_logic;
signal \N_665_0\ : std_logic;
signal \N_301_0_cascade_\ : std_logic;
signal \N_668_0_cascade_\ : std_logic;
signal \ALU.m300_nsZ0Z_1\ : std_logic;
signal \N_662_0\ : std_logic;
signal \N_670_0_cascade_\ : std_logic;
signal \CONTROL.results_cnvZ0Z_0\ : std_logic;
signal \ALU.un2_addsub_axb_14\ : std_logic;
signal \ALU.un2_addsub_axb_9_cascade_\ : std_logic;
signal \ALU.a13_b_1_cascade_\ : std_logic;
signal \ALU.a11_b_3\ : std_logic;
signal \ALU.a11_b_3_cascade_\ : std_logic;
signal \ctrlOut_14\ : std_logic;
signal \RXbuffer_6\ : std_logic;
signal \testWordZ0Z_14\ : std_logic;
signal \ALU.a7_b_6_cascade_\ : std_logic;
signal \ALU.a6_b_7\ : std_logic;
signal \ALU.a7_b_6\ : std_logic;
signal \ALU.madd_324_0\ : std_logic;
signal \ALU.madd_324_0_cascade_\ : std_logic;
signal \ALU.madd_372\ : std_logic;
signal \ALU.madd_396\ : std_logic;
signal \ALU.madd_484_21\ : std_logic;
signal \ALU.madd_411_cascade_\ : std_logic;
signal \ALU.madd_484_24\ : std_logic;
signal \ALU.a8_b_6\ : std_logic;
signal \ALU.a9_b_5\ : std_logic;
signal \ALU.madd_377\ : std_logic;
signal \ALU.madd_372_0\ : std_logic;
signal \ALU.madd_382\ : std_logic;
signal \ALU.madd_377_cascade_\ : std_logic;
signal \ALU.a13_b_1\ : std_logic;
signal \ALU.madd_397\ : std_logic;
signal \ALU.madd_392\ : std_logic;
signal \ALU.madd_397_cascade_\ : std_logic;
signal \ALU.madd_339\ : std_logic;
signal \ALU.madd_406\ : std_logic;
signal \ALU.a5_b_8_cascade_\ : std_logic;
signal \ALU.madd_387\ : std_logic;
signal \ALU.madd_329_0\ : std_logic;
signal \ALU.madd_387_cascade_\ : std_logic;
signal \ALU.madd_402\ : std_logic;
signal \ALU.madd_402_cascade_\ : std_logic;
signal \ALU.madd_354\ : std_logic;
signal \ALU.madd_412_cascade_\ : std_logic;
signal \ALU.madd_329\ : std_logic;
signal \ALU.madd_407\ : std_logic;
signal \ALU.madd_412\ : std_logic;
signal \ALU.madd_i3_mux_1\ : std_logic;
signal \ALU.madd_330\ : std_logic;
signal \ALU.madd_141_1\ : std_logic;
signal \ALU.madd_270_0\ : std_logic;
signal \ALU.madd_250_0\ : std_logic;
signal \ALU.madd_250_0_cascade_\ : std_logic;
signal \ALU.madd_250\ : std_logic;
signal \ALU.a3_b_9\ : std_logic;
signal \ALU.madd_250_cascade_\ : std_logic;
signal \ALU.madd_207\ : std_logic;
signal \ALU.madd_274\ : std_logic;
signal \ALU.madd_320\ : std_logic;
signal \ALU.madd_325_0\ : std_logic;
signal \ALU.madd_274_cascade_\ : std_logic;
signal \ALU.madd_254\ : std_logic;
signal \ALU.madd_344\ : std_logic;
signal \ALU.madd_29_cascade_\ : std_logic;
signal \ALU.madd_47_cascade_\ : std_logic;
signal \ALU.madd_265_0\ : std_logic;
signal \ALU.madd_260\ : std_logic;
signal \ALU.a2_b_6\ : std_logic;
signal \ALU.a0_b_8\ : std_logic;
signal \ALU.a2_b_6_cascade_\ : std_logic;
signal \ALU.a5_b_6_cascade_\ : std_logic;
signal \ALU.operand2_5_cascade_\ : std_logic;
signal \ALU.madd_176_0\ : std_logic;
signal \ALU.madd_218_0\ : std_logic;
signal \ALU.a7_b_4\ : std_logic;
signal \ALU.a6_b_5\ : std_logic;
signal \ALU.a5_b_6\ : std_logic;
signal \ALU.madd_275_0\ : std_logic;
signal \ALU.madd_42_cascade_\ : std_logic;
signal \ALU.madd_42_0\ : std_logic;
signal \ALU.e_RNIM09HZ0Z_7_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_7_cascade_\ : std_logic;
signal \ALU.g1_2_cascade_\ : std_logic;
signal \ALU.a4_b_0_7\ : std_logic;
signal \ALU.g2_0_0_0\ : std_logic;
signal \ALU.un2_addsub_axb_5_cascade_\ : std_logic;
signal \ALU.a6_b_0_7\ : std_logic;
signal \ALU.a6_b_0_cascade_\ : std_logic;
signal \ALU.madd_41_cascade_\ : std_logic;
signal \ALU.madd_46_cascade_\ : std_logic;
signal \ALU.madd_39_cascade_\ : std_logic;
signal \ALU.a6_b_3\ : std_logic;
signal \ALU.madd_78_0_tz_cascade_\ : std_logic;
signal \ALU.madd_78_0\ : std_logic;
signal \ALU.madd_39\ : std_logic;
signal \ALU.madd_78_0_cascade_\ : std_logic;
signal \ALU.madd_114_cascade_\ : std_logic;
signal \testClock_0_cascade_\ : std_logic;
signal \ALU.a_cnv_0Z0Z_0_cascade_\ : std_logic;
signal \ALU.N_53_0\ : std_logic;
signal \aluResults_0\ : std_logic;
signal \testClock_0\ : std_logic;
signal \testClockZ0\ : std_logic;
signal \ALU.a_cnv_0Z0Z_0\ : std_logic;
signal \aluResults_1\ : std_logic;
signal \ALU.b_cnv_0Z0Z_0\ : std_logic;
signal \aluResults_2\ : std_logic;
signal \ALU.N_169_0\ : std_logic;
signal \ALU.c_RNIEP354Z0Z_14_cascade_\ : std_logic;
signal \ALU.c_RNIJENJ8_0Z0Z_15\ : std_logic;
signal \ALU.rshift_3_ns_1_6_cascade_\ : std_logic;
signal \ALU.N_474_cascade_\ : std_logic;
signal \ALU.rshift_15_ns_1_6\ : std_logic;
signal \ALU.rshift_6_cascade_\ : std_logic;
signal \ALU.N_291_0\ : std_logic;
signal \ALU.dout_6_ns_1_14_cascade_\ : std_logic;
signal \ALU.aluOut_15_cascade_\ : std_logic;
signal \ALU.N_761\ : std_logic;
signal \ALU.N_713\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_14_cascade_\ : std_logic;
signal \ALU.lshift_15_ns_1_14_cascade_\ : std_logic;
signal \ALU.lshift_14_cascade_\ : std_logic;
signal \ALU.a_15_m2_14\ : std_logic;
signal \ALU.a_15_m4_14_cascade_\ : std_logic;
signal \ALU.a_15_m3_14\ : std_logic;
signal \ALU.dout_3_ns_1_12_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_12_cascade_\ : std_logic;
signal \ALU.N_711\ : std_logic;
signal \ALU.N_759_cascade_\ : std_logic;
signal \ALU.aluOut_12_cascade_\ : std_logic;
signal \ALU.a12_b_2\ : std_logic;
signal \ALU.N_90_0\ : std_logic;
signal \ctrlOut_3\ : std_logic;
signal \ALU.N_235_0_cascade_\ : std_logic;
signal \ALU.a12_b_3_cascade_\ : std_logic;
signal \ctrlOut_4\ : std_logic;
signal \ALU.a9_b_4\ : std_logic;
signal \ALU.a10_b_3_cascade_\ : std_logic;
signal \ALU.madd_319\ : std_logic;
signal \ALU.madd_366\ : std_logic;
signal \ALU.madd_484_11\ : std_logic;
signal \ALU.madd_376\ : std_logic;
signal \ALU.madd_484_17_cascade_\ : std_logic;
signal \ALU.madd_484_15\ : std_logic;
signal \ALU.madd_484_20\ : std_logic;
signal \ALU.madd_309\ : std_logic;
signal \ALU.madd_362\ : std_logic;
signal \ALU.madd_391\ : std_logic;
signal \ALU.a5_b_9\ : std_logic;
signal \ALU.a6_b_8\ : std_logic;
signal \ALU.a7_b_7_cascade_\ : std_logic;
signal \ALU.madd_381\ : std_logic;
signal \ALU.madd_484_16\ : std_logic;
signal \ALU.un9_addsub_axb_12_cascade_\ : std_logic;
signal \ALU.d_RNIV96U8Z0Z_13_cascade_\ : std_logic;
signal \ALU.madd_314\ : std_logic;
signal \ALU.madd_310_0_cascade_\ : std_logic;
signal \ALU.madd_334\ : std_logic;
signal \ALU.a1_b_12\ : std_logic;
signal \ALU.a2_b_9_cascade_\ : std_logic;
signal \ALU.operand2_8\ : std_logic;
signal \ALU.N_199_0\ : std_logic;
signal \ALU.a3_b_8\ : std_logic;
signal \ALU.madd_275\ : std_logic;
signal \ALU.madd_217\ : std_logic;
signal \ALU.madd_222\ : std_logic;
signal \ALU.madd_212\ : std_logic;
signal \ALU.madd_284\ : std_logic;
signal \ALU.madd_279_cascade_\ : std_logic;
signal \ALU.madd_349\ : std_logic;
signal \ALU.d_RNIV96U8Z0Z_13\ : std_logic;
signal \ALU.madd_310_0\ : std_logic;
signal \ALU.madd_330_0\ : std_logic;
signal \ALU.c_RNIF549Z0Z_10_cascade_\ : std_logic;
signal \ALU.a_RNIBLBOZ0Z_10\ : std_logic;
signal \ALU.operand2_7_ns_1_10_cascade_\ : std_logic;
signal \ALU.operand2_10_cascade_\ : std_logic;
signal \ALU.a4_b_10\ : std_logic;
signal \ALU.a3_b_10\ : std_logic;
signal \ALU.a3_b_10_cascade_\ : std_logic;
signal \ALU.madd_305\ : std_logic;
signal \ALU.madd_5_cascade_\ : std_logic;
signal \ALU.madd_19\ : std_logic;
signal \ALU.madd_17\ : std_logic;
signal \ALU.madd_19_cascade_\ : std_logic;
signal \ALU.madd_47\ : std_logic;
signal \ALU.g0_0_a3_0\ : std_logic;
signal \ALU.a8_b_0_cascade_\ : std_logic;
signal \ALU.madd_10_cascade_\ : std_logic;
signal \ALU.madd_24\ : std_logic;
signal \ALU.madd_29\ : std_logic;
signal \ALU.madd_24_cascade_\ : std_logic;
signal \ALU.madd_i1_mux_1\ : std_logic;
signal \ALU.madd_i3_mux_0\ : std_logic;
signal \ALU.a4_b_2\ : std_logic;
signal \ALU.a6_b_0\ : std_logic;
signal \ALU.madd_12_cascade_\ : std_logic;
signal \ALU.madd_34\ : std_logic;
signal \ALU.madd_42\ : std_logic;
signal \ALU.madd_34_cascade_\ : std_logic;
signal \ALU.madd_37\ : std_logic;
signal \ALU.madd_56_cascade_\ : std_logic;
signal \ALU.madd_52_0\ : std_logic;
signal \ALU.madd_25\ : std_logic;
signal \ALU.madd_12\ : std_logic;
signal \ALU.un2_addsub_axb_6_cascade_\ : std_logic;
signal \ALU.madd_64_0\ : std_logic;
signal \ALU.madd_74_0_cascade_\ : std_logic;
signal \ALU.madd_83\ : std_logic;
signal \ALU.madd_46\ : std_logic;
signal \ALU.madd_69\ : std_logic;
signal \ALU.madd_74_0\ : std_logic;
signal \ALU.madd_79_0\ : std_logic;
signal \ALU.madd_51\ : std_logic;
signal \ALU.madd_58\ : std_logic;
signal \ALU.madd_79_0_cascade_\ : std_logic;
signal \ALU.madd_56\ : std_logic;
signal \ALU.madd_88_cascade_\ : std_logic;
signal \ALU.madd_114\ : std_logic;
signal \ALU.madd_41\ : std_logic;
signal \ALU.madd_73_cascade_\ : std_logic;
signal \ALU.operand2_7\ : std_logic;
signal \ALU.a0_b_7\ : std_logic;
signal \ALU.madd_144\ : std_logic;
signal \ALU.madd_113\ : std_logic;
signal \ALU.madd_154_cascade_\ : std_logic;
signal \ALU.madd_99\ : std_logic;
signal \ALU.madd_73\ : std_logic;
signal \ALU.madd_109\ : std_logic;
signal \ALU.madd_154\ : std_logic;
signal \ALU.madd_118\ : std_logic;
signal \ALU.m641_nsZ0Z_1\ : std_logic;
signal \ALU.m645_nsZ0Z_1\ : std_logic;
signal \ALU.N_283_0_cascade_\ : std_logic;
signal \ALU.m55_bmZ0\ : std_logic;
signal \ALU.m55_amZ0\ : std_logic;
signal \ALU.m650_nsZ0Z_1_cascade_\ : std_logic;
signal \ALU.N_15_0\ : std_logic;
signal \N_727\ : std_logic;
signal \ALU.N_577_cascade_\ : std_logic;
signal \ALU.N_528_cascade_\ : std_logic;
signal \ALU.N_633\ : std_logic;
signal \ALU.d_RNI8DL9U1Z0Z_3_cascade_\ : std_logic;
signal \ALU.N_221_cascade_\ : std_logic;
signal \ALU.N_588_cascade_\ : std_logic;
signal \ALU.N_575\ : std_logic;
signal \ALU.N_575_cascade_\ : std_logic;
signal \ALU.rshift_3_ns_1_8\ : std_logic;
signal \ALU.lshift_3_ns_1_15\ : std_logic;
signal \ALU.dout_3_ns_1_14\ : std_logic;
signal \ALU.lshift_3_ns_1_14_cascade_\ : std_logic;
signal \ALU.N_256\ : std_logic;
signal \ALU.N_224_cascade_\ : std_logic;
signal \ALU.N_220_cascade_\ : std_logic;
signal \ALU.N_222\ : std_logic;
signal \ALU.madd_484_4\ : std_logic;
signal \ALU.N_241_0\ : std_logic;
signal \ALU.N_240_0_i_cascade_\ : std_logic;
signal \ALU.N_9_0\ : std_logic;
signal \ALU.N_10_0\ : std_logic;
signal \ALU.N_253_0\ : std_logic;
signal \ALU.d_RNIUV3H4Z0Z_0\ : std_logic;
signal \ALU.N_635_0\ : std_logic;
signal \ALU.N_724\ : std_logic;
signal \ALU.N_283_0\ : std_logic;
signal \ctrlOut_7\ : std_logic;
signal \ALU.N_211_0\ : std_logic;
signal \ctrlOut_9\ : std_logic;
signal \ALU.madd_367\ : std_logic;
signal \ALU.d_RNIRV558Z0Z_13\ : std_logic;
signal \ALU.d_RNIRV558Z0Z_13_cascade_\ : std_logic;
signal \ALU.madd_371\ : std_logic;
signal \ALU.a2_b_12\ : std_logic;
signal \ALU.madd_259\ : std_logic;
signal \ALU.N_186_0_cascade_\ : std_logic;
signal \ALU.a1_b_11\ : std_logic;
signal \ALU.a0_b_12\ : std_logic;
signal \ALU.a1_b_11_cascade_\ : std_logic;
signal \ALU.madd_255\ : std_logic;
signal \ALU.dout_6_ns_1_8_cascade_\ : std_logic;
signal \ALU.dout_3_ns_1_8\ : std_logic;
signal \ALU.N_707_cascade_\ : std_logic;
signal \ALU.N_755\ : std_logic;
signal \ALU.m272_nsZ0Z_1_cascade_\ : std_logic;
signal \ALU.N_191_0_0\ : std_logic;
signal \ctrlOut_10\ : std_logic;
signal \ALU.N_191_0\ : std_logic;
signal \ALU.N_191_0_cascade_\ : std_logic;
signal \ALU.operand2_10\ : std_logic;
signal \ALU.a1_b_10\ : std_logic;
signal \ALU.a1_b_10_cascade_\ : std_logic;
signal \ALU.madd_203\ : std_logic;
signal \ALU.a9_b_2\ : std_logic;
signal \ALU.dout_3_ns_1_9_cascade_\ : std_logic;
signal \ALU.N_708_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_9_cascade_\ : std_logic;
signal \ALU.N_756\ : std_logic;
signal \ALU.N_751_cascade_\ : std_logic;
signal \ALU.N_703\ : std_logic;
signal \ALU.rshift_3_ns_1_4_cascade_\ : std_logic;
signal \ALU.N_472\ : std_logic;
signal \ALU.N_472_cascade_\ : std_logic;
signal \ALU.N_476\ : std_logic;
signal \ALU.N_706_cascade_\ : std_logic;
signal \ALU.N_754\ : std_logic;
signal \ALU.aluOut_7_cascade_\ : std_logic;
signal \ALU.a7_b_0_6\ : std_logic;
signal \ALU.m271_nsZ0Z_1\ : std_logic;
signal \ALU.madd_20_0_cascade_\ : std_logic;
signal \ALU.madd_20\ : std_logic;
signal \ctrlOut_2\ : std_logic;
signal \ALU.N_5_0_cascade_\ : std_logic;
signal \ALU.N_240_0_cascade_\ : std_logic;
signal \ALU.madd_24_0_tz\ : std_logic;
signal \ALU.madd_8_0\ : std_logic;
signal \ALU.madd_5\ : std_logic;
signal \ALU.madd_8_0_cascade_\ : std_logic;
signal \ALU.a7_b_0_cascade_\ : std_logic;
signal \ALU.madd_59\ : std_logic;
signal \ALU.madd_484_5\ : std_logic;
signal \ALU.madd_128_0_tz_0\ : std_logic;
signal \ALU.madd_104\ : std_logic;
signal \ALU.madd_149\ : std_logic;
signal \ALU.madd_128_0_tz\ : std_logic;
signal \ALU.madd_128_0\ : std_logic;
signal \ALU.madd_N_1_i\ : std_logic;
signal \ALU.madd_33\ : std_logic;
signal \ALU.madd_68_0_tz\ : std_logic;
signal \ALU.madd_68\ : std_logic;
signal \ALU.madd_89_0\ : std_logic;
signal \ALU.madd_68_cascade_\ : std_logic;
signal \ALU.a7_b_1\ : std_logic;
signal \ALU.madd_108\ : std_logic;
signal \ALU.madd_108_cascade_\ : std_logic;
signal \ALU.madd_134\ : std_logic;
signal \ALU.madd_153\ : std_logic;
signal \FTDI.N_201_2\ : std_logic;
signal \INVFTDI.RXreadyC_net\ : std_logic;
signal \aluOperation_3\ : std_logic;
signal \ALU.m681Z0Z_1_cascade_\ : std_logic;
signal \ALU.N_730_mux\ : std_logic;
signal \FTDI.N_28\ : std_logic;
signal \ALU.a_15_m1_0\ : std_logic;
signal \ALU.a_15_m4_ns_1_0_cascade_\ : std_logic;
signal \ALU.a_15_m4_0_cascade_\ : std_logic;
signal \ALU.a_15_m3_0\ : std_logic;
signal \ALU.a_15_m4_bm_1Z0Z_8\ : std_logic;
signal \ALU.a_15_m0_0\ : std_logic;
signal i53_mux_0 : std_logic;
signal \ALU.N_273_0\ : std_logic;
signal \ALU.N_461\ : std_logic;
signal \ALU.N_474\ : std_logic;
signal \ALU.N_530_cascade_\ : std_logic;
signal \ALU.N_635\ : std_logic;
signal \ALU.d_RNIP8ITN1Z0Z_5_cascade_\ : std_logic;
signal \ALU.d_RNILBFG4Z0Z_2\ : std_logic;
signal \ALU.a_15_m3_2_cascade_\ : std_logic;
signal \ALU.d_RNIE937BZ0Z_0_cascade_\ : std_logic;
signal \ALU.a_15_m4_2\ : std_logic;
signal \ALU.N_257\ : std_logic;
signal \ALU.N_249_cascade_\ : std_logic;
signal \ALU.N_253\ : std_logic;
signal \ALU.c_RNIUGCLVZ0Z_11_cascade_\ : std_logic;
signal \ALU.N_415\ : std_logic;
signal \ALU.N_310\ : std_logic;
signal \ALU.lshift_3_ns_1_4_cascade_\ : std_logic;
signal \ALU.N_220\ : std_logic;
signal \ALU.N_250\ : std_logic;
signal \ALU.N_250_cascade_\ : std_logic;
signal \ALU.N_254\ : std_logic;
signal \ALU.N_218\ : std_logic;
signal \ALU.N_218_cascade_\ : std_logic;
signal \ALU.N_361_cascade_\ : std_logic;
signal \ALU.N_252\ : std_logic;
signal \ALU.m270_nsZ0Z_1_cascade_\ : std_logic;
signal \ctrlOut_12\ : std_logic;
signal \ctrlOut_15\ : std_logic;
signal \ALU.N_7_0_cascade_\ : std_logic;
signal \ALU.N_179_0\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_13_cascade_\ : std_logic;
signal \ALU.operand2_9\ : std_logic;
signal \ALU.N_205_0\ : std_logic;
signal \ALU.operand2_9_cascade_\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_9_cascade_\ : std_logic;
signal \ALU.d_RNIO7LUZ0Z_13_cascade_\ : std_logic;
signal \ALU.operand2_13_cascade_\ : std_logic;
signal \ALU.N_177_0_cascade_\ : std_logic;
signal \ALU.madd_484_3\ : std_logic;
signal \ALU.madd_484_1\ : std_logic;
signal \ALU.madd_484_2_cascade_\ : std_logic;
signal \ALU.madd_484_0\ : std_logic;
signal \ALU.madd_484_12\ : std_logic;
signal \ALU.a0_b_11\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \ALU.un2_addsub_cry_0\ : std_logic;
signal \ALU.d_RNIEDJEAZ0Z_2\ : std_logic;
signal \ALU.N_240_0_i\ : std_logic;
signal \ALU.un2_addsub_cry_1\ : std_logic;
signal \ALU.un2_addsub_cry_2\ : std_logic;
signal \ALU.un2_addsub_cry_3\ : std_logic;
signal \ALU.d_RNIVR3QAZ0Z_5\ : std_logic;
signal \ALU.un2_addsub_cry_4\ : std_logic;
signal \ALU.d_RNIGLK5BZ0Z_6\ : std_logic;
signal \ALU.un2_addsub_cry_5\ : std_logic;
signal \ALU.d_RNITAM9DZ0Z_7\ : std_logic;
signal \ALU.un2_addsub_cry_6\ : std_logic;
signal \ALU.un2_addsub_cry_7\ : std_logic;
signal \ALU.N_201_0\ : std_logic;
signal \ALU.d_RNIQ74VBZ0Z_8\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \ALU.d_RNI6B7KDZ0Z_9\ : std_logic;
signal \ALU.un2_addsub_cry_8\ : std_logic;
signal \ALU.N_192_0_i\ : std_logic;
signal \ALU.un2_addsub_cry_9\ : std_logic;
signal \ALU.un2_addsub_cry_10\ : std_logic;
signal \ALU.N_180_0_i\ : std_logic;
signal \ALU.un2_addsub_cry_11\ : std_logic;
signal \ALU.un2_addsub_cry_12\ : std_logic;
signal \ALU.N_171_0\ : std_logic;
signal \ALU.d_RNI1M3JEZ0Z_14\ : std_logic;
signal \ALU.un2_addsub_cry_13\ : std_logic;
signal \ALU.un2_addsub_cry_14\ : std_logic;
signal \ALU.g0_7_a3_0Z0Z_0\ : std_logic;
signal \ALU.N_8_1_cascade_\ : std_logic;
signal \ALU.g0_2Z0Z_1\ : std_logic;
signal \ALU.g0_7_m4_0_1_cascade_\ : std_logic;
signal \ALU.N_9_2\ : std_logic;
signal \ALU.dout_3_ns_1_0_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_0_cascade_\ : std_logic;
signal \ALU.N_747_cascade_\ : std_logic;
signal \ALU.aluOut_0_cascade_\ : std_logic;
signal \ALU.g0_0_0_N_2L1\ : std_logic;
signal \ALU.dout_3_ns_1_7\ : std_logic;
signal \ALU.a_15_m5_0\ : std_logic;
signal \ALU.d_RNI9BO713Z0Z_0_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_0_cascade_\ : std_logic;
signal \ctrlOut_0\ : std_logic;
signal \ALU.operand2_0_cascade_\ : std_logic;
signal \ALU.hZ0Z_0\ : std_logic;
signal \ALU.d_RNIE4R7Z0Z_0\ : std_logic;
signal \ALU.g_RNIT0COZ0Z_1_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_1_cascade_\ : std_logic;
signal \ALU.e_RNIPKVJZ0Z_1\ : std_logic;
signal \ALU.madd_4\ : std_logic;
signal \ALU.madd_12_0_tz\ : std_logic;
signal \ALU.dout_6_ns_1_15_cascade_\ : std_logic;
signal \ALU.N_752_cascade_\ : std_logic;
signal \ALU.dout_3_ns_1_5_cascade_\ : std_logic;
signal \ALU.N_704\ : std_logic;
signal \ALU.un2_addsub_axb_4_cascade_\ : std_logic;
signal \ALU.d_RNI312TBZ0Z_4\ : std_logic;
signal \ALU.N_223_0\ : std_logic;
signal \ALU.operand2_5\ : std_logic;
signal \ALU.a3_b_5_cascade_\ : std_logic;
signal \ALU.madd_94\ : std_logic;
signal \ALU.a4_b_4\ : std_logic;
signal \ALU.a3_b_5\ : std_logic;
signal \ALU.a4_b_4_cascade_\ : std_logic;
signal \ALU.madd_98\ : std_logic;
signal \ALU.N_207_0\ : std_logic;
signal \ALU.madd_98_cascade_\ : std_logic;
signal \ALU.madd_93\ : std_logic;
signal \ALU.madd_139\ : std_logic;
signal \RX_c\ : std_logic;
signal \RXready\ : std_logic;
signal \ctrlOut_1\ : std_logic;
signal \ALU.N_41_0_0_cascade_\ : std_logic;
signal \ALU.rshift_3_ns_1_5\ : std_logic;
signal \ALU.N_473_cascade_\ : std_logic;
signal \ALU.m42_nsZ0Z_1\ : std_logic;
signal \testWordZ0Z_1\ : std_logic;
signal \testWordZ0Z_4\ : std_logic;
signal \testWordZ0Z_2\ : std_logic;
signal \testWordZ0Z_3\ : std_logic;
signal \ALU.N_469_cascade_\ : std_logic;
signal \ALU.N_473\ : std_logic;
signal \ALU.rshift_15_ns_1_1_cascade_\ : std_logic;
signal \N_305_0\ : std_logic;
signal \CONTROL.aluParams_cnvZ0Z_0\ : std_logic;
signal \ALU.rshift_3_ns_1_9_cascade_\ : std_logic;
signal \ALU.rshift_3_ns_1_1\ : std_logic;
signal \ALU.d_RNINEO9E_0Z0Z_1\ : std_logic;
signal \ALU.N_217\ : std_logic;
signal \ALU.lshift_7_ns_1_9\ : std_logic;
signal \ALU.N_311_cascade_\ : std_logic;
signal \ALU.lshift_9_cascade_\ : std_logic;
signal \ALU.a_15_m2_9\ : std_logic;
signal \ALU.N_292_0\ : std_logic;
signal \ALU.rshift_1\ : std_logic;
signal \ALU.d_RNIA28GU1Z0Z_1_cascade_\ : std_logic;
signal \ALU.d_RNIJ1PCQZ0Z_1\ : std_logic;
signal \ALU.N_225\ : std_logic;
signal \ALU.N_223\ : std_logic;
signal \ALU.N_221\ : std_logic;
signal \ALU.lshift_7_ns_1_13_cascade_\ : std_logic;
signal \ALU.N_219\ : std_logic;
signal \ALU.N_315_cascade_\ : std_logic;
signal \ALU.lshift_13_cascade_\ : std_logic;
signal \ALU.a_15_m2_13\ : std_logic;
signal \ALU.a_15_m4_13_cascade_\ : std_logic;
signal \ALU.N_247\ : std_logic;
signal \ALU.lshift_15_ns_1_15\ : std_logic;
signal \ALU.N_416\ : std_logic;
signal \ALU.N_377\ : std_logic;
signal \ALU.N_377_cascade_\ : std_logic;
signal \ALU.N_216\ : std_logic;
signal \ALU.N_404\ : std_logic;
signal \ALU.N_246\ : std_logic;
signal \ALU.N_376_cascade_\ : std_logic;
signal \ALU.d_RNIEBMRAZ0Z_0_cascade_\ : std_logic;
signal \ALU.d_RNI1GH4VZ0Z_7\ : std_logic;
signal \ALU.N_468\ : std_logic;
signal \ALU.a1_b_3\ : std_logic;
signal \ALU.a0_b_4\ : std_logic;
signal \ALU.a1_b_3_cascade_\ : std_logic;
signal \ALU.madd_0\ : std_logic;
signal \ALU.a0_b_3\ : std_logic;
signal \ALU.N_375\ : std_logic;
signal \ALU.rshift_3_ns_1_0\ : std_logic;
signal \ALU.N_249\ : std_logic;
signal \ALU.N_245\ : std_logic;
signal \ALU.lshift_10\ : std_logic;
signal \ALU.a_15_m3_10\ : std_logic;
signal \ALU.a_15_m4_10_cascade_\ : std_logic;
signal \ALU.a_15_m2_10\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_10\ : std_logic;
signal \ALU.un2_addsub_cry_9_c_RNIVCOFAZ0\ : std_logic;
signal \un9_addsub_cry_9_c_RNI8H83V_cascade_\ : std_logic;
signal \c_RNI5V90O2_10\ : std_logic;
signal \aluOperation_RNINNN4N3_0_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_11_cascade_\ : std_logic;
signal \ALU.dout_3_ns_1_11_cascade_\ : std_logic;
signal \ALU.N_758\ : std_logic;
signal \ALU.N_710_cascade_\ : std_logic;
signal \ALU.aluOut_11_cascade_\ : std_logic;
signal \ALU.madd_484_6\ : std_logic;
signal \ALU.un2_addsub_axb_1_cascade_\ : std_logic;
signal \ALU.d_RNIC4AT9Z0Z_1\ : std_logic;
signal \ALU.dout_7_ns_1_1_cascade_\ : std_logic;
signal \ALU.N_247_0\ : std_logic;
signal \ALU.operand2_1\ : std_logic;
signal \ALU.N_249_0\ : std_logic;
signal \ALU.N_249_0_cascade_\ : std_logic;
signal \ALU.d_RNI61SHAZ0Z_1_cascade_\ : std_logic;
signal \ALU.d_RNIJM067Z0Z_1\ : std_logic;
signal \ALU.a_15_m2_1\ : std_logic;
signal \ALU.g_RNIK6LLZ0Z_4_cascade_\ : std_logic;
signal \ALU.e_RNIGQ8HZ0Z_4\ : std_logic;
signal \ALU.a1_b_4\ : std_logic;
signal \ALU.a2_b_4\ : std_logic;
signal \ALU.operand2_7_ns_1_4\ : std_logic;
signal \ALU.operand2_4\ : std_logic;
signal \ALU.N_229_0\ : std_logic;
signal \ALU.operand2_4_cascade_\ : std_logic;
signal \ALU.N_231_0_cascade_\ : std_logic;
signal \ALU.madd_93_0\ : std_logic;
signal \ALU.aZ0Z_10\ : std_logic;
signal \ALU.dout_3_ns_1_10_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_10_cascade_\ : std_logic;
signal \ALU.N_757_cascade_\ : std_logic;
signal \ALU.N_709\ : std_logic;
signal \ALU.dout_6_ns_1_5\ : std_logic;
signal \ALU.N_865_cascade_\ : std_logic;
signal \ALU.operand2_3_ns_1_6_cascade_\ : std_logic;
signal \ALU.N_817\ : std_logic;
signal \ALU.a6_b_6\ : std_logic;
signal \ALU.a3_b_6\ : std_logic;
signal \ALU.operand2_6_ns_1_6\ : std_logic;
signal \ALU.N_750_cascade_\ : std_logic;
signal \ALU.operand2_3_cascade_\ : std_logic;
signal \ALU.a3_b_3\ : std_logic;
signal \aluReadBus_rep1\ : std_logic;
signal \ALU.a2_b_3\ : std_logic;
signal \ALU.operand2_3\ : std_logic;
signal \ALU.N_235_0\ : std_logic;
signal \ALU.un2_addsub_axb_3\ : std_logic;
signal \ALU.d_RNIDK21BZ0Z_3\ : std_logic;
signal \ALU.dout_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.N_702\ : std_logic;
signal \ALU.g_RNII4LLZ0Z_3\ : std_logic;
signal \ALU.e_RNITOVJZ0Z_3_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_3\ : std_logic;
signal \ALU.un2_addsub_cry_6_c_RNIL4LMIZ0\ : std_logic;
signal \ALU.a7_b_0\ : std_logic;
signal \ALU.a5_b_2\ : std_logic;
signal \ALU.madd_63\ : std_logic;
signal \ALU.a2_b_1\ : std_logic;
signal \ALU.a3_b_0\ : std_logic;
signal \ALU.a1_b_2\ : std_logic;
signal \ALU.d_RNI2B0LZ0Z_9\ : std_logic;
signal \ALU.hZ0Z_10\ : std_logic;
signal \ALU.d_RNII1LUZ0Z_10\ : std_logic;
signal \ALU.d_RNIO00LZ0Z_4\ : std_logic;
signal \FTDI.RXstateZ0Z_2\ : std_logic;
signal \FTDI.N_23_cascade_\ : std_logic;
signal \FTDI.RXstateZ0Z_1\ : std_logic;
signal \FTDI.m13_ns_1\ : std_logic;
signal \FTDI.RXstateZ0Z_0\ : std_logic;
signal \FTDI.RXstateZ0Z_3\ : std_logic;
signal \INVFTDI.gap_0C_net\ : std_logic;
signal \ALU.a_15_sm0_cascade_\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_12_cascade_\ : std_logic;
signal \ALU.log_2_sqmuxa\ : std_logic;
signal \ALU.a_15_m4_bm_1Z0Z_2_cascade_\ : std_logic;
signal \ALU.d_RNIII58AZ0Z_2\ : std_logic;
signal \ALU.rshift_3_ns_1_2_cascade_\ : std_logic;
signal \ALU.N_470\ : std_logic;
signal \ALU.N_376\ : std_logic;
signal \ALU.N_589_cascade_\ : std_logic;
signal \ALU.rshift_1_13_cascade_\ : std_logic;
signal \ALU.a_15_m3_13\ : std_logic;
signal \ALU.N_576_cascade_\ : std_logic;
signal \ALU.N_636_cascade_\ : std_logic;
signal \ALU.N_272_0\ : std_logic;
signal \ALU.N_264_0\ : std_logic;
signal \ALU.aluOut_12\ : std_logic;
signal \ALU.N_462\ : std_logic;
signal \ALU.N_270_0\ : std_logic;
signal \aluReadBus_fast\ : std_logic;
signal \ALU.N_175_0\ : std_logic;
signal \ALU.N_175_0_cascade_\ : std_logic;
signal \ALU.operand2_13\ : std_logic;
signal \ALU.un2_addsub_axb_13_cascade_\ : std_logic;
signal \ALU.N_177_0\ : std_logic;
signal \ALU.d_RNI9FOTEZ0Z_13\ : std_logic;
signal \ctrlOut_11\ : std_logic;
signal \ALU.N_186_0_i\ : std_logic;
signal \ALU.N_186_0_i_cascade_\ : std_logic;
signal \ALU.c_RNIA7OEEZ0Z_11\ : std_logic;
signal \RXbuffer_5\ : std_logic;
signal \ALU.hZ0Z_12\ : std_logic;
signal \ALU.c_RNIJ949Z0Z_12_cascade_\ : std_logic;
signal \ALU.a_RNIFPBOZ0Z_12\ : std_logic;
signal \ALU.d_RNIM5LUZ0Z_12\ : std_logic;
signal \ALU.operand2_7_ns_1_12_cascade_\ : std_logic;
signal \ALU.operand2_12\ : std_logic;
signal \ALU.d_RNICJE9BZ0Z_8\ : std_logic;
signal \ALU.d_RNIEUKR11Z0Z_0\ : std_logic;
signal \ALU.a_15_m3_8\ : std_logic;
signal \ALU.a_15_m4_8_cascade_\ : std_logic;
signal \ALU.a_15_m5_8\ : std_logic;
signal \ALU.fZ0Z_8\ : std_logic;
signal \ALU.dZ0Z_8\ : std_logic;
signal \ALU.operand2_6_ns_1_8_cascade_\ : std_logic;
signal \ALU.N_867\ : std_logic;
signal \ALU.hZ0Z_8\ : std_logic;
signal \ALU.fZ0Z_15\ : std_logic;
signal \ALU.madd_cry_0_ma\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \ALU.madd_cry_1_ma\ : std_logic;
signal \ALU.madd_cry_0\ : std_logic;
signal \ALU.madd_axb_2_l_fx\ : std_logic;
signal \ALU.madd_6\ : std_logic;
signal \ALU.madd_cry_1\ : std_logic;
signal \ALU.madd_13\ : std_logic;
signal \ALU.madd_18\ : std_logic;
signal \ALU.madd_cry_2\ : std_logic;
signal \ALU.madd_axb_4_l_fx\ : std_logic;
signal \ALU.madd_30\ : std_logic;
signal \ALU.madd_cry_3\ : std_logic;
signal \ALU.madd_52\ : std_logic;
signal \ALU.madd_axb_5_l_fx\ : std_logic;
signal \ALU.madd_cry_4\ : std_logic;
signal \ALU.madd_cry_5\ : std_logic;
signal \ALU.madd_axb_7\ : std_logic;
signal \ALU.madd_cry_6_THRU_CO\ : std_logic;
signal \ALU.madd_cry_6\ : std_logic;
signal \ALU.madd_cry_7\ : std_logic;
signal \ALU.madd_axb_8_l_fx\ : std_logic;
signal \ALU.madd_159\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \ALU.madd_cry_9_ma\ : std_logic;
signal \ALU.madd_axb_9_l_ofx\ : std_logic;
signal \ALU.madd_cry_8\ : std_logic;
signal \ALU.madd_cry_10_ma\ : std_logic;
signal \ALU.madd_axb_10_l_ofx\ : std_logic;
signal \ALU.madd_cry_9\ : std_logic;
signal \ALU.madd_axb_11\ : std_logic;
signal \ALU.madd_cry_10\ : std_logic;
signal \ALU.madd_axb_12_l_fx\ : std_logic;
signal \ALU.madd_360\ : std_logic;
signal \ALU.madd_cry_11\ : std_logic;
signal \ALU.madd_cry_13_ma\ : std_logic;
signal \ALU.madd_axb_13_l_ofx\ : std_logic;
signal \ALU.madd_cry_12\ : std_logic;
signal \ALU.madd_axb_14\ : std_logic;
signal \ALU.madd_cry_13\ : std_logic;
signal \ALU.operand2_6\ : std_logic;
signal \aluReadBus\ : std_logic;
signal \ALU.N_217_0\ : std_logic;
signal \ALU.dout_3_ns_1_15_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_2_cascade_\ : std_logic;
signal \ALU.N_749_cascade_\ : std_logic;
signal \ALU.N_701\ : std_logic;
signal \ALU.dout_3_ns_1_2\ : std_logic;
signal \ALU.dout_6_ns_1_7\ : std_logic;
signal \ALU.f_RNIQQJ01Z0Z_7\ : std_logic;
signal \testWordZ0Z_8\ : std_logic;
signal \ALU.fZ0Z_10\ : std_logic;
signal \ALU.b_RNIEHSD1Z0Z_10\ : std_logic;
signal \ALU.dout_3_ns_1_4\ : std_logic;
signal \ALU.eZ0Z_4\ : std_logic;
signal \ALU.e_RNIS97JZ0Z_1\ : std_logic;
signal \ALU.eZ0Z_1\ : std_logic;
signal \ALU.g_RNI0MJNZ0Z_1\ : std_logic;
signal \ALU.dout_6_ns_1_3\ : std_logic;
signal \aluOperand1_2_rep1\ : std_logic;
signal \ALU.dout_6_ns_1_4\ : std_logic;
signal \ALU.N_747\ : std_logic;
signal \ALU.N_699\ : std_logic;
signal \ALU.N_404_1\ : std_logic;
signal \ALU.dout_6_ns_1_6\ : std_logic;
signal \ALU.N_753_cascade_\ : std_logic;
signal \testWordZ0Z_9\ : std_logic;
signal \aluOperand1_fast_1\ : std_logic;
signal \aluOperand1_fast_2\ : std_logic;
signal \ALU.dout_3_ns_1_6_cascade_\ : std_logic;
signal \ALU.N_705\ : std_logic;
signal \testWordZ0Z_7\ : std_logic;
signal \CONTROL.operand1_cnvZ0Z_0\ : std_logic;
signal \ALU.c_RNI72MICZ0Z_15_cascade_\ : std_logic;
signal \ALU.d_RNI4HG101Z0Z_7\ : std_logic;
signal \INVFTDI.baudAcc_0C_net\ : std_logic;
signal \ALU.aluOut_10\ : std_logic;
signal \ALU.N_475_cascade_\ : std_logic;
signal \ALU.rshift_7\ : std_logic;
signal \ALU.rshift_15_ns_1_7\ : std_logic;
signal \ALU.rshift_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.N_471_cascade_\ : std_logic;
signal \ALU.N_475\ : std_logic;
signal \ALU.rshift_3_ns_1_7\ : std_logic;
signal \ALU.N_576\ : std_logic;
signal \ALU.a_15_m5_5_cascade_\ : std_logic;
signal \ALU.mult_5\ : std_logic;
signal \ALU.d_RNIPFIBI1Z0Z_9\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_5_cascade_\ : std_logic;
signal \ALU.N_225_0\ : std_logic;
signal \ALU.a_15_m2_5_cascade_\ : std_logic;
signal \ALU.N_420\ : std_logic;
signal \ALU.a_15_m4_5\ : std_logic;
signal a_4 : std_logic;
signal a_6 : std_logic;
signal a_7 : std_logic;
signal \ALU.a_15_m2_12\ : std_logic;
signal \ALU.a_15_m4_12_cascade_\ : std_logic;
signal \ALU.un2_addsub_cry_11_c_RNII7OFZ0Z9\ : std_logic;
signal \un2_addsub_cry_11_c_RNIQ9LMU_cascade_\ : std_logic;
signal \c_RNIC8RDN2_12\ : std_logic;
signal \aluOperation_RNIGPL5M3_0_cascade_\ : std_logic;
signal \ALU.aZ0Z_12\ : std_logic;
signal \ALU.N_271_0\ : std_logic;
signal \ALU.a_15_m3_12\ : std_logic;
signal \ALU.N_314\ : std_logic;
signal \ALU.lshift_12\ : std_logic;
signal \ALU.fZ0Z_9\ : std_logic;
signal \ALU.bZ0Z_9\ : std_logic;
signal \ALU.f_RNIUUJ01Z0Z_9\ : std_logic;
signal \ALU.bZ0Z_12\ : std_logic;
signal \ALU.fZ0Z_12\ : std_logic;
signal \ALU.b_RNIILSD1Z0Z_12\ : std_logic;
signal \ALU.fZ0Z_14\ : std_logic;
signal \ALU.bZ0Z_14\ : std_logic;
signal \ALU.g0_3_1_cascade_\ : std_logic;
signal \ALU.N_703_0_0\ : std_logic;
signal \ALU.N_4\ : std_logic;
signal \ALU.N_5\ : std_logic;
signal \ALU.fZ0Z_11\ : std_logic;
signal \ALU.bZ0Z_11\ : std_logic;
signal \ALU.b_RNIKNSD1Z0Z_13\ : std_logic;
signal \ALU.dZ0Z_10\ : std_logic;
signal \ALU.dZ0Z_12\ : std_logic;
signal \ALU.eZ0Z_10\ : std_logic;
signal \ALU.eZ0Z_12\ : std_logic;
signal \ALU.d_RNIPER7Z0Z_5\ : std_logic;
signal \ALU.bZ0Z_10\ : std_logic;
signal \ALU.bZ0Z_15\ : std_logic;
signal \ALU.un2_addsub_cry_12_c_RNIUL1GKZ0\ : std_logic;
signal \un2_addsub_cry_12_c_RNIG3PMU_cascade_\ : std_logic;
signal \c_RNI88B4N2_13\ : std_logic;
signal \aluOperation_RNI2J9SL3_0_cascade_\ : std_logic;
signal \ALU.mult_2\ : std_logic;
signal \ALU.a_15_m5_2\ : std_logic;
signal \ALU.d_RNIIFMN04Z0Z_2_cascade_\ : std_logic;
signal \ALU.eZ0Z_3\ : std_logic;
signal \ALU.eZ0Z_6\ : std_logic;
signal \ALU.eZ0Z_7\ : std_logic;
signal \ALU.eZ0Z_2\ : std_logic;
signal a_2 : std_logic;
signal \ALU.g_RNIV2COZ0Z_2_cascade_\ : std_logic;
signal \ALU.e_RNIRMVJZ0Z_2\ : std_logic;
signal \ALU.operand2_7_ns_1_2_cascade_\ : std_logic;
signal \ALU.operand2_2\ : std_logic;
signal \ALU.eZ0Z_0\ : std_logic;
signal a_0 : std_logic;
signal \ALU.e_RNINIVJZ0Z_0\ : std_logic;
signal \ALU.g_RNIM8LLZ0Z_5\ : std_logic;
signal \ALU.e_RNI1TVJZ0Z_5_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_5\ : std_logic;
signal \ALU.eZ0Z_5\ : std_logic;
signal \ALU.g_RNIRUBOZ0Z_0\ : std_logic;
signal \ALU.d_RNIG6R7Z0Z_1\ : std_logic;
signal \ALU.d_RNI45J9Z0Z_1\ : std_logic;
signal \ALU.d_RNII8R7Z0Z_2\ : std_logic;
signal \ALU.cZ0Z_0\ : std_logic;
signal \ALU.cZ0Z_1\ : std_logic;
signal \ALU.cZ0Z_2\ : std_logic;
signal \ALU.cZ0Z_3\ : std_logic;
signal \ALU.cZ0Z_4\ : std_logic;
signal \ALU.cZ0Z_5\ : std_logic;
signal \ALU.cZ0Z_6\ : std_logic;
signal \ALU.dZ0Z_4\ : std_logic;
signal \ALU.gZ0Z_6\ : std_logic;
signal \FTDI.gapZ0Z_2\ : std_logic;
signal \FTDI.gapZ0Z_0\ : std_logic;
signal \FTDI.gap8\ : std_logic;
signal \FTDI.gapZ0Z_1\ : std_logic;
signal \INVFTDI.gap_2C_net\ : std_logic;
signal \FTDI.TXstate_e_1_0\ : std_logic;
signal \FTDI.N_169_0_cascade_\ : std_logic;
signal \FTDI.N_169_0\ : std_logic;
signal \FTDI.TXstate_cnst_0_0_2_cascade_\ : std_logic;
signal \INVFTDI.TXstate_0C_net\ : std_logic;
signal \FTDI.N_217_0_cascade_\ : std_logic;
signal \FTDI.N_216_0\ : std_logic;
signal \FTDI.TXready_cascade_\ : std_logic;
signal \FTDI.baudAccZ0Z_0\ : std_logic;
signal \FTDI.baudAccZ0Z_1\ : std_logic;
signal \ALU.N_290_0\ : std_logic;
signal \ALU.rshift_5\ : std_logic;
signal \ALU.a_15_m3_5\ : std_logic;
signal \FTDI.TXstateZ1Z_0\ : std_logic;
signal \FTDI.TXstateZ1Z_1\ : std_logic;
signal \FTDI.N_170_0\ : std_logic;
signal \FTDI.TXstate_e_1_3_cascade_\ : std_logic;
signal \INVFTDI.baudAcc_1C_net\ : std_logic;
signal \ALU.N_11_0\ : std_logic;
signal \ALU.N_5_0\ : std_logic;
signal \ALU.c_RNI1OCN4Z0Z_15_cascade_\ : std_logic;
signal \ALU.N_762\ : std_logic;
signal \ALU.N_714\ : std_logic;
signal \ALU.N_621_1_cascade_\ : std_logic;
signal \ALU.N_589\ : std_logic;
signal \ALU.N_621_1\ : std_logic;
signal \ALU.c_RNI4JFV4_0Z0Z_15\ : std_logic;
signal \ALU.N_274_0\ : std_logic;
signal \ALU.d_RNI36KJ21Z0Z_9\ : std_logic;
signal \FTDI.TXready\ : std_logic;
signal \FTDI.baudAccZ0Z_2\ : std_logic;
signal \TXstartZ0\ : std_logic;
signal \testStateZ0Z_0\ : std_logic;
signal \ctrlOut_13\ : std_logic;
signal \busState_2\ : std_logic;
signal \aluReadBus_rep2\ : std_logic;
signal \busState_0\ : std_logic;
signal \ALU.N_9_1\ : std_logic;
signal \testStateZ0Z_2\ : std_logic;
signal \testState_i_2\ : std_logic;
signal \ALU.eZ0Z_14\ : std_logic;
signal \ALU.un2_addsub_cry_13_c_RNINVE5KZ0\ : std_logic;
signal \un2_addsub_cry_13_c_RNI2LH1U_cascade_\ : std_logic;
signal \c_RNIFCGVL2_14\ : std_logic;
signal \aluOperation_RNIR872K3_0_cascade_\ : std_logic;
signal \ALU.a_RNIJTBOZ0Z_14\ : std_logic;
signal \ALU.operand2_7_ns_1_14_cascade_\ : std_logic;
signal \ALU.b_RNIMPSD1Z0Z_14\ : std_logic;
signal \ALU.operand2_14\ : std_logic;
signal \ALU.hZ0Z_14\ : std_logic;
signal \ALU.dZ0Z_14\ : std_logic;
signal \ALU.d_RNIQ9LUZ0Z_14\ : std_logic;
signal \ALU.un2_addsub_cry_7_c_RNIL8JHGZ0\ : std_logic;
signal \ALU.aZ0Z_8\ : std_logic;
signal \aluOperand2_fast_1\ : std_logic;
signal \ALU.eZ0Z_8\ : std_logic;
signal \ALU.gZ0Z_8\ : std_logic;
signal \ALU.cZ0Z_8\ : std_logic;
signal \ALU.operand2_3_ns_1_8_cascade_\ : std_logic;
signal \ALU.N_819\ : std_logic;
signal \ALU.addsub_0_sqmuxa_cascade_\ : std_logic;
signal \ALU.un2_addsub_cry_8_c_RNIKR81JZ0\ : std_logic;
signal \ALU.un9_addsub_cry_8_c_RNIKTS9SZ0_cascade_\ : std_logic;
signal \ALU.a_15_m5_9\ : std_logic;
signal \ALU.a_15_ns_1_9_cascade_\ : std_logic;
signal \ALU.eZ0Z_11\ : std_logic;
signal \aluOperand2_0_rep1\ : std_logic;
signal \ALU.a_RNICNBOZ0Z_11_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_11_cascade_\ : std_logic;
signal \ALU.b_RNIGJSD1Z0Z_11\ : std_logic;
signal \ALU.operand2_11\ : std_logic;
signal \ALU.dZ0Z_11\ : std_logic;
signal \ALU.d_RNIK3LUZ0Z_11\ : std_logic;
signal \ALU.hZ0Z_11\ : std_logic;
signal \ALU.c_RNIG749Z0Z_11\ : std_logic;
signal \ALU.a_RNIHRBOZ0Z_13_cascade_\ : std_logic;
signal \ALU.c_RNILB49Z0Z_13\ : std_logic;
signal \ALU.operand2_7_ns_1_13\ : std_logic;
signal \ALU.eZ0Z_15\ : std_logic;
signal \ALU.a_RNILVBOZ0Z_15_cascade_\ : std_logic;
signal \ALU.c_RNIPF49Z0Z_15\ : std_logic;
signal \ALU.operand2_7_ns_1_15_cascade_\ : std_logic;
signal \ALU.b_RNIORSD1Z0Z_15\ : std_logic;
signal \ALU.operand2_15\ : std_logic;
signal \ALU.cZ0Z_11\ : std_logic;
signal \ALU.cZ0Z_12\ : std_logic;
signal \ALU.cZ0Z_14\ : std_logic;
signal \ALU.c_RNIND49Z0Z_14\ : std_logic;
signal \ALU.cZ0Z_15\ : std_logic;
signal \ALU.c_cnvZ0Z_0\ : std_logic;
signal \ALU.hZ0Z_1\ : std_logic;
signal \ALU.hZ0Z_2\ : std_logic;
signal \ALU.hZ0Z_5\ : std_logic;
signal \ALU.aZ0Z_14\ : std_logic;
signal \ALU.aZ0Z_15\ : std_logic;
signal \ALU.f_RNI0P6LZ0Z_1\ : std_logic;
signal \ALU.f_RNICQEJZ0Z_1\ : std_logic;
signal \ALU.cZ0Z_7\ : std_logic;
signal \ALU.g_RNIQCLLZ0Z_7\ : std_logic;
signal \ALU.f_RNIL2FJZ0Z_5\ : std_logic;
signal \ALU.m286_bmZ0\ : std_logic;
signal \ALU.m286_amZ0\ : std_logic;
signal \ALU.f_RNIAOEJZ0Z_0\ : std_logic;
signal \aluOperand2_fast_0\ : std_logic;
signal \aluOperand2_2_rep1\ : std_logic;
signal \ALU.bZ0Z_2\ : std_logic;
signal \ALU.f_RNIESEJZ0Z_2\ : std_logic;
signal \ALU.gZ0Z_0\ : std_logic;
signal \ALU.gZ0Z_1\ : std_logic;
signal \ALU.gZ0Z_2\ : std_logic;
signal \ALU.gZ0Z_3\ : std_logic;
signal \ALU.gZ0Z_4\ : std_logic;
signal \ALU.gZ0Z_5\ : std_logic;
signal \ALU.gZ0Z_7\ : std_logic;
signal \ALU.N_578\ : std_logic;
signal \ALU.N_477\ : std_logic;
signal \ALU.N_634\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \FTDI.un3_TX_0\ : std_logic;
signal \RXbuffer_4\ : std_logic;
signal \testWordZ0Z_12\ : std_logic;
signal \TXbufferZ0Z_0\ : std_logic;
signal \TXbufferZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_5\ : std_logic;
signal \TXbufferZ0Z_4\ : std_logic;
signal \FTDI.TXshiftZ0Z_4\ : std_logic;
signal \FTDI.TXshiftZ0Z_3\ : std_logic;
signal \TXbufferZ0Z_2\ : std_logic;
signal \TXbufferZ0Z_6\ : std_logic;
signal \FTDI.TXshiftZ0Z_6\ : std_logic;
signal \TXbufferZ0Z_7\ : std_logic;
signal \FTDI.TXshiftZ0Z_7\ : std_logic;
signal \INVFTDI.TXshift_0C_net\ : std_logic;
signal \ALU.un2_addsub_cry_10_c_RNIUS1OJZ0\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_11_cascade_\ : std_logic;
signal \ALU.a_15_m2_11_cascade_\ : std_logic;
signal \ALU.lshift_11\ : std_logic;
signal \ALU.a_15_m4_11_cascade_\ : std_logic;
signal \ALU.a_15_m3_11\ : std_logic;
signal \c_RNID7K8N2_11_cascade_\ : std_logic;
signal \un2_addsub_cry_10_c_RNIEBKOT\ : std_logic;
signal \aluOperation_RNI5QD2L3_0_cascade_\ : std_logic;
signal \ALU.aZ0Z_11\ : std_logic;
signal \ALU.e_cnvZ0Z_0\ : std_logic;
signal \ALU.g_RNIVGLLZ0Z_9_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_9\ : std_logic;
signal \ALU.hZ0Z_9\ : std_logic;
signal \ALU.dZ0Z_9\ : std_logic;
signal \ALU.g0_0_0_m2_1\ : std_logic;
signal \ALU.N_11_cascade_\ : std_logic;
signal \ALU.N_13\ : std_logic;
signal \ALU.cZ0Z_9\ : std_logic;
signal \ALU.g0_0_0_m2_0_1\ : std_logic;
signal \ALU.N_12\ : std_logic;
signal \ALU.aluOut_15\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_15_cascade_\ : std_logic;
signal \ALU.N_7_0\ : std_logic;
signal \ALU.a_15_m2_15_cascade_\ : std_logic;
signal \ALU.lshift_15\ : std_logic;
signal \ALU.a_15_m4_15_cascade_\ : std_logic;
signal \ALU.a_15_m3_15\ : std_logic;
signal \ALU.c_RNIR4QHM2Z0Z_15_cascade_\ : std_logic;
signal \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93_cascade_\ : std_logic;
signal \ALU.hZ0Z_15\ : std_logic;
signal \ALU.dZ0Z_15\ : std_logic;
signal \ALU.d_RNISBLUZ0Z_15\ : std_logic;
signal \CONTROL.aluOperation_cnvZ0Z_0\ : std_logic;
signal \N_723\ : std_logic;
signal \testWordZ0Z_5\ : std_logic;
signal \aluOperation_5\ : std_logic;
signal \ALU.a2_b_0\ : std_logic;
signal \ALU.madd_axb_1_l_ofx\ : std_logic;
signal \aluOperand2_0_rep2\ : std_logic;
signal \aluOperand2_0\ : std_logic;
signal \aluOperand2_1_rep1\ : std_logic;
signal \ALU.cZ0Z_10\ : std_logic;
signal \aluOperand2_fast_2\ : std_logic;
signal \ALU.g0_7_m4_1\ : std_logic;
signal \N_287_0\ : std_logic;
signal \G_566\ : std_logic;
signal \testWordZ0Z_11\ : std_logic;
signal \aluOperand2_1\ : std_logic;
signal \ALU.mult_10\ : std_logic;
signal \aluOperation_RNINNN4N3_0\ : std_logic;
signal \ALU.gZ0Z_10\ : std_logic;
signal \aluOperation_RNI5QD2L3_0\ : std_logic;
signal \ALU.mult_11\ : std_logic;
signal \ALU.gZ0Z_11\ : std_logic;
signal \aluOperation_RNIGPL5M3_0\ : std_logic;
signal \ALU.mult_12\ : std_logic;
signal \ALU.gZ0Z_12\ : std_logic;
signal \aluOperation_RNI2J9SL3_0\ : std_logic;
signal \ALU.mult_13\ : std_logic;
signal \aluOperation_RNIR872K3_0\ : std_logic;
signal \ALU.mult_14\ : std_logic;
signal \ALU.gZ0Z_14\ : std_logic;
signal \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93\ : std_logic;
signal \ALU.mult_15\ : std_logic;
signal \ALU.gZ0Z_15\ : std_logic;
signal \ALU.a_15_ns_1_9\ : std_logic;
signal \ALU.mult_9\ : std_logic;
signal \ALU.gZ0Z_9\ : std_logic;
signal \ALU.g_cnvZ0Z_0\ : std_logic;
signal \ALU.eZ0Z_13\ : std_logic;
signal \ALU.aZ0Z_13\ : std_logic;
signal \aluOperand1_2_rep2\ : std_logic;
signal \aluOperand1_1_rep1\ : std_logic;
signal \ALU.cZ0Z_13\ : std_logic;
signal \ALU.dout_3_ns_1_13_cascade_\ : std_logic;
signal \ALU.gZ0Z_13\ : std_logic;
signal \ALU.bZ0Z_13\ : std_logic;
signal \aluOperand1_1_rep2\ : std_logic;
signal \ALU.fZ0Z_13\ : std_logic;
signal \aluOperand1_2\ : std_logic;
signal \ALU.hZ0Z_13\ : std_logic;
signal \ALU.dZ0Z_13\ : std_logic;
signal \ALU.dout_6_ns_1_13_cascade_\ : std_logic;
signal \aluOperand1_1\ : std_logic;
signal \ALU.N_712\ : std_logic;
signal \ALU.N_760_cascade_\ : std_logic;
signal \aluOperand1_0\ : std_logic;
signal \ALU.aluOut_13_cascade_\ : std_logic;
signal \ALU.a13_b_0\ : std_logic;
signal \ALU.fZ0Z_0\ : std_logic;
signal \ALU.fZ0Z_1\ : std_logic;
signal \ALU.fZ0Z_2\ : std_logic;
signal \ALU.fZ0Z_5\ : std_logic;
signal \ALU.fZ0Z_6\ : std_logic;
signal \ALU.fZ0Z_7\ : std_logic;
signal \ALU.f_cnvZ0Z_0\ : std_logic;
signal \ALU.N_1700_i\ : std_logic;
signal \ALU.d_RNIO75MAZ0Z_0_cascade_\ : std_logic;
signal \ALU.bZ0Z_0\ : std_logic;
signal \ALU.madd_axb_0_l_ofx\ : std_logic;
signal \ALU.mult_1_cascade_\ : std_logic;
signal \ALU.a_15_m5_1\ : std_logic;
signal \ALU.d_RNIEICQ63Z0Z_1_cascade_\ : std_logic;
signal \ALU.bZ0Z_1\ : std_logic;
signal \ALU.d_RNIEICQ63Z0Z_1\ : std_logic;
signal \ALU.dZ0Z_1\ : std_logic;
signal \ALU.hZ0Z_4\ : std_logic;
signal \FTDI.un3_TX_0_i\ : std_logic;
signal \bfn_13_2_0_\ : std_logic;
signal \FTDI.un3_TX_axb_3\ : std_logic;
signal \FTDI.un3_TX_cry_2\ : std_logic;
signal \FTDI.TXshiftZ0Z_0\ : std_logic;
signal \FTDI.un3_TX_cry_3\ : std_logic;
signal \FTDI_TX_0_i\ : std_logic;
signal \ALU.N_361\ : std_logic;
signal \ALU.N_244\ : std_logic;
signal \aluParams_1\ : std_logic;
signal \ALU.N_588\ : std_logic;
signal \aluParams_2\ : std_logic;
signal \ALU.N_590\ : std_logic;
signal \ALU.eZ0Z_9\ : std_logic;
signal \ALU.aZ0Z_9\ : std_logic;
signal \ALU.e_RNIR49HZ0Z_9\ : std_logic;
signal \ALU.N_252_0\ : std_logic;
signal \ALU.aluOut_0\ : std_logic;
signal \ALU.a0_b_2\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \ALU.N_249_0_i\ : std_logic;
signal \ALU.aluOut_1\ : std_logic;
signal \ALU.un9_addsub_cry_0\ : std_logic;
signal \ALU.N_240_0\ : std_logic;
signal \ALU.aluOut_2\ : std_logic;
signal \ALU.un9_addsub_cry_1\ : std_logic;
signal \ALU.N_237_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_2\ : std_logic;
signal \ALU.N_231_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_3\ : std_logic;
signal \ALU.aluOut_5\ : std_logic;
signal \ALU.N_225_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_4\ : std_logic;
signal \ALU.N_219_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_5\ : std_logic;
signal \ALU.N_213_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_6_c_RNI2EFHZ0Z8\ : std_logic;
signal \ALU.un9_addsub_cry_6\ : std_logic;
signal \ALU.un9_addsub_cry_7\ : std_logic;
signal \ALU.aluOut_8\ : std_logic;
signal \ALU.N_201_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_7_c_RNIU7FZ0Z18\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \ALU.aluOut_9\ : std_logic;
signal \ALU.N_207_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_8_c_RNIPV1SZ0Z8\ : std_logic;
signal \ALU.un9_addsub_cry_8\ : std_logic;
signal \ALU.N_192_0\ : std_logic;
signal \ALU.a_RNIV2S0FZ0Z_10\ : std_logic;
signal \ALU.un9_addsub_cry_9_c_RNI22U6KZ0\ : std_logic;
signal \ALU.un9_addsub_cry_9\ : std_logic;
signal \ALU.N_186_0\ : std_logic;
signal \ALU.aluOut_11\ : std_logic;
signal \ALU.un9_addsub_cry_10_c_RNI9C0KZ0Z9\ : std_logic;
signal \ALU.un9_addsub_cry_10\ : std_logic;
signal \ALU.N_180_0\ : std_logic;
signal \ALU.d_RNIFKNTEZ0Z_12\ : std_logic;
signal \ALU.un9_addsub_cry_11_c_RNI10BQKZ0\ : std_logic;
signal \ALU.un9_addsub_cry_11\ : std_logic;
signal \ALU.aluOut_13\ : std_logic;
signal \ALU.N_177_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_12_c_RNIBB5QZ0Z9\ : std_logic;
signal \ALU.un9_addsub_cry_12\ : std_logic;
signal \ALU.aluOut_14\ : std_logic;
signal \ALU.N_171_0_i\ : std_logic;
signal \ALU.un9_addsub_cry_13_c_RNI4JGFZ0Z9\ : std_logic;
signal \ALU.un9_addsub_cry_13\ : std_logic;
signal \ALU.un9_addsub_axb_15\ : std_logic;
signal \ALU.un2_addsub_cry_14_c_RNINOKZ0Z69\ : std_logic;
signal \ALU.un9_addsub_cry_14\ : std_logic;
signal \ALU.un9_addsub_cry_14_c_RNIS374JZ0\ : std_logic;
signal \ALU.c_RNIA9V4LZ0Z_15\ : std_logic;
signal \ALU.d_RNI9DPVUZ0Z_6\ : std_logic;
signal \ALU.rshift_3_cascade_\ : std_logic;
signal \ALU.N_293_0\ : std_logic;
signal \ALU.d_RNI3V2CP1Z0Z_3_cascade_\ : std_logic;
signal \ALU.aluOut_3\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_3\ : std_logic;
signal \ALU.N_237_0\ : std_logic;
signal \ALU.a_15_m2_3_cascade_\ : std_logic;
signal \ALU.lshift_1_3\ : std_logic;
signal \ALU.d_RNI95MLPZ0Z_3\ : std_logic;
signal \ALU.mult_3\ : std_logic;
signal \ALU.a_15_m5_3\ : std_logic;
signal \RXbuffer_2\ : std_logic;
signal \testStateZ0Z_1\ : std_logic;
signal \ALU.N_58_0\ : std_logic;
signal \testWordZ0Z_10\ : std_logic;
signal \testState_i_g_2\ : std_logic;
signal \ALU.un9_addsub_cry_0_c_RNI2UZ0Z096\ : std_logic;
signal \ALU.un2_addsub_cry_0_c_RNI5MA0EZ0\ : std_logic;
signal \ALU.un9_addsub_cry_0_c_RNIEMTLKZ0\ : std_logic;
signal \ALU.un9_addsub_cry_1_c_RNI6TDZ0Z17\ : std_logic;
signal \ALU.un2_addsub_cry_1_c_RNI966GEZ0\ : std_logic;
signal \ALU.un9_addsub_cry_2_c_RNIA3LGZ0Z7\ : std_logic;
signal \ALU.un2_addsub_cry_2_c_RNI5IV5FZ0\ : std_logic;
signal \ALU.un2_addsub_cry_3_c_RNIOGGJGZ0\ : std_logic;
signal \ALU.un9_addsub_cry_3_c_RNI525RZ0Z7\ : std_logic;
signal \ALU.un9_addsub_cry_4_c_RNIL4NZ0Z97\ : std_logic;
signal \ALU.un2_addsub_cry_4_c_RNI284VEZ0\ : std_logic;
signal \ALU.un9_addsub_cry_5_c_RNI6SCFZ0Z7\ : std_logic;
signal \ALU.addsub_0_sqmuxa\ : std_logic;
signal \ALU.un2_addsub_cry_5_c_RNIL7IGFZ0\ : std_logic;
signal \ALU.N_422\ : std_logic;
signal \ALU.d_RNIP43E91Z0Z_7_cascade_\ : std_logic;
signal \ALU.d_RNIT87FA1Z0Z_7\ : std_logic;
signal \ALU.madd_cry_5_THRU_CO\ : std_logic;
signal \ALU.a_15_m5_7_cascade_\ : std_logic;
signal \ALU.madd_axb_6\ : std_logic;
signal \ALU.d_RNIO75MAZ0Z_0\ : std_logic;
signal \ALU.d_RNI9BO713Z0Z_0\ : std_logic;
signal \ALU.dZ0Z_0\ : std_logic;
signal \ALU.un9_addsub_cry_1_c_RNIM56ULZ0\ : std_logic;
signal \ALU.d_RNIIFMN04Z0Z_2\ : std_logic;
signal \ALU.dZ0Z_2\ : std_logic;
signal \ALU.dZ0Z_5\ : std_logic;
signal \ALU.dZ0Z_6\ : std_logic;
signal \ALU.d_cnvZ0Z_0\ : std_logic;
signal \ALU.fZ0Z_3\ : std_logic;
signal \ALU.f_RNIHUEJZ0Z_3\ : std_logic;
signal \ALU.rshift_1_12\ : std_logic;
signal \ALU.N_532\ : std_logic;
signal \aluOperation_4\ : std_logic;
signal \ALU.rshift_4_cascade_\ : std_logic;
signal \ALU.N_289_0\ : std_logic;
signal \ALU.a_15_m3_4_cascade_\ : std_logic;
signal \ALU.aluOut_4\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_4\ : std_logic;
signal \ALU.N_231_0\ : std_logic;
signal \ALU.a_15_m2_4_cascade_\ : std_logic;
signal \ALU.N_419\ : std_logic;
signal \ALU.a_15_m4_4\ : std_logic;
signal \ALU.mult_4\ : std_logic;
signal \ALU.a_15_m5_4\ : std_logic;
signal a_3 : std_logic;
signal \ALU.a_cnvZ0Z_0\ : std_logic;
signal \FTDI.TXshiftZ0Z_2\ : std_logic;
signal \FTDI.TXstateZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_1\ : std_logic;
signal \INVFTDI.TXshift_1C_net\ : std_logic;
signal \FTDI.un1_TXstate_0_sqmuxa_0_i\ : std_logic;
signal a_5 : std_logic;
signal \TXbufferZ0Z_5\ : std_logic;
signal a_1 : std_logic;
signal \TXbufferZ0Z_1\ : std_logic;
signal m326dup : std_logic;
signal \aluParams_3\ : std_logic;
signal \ALU.N_308\ : std_logic;
signal \aluOperation_2\ : std_logic;
signal \ALU.log_0_sqmuxa\ : std_logic;
signal \aluParams_0\ : std_logic;
signal \ALU.aluOut_6\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_6_cascade_\ : std_logic;
signal \ALU.N_219_0\ : std_logic;
signal \ALU.a_15_m2_6\ : std_logic;
signal \ALU.a_15_sm3\ : std_logic;
signal \ALU.d_RNIL01TD1Z0Z_6\ : std_logic;
signal \ALU.d_RNIJ75U41Z0Z_6\ : std_logic;
signal \aluOperation_1\ : std_logic;
signal \ALU.a_15_m5_6_cascade_\ : std_logic;
signal \ALU.mult_6\ : std_logic;
signal \ALU.d_RNILPR7TQZ0Z_6_cascade_\ : std_logic;
signal \ALU.hZ0Z_6\ : std_logic;
signal \ALU.h_cnvZ0Z_0\ : std_logic;
signal \ALU.fZ0Z_4\ : std_logic;
signal \ALU.f_RNIJ0FJZ0Z_4\ : std_logic;
signal \ALU.hZ0Z_7\ : std_logic;
signal \ALU.dZ0Z_7\ : std_logic;
signal \aluOperand2_2\ : std_logic;
signal \ALU.d_RNIU60LZ0Z_7\ : std_logic;
signal \ALU.hZ0Z_3\ : std_logic;
signal \ALU.dZ0Z_3\ : std_logic;
signal \aluOperand2_2_rep2\ : std_logic;
signal \ALU.d_RNILAR7Z0Z_3\ : std_logic;
signal \ALU.un9_addsub_cry_2_c_RNIMN63NZ0\ : std_logic;
signal \ALU.d_RNIE8SJN5Z0Z_3\ : std_logic;
signal \ALU.bZ0Z_3\ : std_logic;
signal \ALU.un9_addsub_cry_3_c_RNI4L7ROZ0\ : std_logic;
signal \ALU.d_RNIMA3938Z0Z_4\ : std_logic;
signal \ALU.bZ0Z_4\ : std_logic;
signal \ALU.un9_addsub_cry_4_c_RNIUEDLMZ0\ : std_logic;
signal \ALU.d_RNIH1NE6FZ0Z_5\ : std_logic;
signal \ALU.bZ0Z_5\ : std_logic;
signal \ALU.d_RNILPR7TQZ0Z_6\ : std_logic;
signal \ALU.un9_addsub_cry_5_c_RNI26HCNZ0\ : std_logic;
signal \ALU.bZ0Z_6\ : std_logic;
signal \ALU.un9_addsub_cry_6_c_RNIUKMKRZ0\ : std_logic;
signal \ALU.d_RNIIIPM081Z0Z_7\ : std_logic;
signal \ALU.bZ0Z_7\ : std_logic;
signal \aluOperation_0\ : std_logic;
signal \ALU.un9_addsub_cry_7_c_RNIQIKVOZ0\ : std_logic;
signal \ALU.d_RNI7GCMD22Z0Z_8\ : std_logic;
signal \ALU.bZ0Z_8\ : std_logic;
signal \CLK_0_c_g\ : std_logic;
signal \ALU.b_cnvZ0Z_0\ : std_logic;
signal \ALU.a_15_sm0\ : std_logic;
signal \ALU.N_213_0\ : std_logic;
signal \ALU.a_15_m2_ns_1Z0Z_7\ : std_logic;
signal \ALU.aluOut_7\ : std_logic;
signal \ALU.a_15_m2_7\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \GPIO11_wire\ : std_logic;
signal \GPIO9_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \GPIO3_wire\ : std_logic;
signal \RX_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    GPIO11 <= \GPIO11_wire\;
    GPIO9 <= \GPIO9_wire\;
    TX <= \TX_wire\;
    GPIO3 <= \GPIO3_wire\;
    \RX_wire\ <= RX;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__49533\,
            GLOBALBUFFEROUTPUT => \CLK_0_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49535\,
            DIN => \N__49534\,
            DOUT => \N__49533\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49535\,
            PADOUT => \N__49534\,
            PADIN => \N__49533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO11_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49524\,
            DIN => \N__49523\,
            DOUT => \N__49522\,
            PACKAGEPIN => \GPIO11_wire\
        );

    \GPIO11_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49524\,
            PADOUT => \N__49523\,
            PADIN => \N__49522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO9_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49515\,
            DIN => \N__49514\,
            DOUT => \N__49513\,
            PACKAGEPIN => \GPIO9_wire\
        );

    \GPIO9_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49515\,
            PADOUT => \N__49514\,
            PADIN => \N__49513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32362\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TX_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49506\,
            DIN => \N__49505\,
            DOUT => \N__49504\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49506\,
            PADOUT => \N__49505\,
            PADIN => \N__49504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36485\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49497\,
            DIN => \N__49496\,
            DOUT => \N__49495\,
            PACKAGEPIN => \GPIO3_wire\
        );

    \GPIO3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49497\,
            PADOUT => \N__49496\,
            PADIN => \N__49495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15686\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RX_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49488\,
            DIN => \N__49487\,
            DOUT => \N__49486\,
            PACKAGEPIN => \RX_wire\
        );

    \RX_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49488\,
            PADOUT => \N__49487\,
            PADIN => \N__49486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12697\ : InMux
    port map (
            O => \N__49469\,
            I => \N__49464\
        );

    \I__12696\ : InMux
    port map (
            O => \N__49468\,
            I => \N__49461\
        );

    \I__12695\ : InMux
    port map (
            O => \N__49467\,
            I => \N__49457\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__49464\,
            I => \N__49454\
        );

    \I__12693\ : LocalMux
    port map (
            O => \N__49461\,
            I => \N__49451\
        );

    \I__12692\ : InMux
    port map (
            O => \N__49460\,
            I => \N__49447\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__49457\,
            I => \N__49444\
        );

    \I__12690\ : Span4Mux_h
    port map (
            O => \N__49454\,
            I => \N__49438\
        );

    \I__12689\ : Span4Mux_h
    port map (
            O => \N__49451\,
            I => \N__49435\
        );

    \I__12688\ : InMux
    port map (
            O => \N__49450\,
            I => \N__49432\
        );

    \I__12687\ : LocalMux
    port map (
            O => \N__49447\,
            I => \N__49429\
        );

    \I__12686\ : Span4Mux_v
    port map (
            O => \N__49444\,
            I => \N__49426\
        );

    \I__12685\ : InMux
    port map (
            O => \N__49443\,
            I => \N__49423\
        );

    \I__12684\ : InMux
    port map (
            O => \N__49442\,
            I => \N__49420\
        );

    \I__12683\ : InMux
    port map (
            O => \N__49441\,
            I => \N__49417\
        );

    \I__12682\ : Sp12to4
    port map (
            O => \N__49438\,
            I => \N__49410\
        );

    \I__12681\ : Sp12to4
    port map (
            O => \N__49435\,
            I => \N__49410\
        );

    \I__12680\ : LocalMux
    port map (
            O => \N__49432\,
            I => \N__49410\
        );

    \I__12679\ : Span4Mux_h
    port map (
            O => \N__49429\,
            I => \N__49407\
        );

    \I__12678\ : Span4Mux_h
    port map (
            O => \N__49426\,
            I => \N__49402\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__49423\,
            I => \N__49402\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49397\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__49417\,
            I => \N__49397\
        );

    \I__12674\ : Odrv12
    port map (
            O => \N__49410\,
            I => \ALU.un9_addsub_cry_2_c_RNIMN63NZ0\
        );

    \I__12673\ : Odrv4
    port map (
            O => \N__49407\,
            I => \ALU.un9_addsub_cry_2_c_RNIMN63NZ0\
        );

    \I__12672\ : Odrv4
    port map (
            O => \N__49402\,
            I => \ALU.un9_addsub_cry_2_c_RNIMN63NZ0\
        );

    \I__12671\ : Odrv4
    port map (
            O => \N__49397\,
            I => \ALU.un9_addsub_cry_2_c_RNIMN63NZ0\
        );

    \I__12670\ : InMux
    port map (
            O => \N__49388\,
            I => \N__49384\
        );

    \I__12669\ : InMux
    port map (
            O => \N__49387\,
            I => \N__49379\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__49384\,
            I => \N__49375\
        );

    \I__12667\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49372\
        );

    \I__12666\ : InMux
    port map (
            O => \N__49382\,
            I => \N__49369\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__49379\,
            I => \N__49365\
        );

    \I__12664\ : InMux
    port map (
            O => \N__49378\,
            I => \N__49362\
        );

    \I__12663\ : Sp12to4
    port map (
            O => \N__49375\,
            I => \N__49355\
        );

    \I__12662\ : LocalMux
    port map (
            O => \N__49372\,
            I => \N__49355\
        );

    \I__12661\ : LocalMux
    port map (
            O => \N__49369\,
            I => \N__49352\
        );

    \I__12660\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49349\
        );

    \I__12659\ : Span4Mux_h
    port map (
            O => \N__49365\,
            I => \N__49346\
        );

    \I__12658\ : LocalMux
    port map (
            O => \N__49362\,
            I => \N__49343\
        );

    \I__12657\ : InMux
    port map (
            O => \N__49361\,
            I => \N__49340\
        );

    \I__12656\ : InMux
    port map (
            O => \N__49360\,
            I => \N__49337\
        );

    \I__12655\ : Span12Mux_v
    port map (
            O => \N__49355\,
            I => \N__49334\
        );

    \I__12654\ : Span4Mux_h
    port map (
            O => \N__49352\,
            I => \N__49331\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__49349\,
            I => \N__49328\
        );

    \I__12652\ : Span4Mux_h
    port map (
            O => \N__49346\,
            I => \N__49319\
        );

    \I__12651\ : Span4Mux_v
    port map (
            O => \N__49343\,
            I => \N__49319\
        );

    \I__12650\ : LocalMux
    port map (
            O => \N__49340\,
            I => \N__49319\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49319\
        );

    \I__12648\ : Odrv12
    port map (
            O => \N__49334\,
            I => \ALU.d_RNIE8SJN5Z0Z_3\
        );

    \I__12647\ : Odrv4
    port map (
            O => \N__49331\,
            I => \ALU.d_RNIE8SJN5Z0Z_3\
        );

    \I__12646\ : Odrv4
    port map (
            O => \N__49328\,
            I => \ALU.d_RNIE8SJN5Z0Z_3\
        );

    \I__12645\ : Odrv4
    port map (
            O => \N__49319\,
            I => \ALU.d_RNIE8SJN5Z0Z_3\
        );

    \I__12644\ : InMux
    port map (
            O => \N__49310\,
            I => \N__49307\
        );

    \I__12643\ : LocalMux
    port map (
            O => \N__49307\,
            I => \N__49304\
        );

    \I__12642\ : Span4Mux_h
    port map (
            O => \N__49304\,
            I => \N__49300\
        );

    \I__12641\ : InMux
    port map (
            O => \N__49303\,
            I => \N__49297\
        );

    \I__12640\ : Span4Mux_h
    port map (
            O => \N__49300\,
            I => \N__49294\
        );

    \I__12639\ : LocalMux
    port map (
            O => \N__49297\,
            I => \ALU.bZ0Z_3\
        );

    \I__12638\ : Odrv4
    port map (
            O => \N__49294\,
            I => \ALU.bZ0Z_3\
        );

    \I__12637\ : InMux
    port map (
            O => \N__49289\,
            I => \N__49282\
        );

    \I__12636\ : InMux
    port map (
            O => \N__49288\,
            I => \N__49278\
        );

    \I__12635\ : InMux
    port map (
            O => \N__49287\,
            I => \N__49275\
        );

    \I__12634\ : InMux
    port map (
            O => \N__49286\,
            I => \N__49272\
        );

    \I__12633\ : InMux
    port map (
            O => \N__49285\,
            I => \N__49269\
        );

    \I__12632\ : LocalMux
    port map (
            O => \N__49282\,
            I => \N__49266\
        );

    \I__12631\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49263\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__49278\,
            I => \N__49259\
        );

    \I__12629\ : LocalMux
    port map (
            O => \N__49275\,
            I => \N__49248\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__49272\,
            I => \N__49248\
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__49269\,
            I => \N__49248\
        );

    \I__12626\ : Span4Mux_h
    port map (
            O => \N__49266\,
            I => \N__49248\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__49263\,
            I => \N__49248\
        );

    \I__12624\ : InMux
    port map (
            O => \N__49262\,
            I => \N__49245\
        );

    \I__12623\ : Span4Mux_h
    port map (
            O => \N__49259\,
            I => \N__49241\
        );

    \I__12622\ : Span4Mux_v
    port map (
            O => \N__49248\,
            I => \N__49236\
        );

    \I__12621\ : LocalMux
    port map (
            O => \N__49245\,
            I => \N__49236\
        );

    \I__12620\ : InMux
    port map (
            O => \N__49244\,
            I => \N__49233\
        );

    \I__12619\ : Span4Mux_v
    port map (
            O => \N__49241\,
            I => \N__49230\
        );

    \I__12618\ : Span4Mux_h
    port map (
            O => \N__49236\,
            I => \N__49225\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__49233\,
            I => \N__49225\
        );

    \I__12616\ : Odrv4
    port map (
            O => \N__49230\,
            I => \ALU.un9_addsub_cry_3_c_RNI4L7ROZ0\
        );

    \I__12615\ : Odrv4
    port map (
            O => \N__49225\,
            I => \ALU.un9_addsub_cry_3_c_RNI4L7ROZ0\
        );

    \I__12614\ : InMux
    port map (
            O => \N__49220\,
            I => \N__49214\
        );

    \I__12613\ : InMux
    port map (
            O => \N__49219\,
            I => \N__49208\
        );

    \I__12612\ : InMux
    port map (
            O => \N__49218\,
            I => \N__49205\
        );

    \I__12611\ : InMux
    port map (
            O => \N__49217\,
            I => \N__49201\
        );

    \I__12610\ : LocalMux
    port map (
            O => \N__49214\,
            I => \N__49198\
        );

    \I__12609\ : InMux
    port map (
            O => \N__49213\,
            I => \N__49195\
        );

    \I__12608\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49192\
        );

    \I__12607\ : InMux
    port map (
            O => \N__49211\,
            I => \N__49189\
        );

    \I__12606\ : LocalMux
    port map (
            O => \N__49208\,
            I => \N__49184\
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__49205\,
            I => \N__49184\
        );

    \I__12604\ : InMux
    port map (
            O => \N__49204\,
            I => \N__49181\
        );

    \I__12603\ : LocalMux
    port map (
            O => \N__49201\,
            I => \N__49178\
        );

    \I__12602\ : Span4Mux_h
    port map (
            O => \N__49198\,
            I => \N__49173\
        );

    \I__12601\ : LocalMux
    port map (
            O => \N__49195\,
            I => \N__49173\
        );

    \I__12600\ : LocalMux
    port map (
            O => \N__49192\,
            I => \N__49170\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__49189\,
            I => \N__49167\
        );

    \I__12598\ : Span4Mux_v
    port map (
            O => \N__49184\,
            I => \N__49162\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__49181\,
            I => \N__49162\
        );

    \I__12596\ : Odrv12
    port map (
            O => \N__49178\,
            I => \ALU.d_RNIMA3938Z0Z_4\
        );

    \I__12595\ : Odrv4
    port map (
            O => \N__49173\,
            I => \ALU.d_RNIMA3938Z0Z_4\
        );

    \I__12594\ : Odrv4
    port map (
            O => \N__49170\,
            I => \ALU.d_RNIMA3938Z0Z_4\
        );

    \I__12593\ : Odrv4
    port map (
            O => \N__49167\,
            I => \ALU.d_RNIMA3938Z0Z_4\
        );

    \I__12592\ : Odrv4
    port map (
            O => \N__49162\,
            I => \ALU.d_RNIMA3938Z0Z_4\
        );

    \I__12591\ : InMux
    port map (
            O => \N__49151\,
            I => \N__49148\
        );

    \I__12590\ : LocalMux
    port map (
            O => \N__49148\,
            I => \N__49145\
        );

    \I__12589\ : Span4Mux_v
    port map (
            O => \N__49145\,
            I => \N__49141\
        );

    \I__12588\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49138\
        );

    \I__12587\ : Span4Mux_h
    port map (
            O => \N__49141\,
            I => \N__49133\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__49138\,
            I => \N__49133\
        );

    \I__12585\ : Odrv4
    port map (
            O => \N__49133\,
            I => \ALU.bZ0Z_4\
        );

    \I__12584\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49127\
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__49127\,
            I => \N__49124\
        );

    \I__12582\ : Span4Mux_h
    port map (
            O => \N__49124\,
            I => \N__49119\
        );

    \I__12581\ : InMux
    port map (
            O => \N__49123\,
            I => \N__49116\
        );

    \I__12580\ : InMux
    port map (
            O => \N__49122\,
            I => \N__49113\
        );

    \I__12579\ : Span4Mux_h
    port map (
            O => \N__49119\,
            I => \N__49105\
        );

    \I__12578\ : LocalMux
    port map (
            O => \N__49116\,
            I => \N__49105\
        );

    \I__12577\ : LocalMux
    port map (
            O => \N__49113\,
            I => \N__49105\
        );

    \I__12576\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49102\
        );

    \I__12575\ : Span4Mux_v
    port map (
            O => \N__49105\,
            I => \N__49098\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__49102\,
            I => \N__49095\
        );

    \I__12573\ : InMux
    port map (
            O => \N__49101\,
            I => \N__49091\
        );

    \I__12572\ : Span4Mux_h
    port map (
            O => \N__49098\,
            I => \N__49086\
        );

    \I__12571\ : Span4Mux_v
    port map (
            O => \N__49095\,
            I => \N__49083\
        );

    \I__12570\ : InMux
    port map (
            O => \N__49094\,
            I => \N__49080\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__49091\,
            I => \N__49077\
        );

    \I__12568\ : InMux
    port map (
            O => \N__49090\,
            I => \N__49074\
        );

    \I__12567\ : InMux
    port map (
            O => \N__49089\,
            I => \N__49071\
        );

    \I__12566\ : Sp12to4
    port map (
            O => \N__49086\,
            I => \N__49068\
        );

    \I__12565\ : Span4Mux_h
    port map (
            O => \N__49083\,
            I => \N__49063\
        );

    \I__12564\ : LocalMux
    port map (
            O => \N__49080\,
            I => \N__49063\
        );

    \I__12563\ : Span4Mux_h
    port map (
            O => \N__49077\,
            I => \N__49056\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__49074\,
            I => \N__49056\
        );

    \I__12561\ : LocalMux
    port map (
            O => \N__49071\,
            I => \N__49056\
        );

    \I__12560\ : Odrv12
    port map (
            O => \N__49068\,
            I => \ALU.un9_addsub_cry_4_c_RNIUEDLMZ0\
        );

    \I__12559\ : Odrv4
    port map (
            O => \N__49063\,
            I => \ALU.un9_addsub_cry_4_c_RNIUEDLMZ0\
        );

    \I__12558\ : Odrv4
    port map (
            O => \N__49056\,
            I => \ALU.un9_addsub_cry_4_c_RNIUEDLMZ0\
        );

    \I__12557\ : InMux
    port map (
            O => \N__49049\,
            I => \N__49040\
        );

    \I__12556\ : InMux
    port map (
            O => \N__49048\,
            I => \N__49037\
        );

    \I__12555\ : InMux
    port map (
            O => \N__49047\,
            I => \N__49034\
        );

    \I__12554\ : InMux
    port map (
            O => \N__49046\,
            I => \N__49031\
        );

    \I__12553\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49028\
        );

    \I__12552\ : InMux
    port map (
            O => \N__49044\,
            I => \N__49024\
        );

    \I__12551\ : InMux
    port map (
            O => \N__49043\,
            I => \N__49021\
        );

    \I__12550\ : LocalMux
    port map (
            O => \N__49040\,
            I => \N__49018\
        );

    \I__12549\ : LocalMux
    port map (
            O => \N__49037\,
            I => \N__49013\
        );

    \I__12548\ : LocalMux
    port map (
            O => \N__49034\,
            I => \N__49013\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__49031\,
            I => \N__49010\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__49028\,
            I => \N__49007\
        );

    \I__12545\ : InMux
    port map (
            O => \N__49027\,
            I => \N__49004\
        );

    \I__12544\ : LocalMux
    port map (
            O => \N__49024\,
            I => \N__48999\
        );

    \I__12543\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__48999\
        );

    \I__12542\ : Span4Mux_v
    port map (
            O => \N__49018\,
            I => \N__48996\
        );

    \I__12541\ : Span4Mux_v
    port map (
            O => \N__49013\,
            I => \N__48991\
        );

    \I__12540\ : Span4Mux_h
    port map (
            O => \N__49010\,
            I => \N__48991\
        );

    \I__12539\ : Span4Mux_v
    port map (
            O => \N__49007\,
            I => \N__48986\
        );

    \I__12538\ : LocalMux
    port map (
            O => \N__49004\,
            I => \N__48986\
        );

    \I__12537\ : Span4Mux_v
    port map (
            O => \N__48999\,
            I => \N__48983\
        );

    \I__12536\ : Span4Mux_h
    port map (
            O => \N__48996\,
            I => \N__48976\
        );

    \I__12535\ : Span4Mux_v
    port map (
            O => \N__48991\,
            I => \N__48976\
        );

    \I__12534\ : Span4Mux_v
    port map (
            O => \N__48986\,
            I => \N__48976\
        );

    \I__12533\ : Span4Mux_v
    port map (
            O => \N__48983\,
            I => \N__48973\
        );

    \I__12532\ : Span4Mux_v
    port map (
            O => \N__48976\,
            I => \N__48970\
        );

    \I__12531\ : Odrv4
    port map (
            O => \N__48973\,
            I => \ALU.d_RNIH1NE6FZ0Z_5\
        );

    \I__12530\ : Odrv4
    port map (
            O => \N__48970\,
            I => \ALU.d_RNIH1NE6FZ0Z_5\
        );

    \I__12529\ : InMux
    port map (
            O => \N__48965\,
            I => \N__48961\
        );

    \I__12528\ : InMux
    port map (
            O => \N__48964\,
            I => \N__48958\
        );

    \I__12527\ : LocalMux
    port map (
            O => \N__48961\,
            I => \N__48955\
        );

    \I__12526\ : LocalMux
    port map (
            O => \N__48958\,
            I => \N__48950\
        );

    \I__12525\ : Span4Mux_h
    port map (
            O => \N__48955\,
            I => \N__48950\
        );

    \I__12524\ : Odrv4
    port map (
            O => \N__48950\,
            I => \ALU.bZ0Z_5\
        );

    \I__12523\ : InMux
    port map (
            O => \N__48947\,
            I => \N__48944\
        );

    \I__12522\ : LocalMux
    port map (
            O => \N__48944\,
            I => \N__48939\
        );

    \I__12521\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48936\
        );

    \I__12520\ : InMux
    port map (
            O => \N__48942\,
            I => \N__48933\
        );

    \I__12519\ : Span4Mux_v
    port map (
            O => \N__48939\,
            I => \N__48924\
        );

    \I__12518\ : LocalMux
    port map (
            O => \N__48936\,
            I => \N__48924\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__48933\,
            I => \N__48924\
        );

    \I__12516\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48921\
        );

    \I__12515\ : InMux
    port map (
            O => \N__48931\,
            I => \N__48918\
        );

    \I__12514\ : Span4Mux_v
    port map (
            O => \N__48924\,
            I => \N__48909\
        );

    \I__12513\ : LocalMux
    port map (
            O => \N__48921\,
            I => \N__48909\
        );

    \I__12512\ : LocalMux
    port map (
            O => \N__48918\,
            I => \N__48909\
        );

    \I__12511\ : InMux
    port map (
            O => \N__48917\,
            I => \N__48906\
        );

    \I__12510\ : InMux
    port map (
            O => \N__48916\,
            I => \N__48903\
        );

    \I__12509\ : Span4Mux_h
    port map (
            O => \N__48909\,
            I => \N__48896\
        );

    \I__12508\ : LocalMux
    port map (
            O => \N__48906\,
            I => \N__48896\
        );

    \I__12507\ : LocalMux
    port map (
            O => \N__48903\,
            I => \N__48896\
        );

    \I__12506\ : Odrv4
    port map (
            O => \N__48896\,
            I => \ALU.d_RNILPR7TQZ0Z_6\
        );

    \I__12505\ : InMux
    port map (
            O => \N__48893\,
            I => \N__48888\
        );

    \I__12504\ : InMux
    port map (
            O => \N__48892\,
            I => \N__48885\
        );

    \I__12503\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48882\
        );

    \I__12502\ : LocalMux
    port map (
            O => \N__48888\,
            I => \N__48877\
        );

    \I__12501\ : LocalMux
    port map (
            O => \N__48885\,
            I => \N__48874\
        );

    \I__12500\ : LocalMux
    port map (
            O => \N__48882\,
            I => \N__48871\
        );

    \I__12499\ : InMux
    port map (
            O => \N__48881\,
            I => \N__48868\
        );

    \I__12498\ : InMux
    port map (
            O => \N__48880\,
            I => \N__48864\
        );

    \I__12497\ : Span4Mux_h
    port map (
            O => \N__48877\,
            I => \N__48860\
        );

    \I__12496\ : Span4Mux_h
    port map (
            O => \N__48874\,
            I => \N__48857\
        );

    \I__12495\ : Span4Mux_v
    port map (
            O => \N__48871\,
            I => \N__48851\
        );

    \I__12494\ : LocalMux
    port map (
            O => \N__48868\,
            I => \N__48851\
        );

    \I__12493\ : InMux
    port map (
            O => \N__48867\,
            I => \N__48848\
        );

    \I__12492\ : LocalMux
    port map (
            O => \N__48864\,
            I => \N__48845\
        );

    \I__12491\ : InMux
    port map (
            O => \N__48863\,
            I => \N__48842\
        );

    \I__12490\ : Span4Mux_v
    port map (
            O => \N__48860\,
            I => \N__48839\
        );

    \I__12489\ : Span4Mux_v
    port map (
            O => \N__48857\,
            I => \N__48836\
        );

    \I__12488\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48833\
        );

    \I__12487\ : Span4Mux_h
    port map (
            O => \N__48851\,
            I => \N__48824\
        );

    \I__12486\ : LocalMux
    port map (
            O => \N__48848\,
            I => \N__48824\
        );

    \I__12485\ : Span4Mux_h
    port map (
            O => \N__48845\,
            I => \N__48824\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__48842\,
            I => \N__48824\
        );

    \I__12483\ : Odrv4
    port map (
            O => \N__48839\,
            I => \ALU.un9_addsub_cry_5_c_RNI26HCNZ0\
        );

    \I__12482\ : Odrv4
    port map (
            O => \N__48836\,
            I => \ALU.un9_addsub_cry_5_c_RNI26HCNZ0\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__48833\,
            I => \ALU.un9_addsub_cry_5_c_RNI26HCNZ0\
        );

    \I__12480\ : Odrv4
    port map (
            O => \N__48824\,
            I => \ALU.un9_addsub_cry_5_c_RNI26HCNZ0\
        );

    \I__12479\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48812\
        );

    \I__12478\ : LocalMux
    port map (
            O => \N__48812\,
            I => \N__48808\
        );

    \I__12477\ : InMux
    port map (
            O => \N__48811\,
            I => \N__48805\
        );

    \I__12476\ : Span4Mux_h
    port map (
            O => \N__48808\,
            I => \N__48802\
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__48805\,
            I => \N__48799\
        );

    \I__12474\ : Span4Mux_h
    port map (
            O => \N__48802\,
            I => \N__48796\
        );

    \I__12473\ : Odrv12
    port map (
            O => \N__48799\,
            I => \ALU.bZ0Z_6\
        );

    \I__12472\ : Odrv4
    port map (
            O => \N__48796\,
            I => \ALU.bZ0Z_6\
        );

    \I__12471\ : InMux
    port map (
            O => \N__48791\,
            I => \N__48784\
        );

    \I__12470\ : InMux
    port map (
            O => \N__48790\,
            I => \N__48781\
        );

    \I__12469\ : InMux
    port map (
            O => \N__48789\,
            I => \N__48778\
        );

    \I__12468\ : InMux
    port map (
            O => \N__48788\,
            I => \N__48774\
        );

    \I__12467\ : InMux
    port map (
            O => \N__48787\,
            I => \N__48771\
        );

    \I__12466\ : LocalMux
    port map (
            O => \N__48784\,
            I => \N__48765\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48765\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__48778\,
            I => \N__48762\
        );

    \I__12463\ : InMux
    port map (
            O => \N__48777\,
            I => \N__48759\
        );

    \I__12462\ : LocalMux
    port map (
            O => \N__48774\,
            I => \N__48756\
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__48771\,
            I => \N__48753\
        );

    \I__12460\ : InMux
    port map (
            O => \N__48770\,
            I => \N__48750\
        );

    \I__12459\ : Span4Mux_h
    port map (
            O => \N__48765\,
            I => \N__48742\
        );

    \I__12458\ : Span4Mux_h
    port map (
            O => \N__48762\,
            I => \N__48742\
        );

    \I__12457\ : LocalMux
    port map (
            O => \N__48759\,
            I => \N__48742\
        );

    \I__12456\ : Span4Mux_v
    port map (
            O => \N__48756\,
            I => \N__48735\
        );

    \I__12455\ : Span4Mux_v
    port map (
            O => \N__48753\,
            I => \N__48735\
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__48750\,
            I => \N__48735\
        );

    \I__12453\ : InMux
    port map (
            O => \N__48749\,
            I => \N__48732\
        );

    \I__12452\ : Span4Mux_h
    port map (
            O => \N__48742\,
            I => \N__48729\
        );

    \I__12451\ : Span4Mux_h
    port map (
            O => \N__48735\,
            I => \N__48726\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__48732\,
            I => \N__48723\
        );

    \I__12449\ : Odrv4
    port map (
            O => \N__48729\,
            I => \ALU.un9_addsub_cry_6_c_RNIUKMKRZ0\
        );

    \I__12448\ : Odrv4
    port map (
            O => \N__48726\,
            I => \ALU.un9_addsub_cry_6_c_RNIUKMKRZ0\
        );

    \I__12447\ : Odrv12
    port map (
            O => \N__48723\,
            I => \ALU.un9_addsub_cry_6_c_RNIUKMKRZ0\
        );

    \I__12446\ : InMux
    port map (
            O => \N__48716\,
            I => \N__48710\
        );

    \I__12445\ : InMux
    port map (
            O => \N__48715\,
            I => \N__48707\
        );

    \I__12444\ : InMux
    port map (
            O => \N__48714\,
            I => \N__48704\
        );

    \I__12443\ : InMux
    port map (
            O => \N__48713\,
            I => \N__48701\
        );

    \I__12442\ : LocalMux
    port map (
            O => \N__48710\,
            I => \N__48697\
        );

    \I__12441\ : LocalMux
    port map (
            O => \N__48707\,
            I => \N__48688\
        );

    \I__12440\ : LocalMux
    port map (
            O => \N__48704\,
            I => \N__48688\
        );

    \I__12439\ : LocalMux
    port map (
            O => \N__48701\,
            I => \N__48688\
        );

    \I__12438\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48685\
        );

    \I__12437\ : Span4Mux_h
    port map (
            O => \N__48697\,
            I => \N__48681\
        );

    \I__12436\ : InMux
    port map (
            O => \N__48696\,
            I => \N__48678\
        );

    \I__12435\ : InMux
    port map (
            O => \N__48695\,
            I => \N__48675\
        );

    \I__12434\ : Span4Mux_v
    port map (
            O => \N__48688\,
            I => \N__48670\
        );

    \I__12433\ : LocalMux
    port map (
            O => \N__48685\,
            I => \N__48670\
        );

    \I__12432\ : InMux
    port map (
            O => \N__48684\,
            I => \N__48667\
        );

    \I__12431\ : Odrv4
    port map (
            O => \N__48681\,
            I => \ALU.d_RNIIIPM081Z0Z_7\
        );

    \I__12430\ : LocalMux
    port map (
            O => \N__48678\,
            I => \ALU.d_RNIIIPM081Z0Z_7\
        );

    \I__12429\ : LocalMux
    port map (
            O => \N__48675\,
            I => \ALU.d_RNIIIPM081Z0Z_7\
        );

    \I__12428\ : Odrv4
    port map (
            O => \N__48670\,
            I => \ALU.d_RNIIIPM081Z0Z_7\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__48667\,
            I => \ALU.d_RNIIIPM081Z0Z_7\
        );

    \I__12426\ : InMux
    port map (
            O => \N__48656\,
            I => \N__48650\
        );

    \I__12425\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48650\
        );

    \I__12424\ : LocalMux
    port map (
            O => \N__48650\,
            I => \N__48647\
        );

    \I__12423\ : Span4Mux_h
    port map (
            O => \N__48647\,
            I => \N__48644\
        );

    \I__12422\ : Odrv4
    port map (
            O => \N__48644\,
            I => \ALU.bZ0Z_7\
        );

    \I__12421\ : InMux
    port map (
            O => \N__48641\,
            I => \N__48606\
        );

    \I__12420\ : InMux
    port map (
            O => \N__48640\,
            I => \N__48606\
        );

    \I__12419\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48606\
        );

    \I__12418\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48606\
        );

    \I__12417\ : InMux
    port map (
            O => \N__48637\,
            I => \N__48599\
        );

    \I__12416\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48599\
        );

    \I__12415\ : InMux
    port map (
            O => \N__48635\,
            I => \N__48599\
        );

    \I__12414\ : CascadeMux
    port map (
            O => \N__48634\,
            I => \N__48557\
        );

    \I__12413\ : InMux
    port map (
            O => \N__48633\,
            I => \N__48548\
        );

    \I__12412\ : InMux
    port map (
            O => \N__48632\,
            I => \N__48548\
        );

    \I__12411\ : InMux
    port map (
            O => \N__48631\,
            I => \N__48548\
        );

    \I__12410\ : InMux
    port map (
            O => \N__48630\,
            I => \N__48545\
        );

    \I__12409\ : InMux
    port map (
            O => \N__48629\,
            I => \N__48542\
        );

    \I__12408\ : InMux
    port map (
            O => \N__48628\,
            I => \N__48535\
        );

    \I__12407\ : InMux
    port map (
            O => \N__48627\,
            I => \N__48535\
        );

    \I__12406\ : InMux
    port map (
            O => \N__48626\,
            I => \N__48535\
        );

    \I__12405\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48526\
        );

    \I__12404\ : InMux
    port map (
            O => \N__48624\,
            I => \N__48526\
        );

    \I__12403\ : InMux
    port map (
            O => \N__48623\,
            I => \N__48526\
        );

    \I__12402\ : InMux
    port map (
            O => \N__48622\,
            I => \N__48526\
        );

    \I__12401\ : InMux
    port map (
            O => \N__48621\,
            I => \N__48517\
        );

    \I__12400\ : InMux
    port map (
            O => \N__48620\,
            I => \N__48517\
        );

    \I__12399\ : InMux
    port map (
            O => \N__48619\,
            I => \N__48517\
        );

    \I__12398\ : InMux
    port map (
            O => \N__48618\,
            I => \N__48517\
        );

    \I__12397\ : InMux
    port map (
            O => \N__48617\,
            I => \N__48510\
        );

    \I__12396\ : InMux
    port map (
            O => \N__48616\,
            I => \N__48510\
        );

    \I__12395\ : InMux
    port map (
            O => \N__48615\,
            I => \N__48510\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__48606\,
            I => \N__48504\
        );

    \I__12393\ : LocalMux
    port map (
            O => \N__48599\,
            I => \N__48504\
        );

    \I__12392\ : InMux
    port map (
            O => \N__48598\,
            I => \N__48501\
        );

    \I__12391\ : InMux
    port map (
            O => \N__48597\,
            I => \N__48498\
        );

    \I__12390\ : InMux
    port map (
            O => \N__48596\,
            I => \N__48472\
        );

    \I__12389\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48472\
        );

    \I__12388\ : InMux
    port map (
            O => \N__48594\,
            I => \N__48472\
        );

    \I__12387\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48472\
        );

    \I__12386\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48472\
        );

    \I__12385\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48469\
        );

    \I__12384\ : InMux
    port map (
            O => \N__48590\,
            I => \N__48464\
        );

    \I__12383\ : InMux
    port map (
            O => \N__48589\,
            I => \N__48464\
        );

    \I__12382\ : InMux
    port map (
            O => \N__48588\,
            I => \N__48461\
        );

    \I__12381\ : InMux
    port map (
            O => \N__48587\,
            I => \N__48454\
        );

    \I__12380\ : InMux
    port map (
            O => \N__48586\,
            I => \N__48454\
        );

    \I__12379\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48454\
        );

    \I__12378\ : InMux
    port map (
            O => \N__48584\,
            I => \N__48447\
        );

    \I__12377\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48447\
        );

    \I__12376\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48447\
        );

    \I__12375\ : InMux
    port map (
            O => \N__48581\,
            I => \N__48444\
        );

    \I__12374\ : InMux
    port map (
            O => \N__48580\,
            I => \N__48437\
        );

    \I__12373\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48437\
        );

    \I__12372\ : InMux
    port map (
            O => \N__48578\,
            I => \N__48437\
        );

    \I__12371\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48427\
        );

    \I__12370\ : CascadeMux
    port map (
            O => \N__48576\,
            I => \N__48416\
        );

    \I__12369\ : CascadeMux
    port map (
            O => \N__48575\,
            I => \N__48413\
        );

    \I__12368\ : InMux
    port map (
            O => \N__48574\,
            I => \N__48406\
        );

    \I__12367\ : InMux
    port map (
            O => \N__48573\,
            I => \N__48401\
        );

    \I__12366\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48401\
        );

    \I__12365\ : InMux
    port map (
            O => \N__48571\,
            I => \N__48396\
        );

    \I__12364\ : InMux
    port map (
            O => \N__48570\,
            I => \N__48396\
        );

    \I__12363\ : InMux
    port map (
            O => \N__48569\,
            I => \N__48389\
        );

    \I__12362\ : InMux
    port map (
            O => \N__48568\,
            I => \N__48389\
        );

    \I__12361\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48389\
        );

    \I__12360\ : InMux
    port map (
            O => \N__48566\,
            I => \N__48384\
        );

    \I__12359\ : InMux
    port map (
            O => \N__48565\,
            I => \N__48384\
        );

    \I__12358\ : InMux
    port map (
            O => \N__48564\,
            I => \N__48375\
        );

    \I__12357\ : InMux
    port map (
            O => \N__48563\,
            I => \N__48375\
        );

    \I__12356\ : InMux
    port map (
            O => \N__48562\,
            I => \N__48375\
        );

    \I__12355\ : InMux
    port map (
            O => \N__48561\,
            I => \N__48375\
        );

    \I__12354\ : InMux
    port map (
            O => \N__48560\,
            I => \N__48366\
        );

    \I__12353\ : InMux
    port map (
            O => \N__48557\,
            I => \N__48366\
        );

    \I__12352\ : InMux
    port map (
            O => \N__48556\,
            I => \N__48366\
        );

    \I__12351\ : InMux
    port map (
            O => \N__48555\,
            I => \N__48366\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__48548\,
            I => \N__48363\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__48545\,
            I => \N__48354\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__48542\,
            I => \N__48354\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__48535\,
            I => \N__48354\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__48526\,
            I => \N__48354\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48349\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__48510\,
            I => \N__48349\
        );

    \I__12343\ : InMux
    port map (
            O => \N__48509\,
            I => \N__48341\
        );

    \I__12342\ : Span4Mux_h
    port map (
            O => \N__48504\,
            I => \N__48334\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__48501\,
            I => \N__48334\
        );

    \I__12340\ : LocalMux
    port map (
            O => \N__48498\,
            I => \N__48331\
        );

    \I__12339\ : InMux
    port map (
            O => \N__48497\,
            I => \N__48317\
        );

    \I__12338\ : InMux
    port map (
            O => \N__48496\,
            I => \N__48317\
        );

    \I__12337\ : InMux
    port map (
            O => \N__48495\,
            I => \N__48317\
        );

    \I__12336\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48317\
        );

    \I__12335\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48317\
        );

    \I__12334\ : InMux
    port map (
            O => \N__48492\,
            I => \N__48310\
        );

    \I__12333\ : InMux
    port map (
            O => \N__48491\,
            I => \N__48310\
        );

    \I__12332\ : InMux
    port map (
            O => \N__48490\,
            I => \N__48310\
        );

    \I__12331\ : InMux
    port map (
            O => \N__48489\,
            I => \N__48301\
        );

    \I__12330\ : InMux
    port map (
            O => \N__48488\,
            I => \N__48301\
        );

    \I__12329\ : InMux
    port map (
            O => \N__48487\,
            I => \N__48301\
        );

    \I__12328\ : InMux
    port map (
            O => \N__48486\,
            I => \N__48301\
        );

    \I__12327\ : InMux
    port map (
            O => \N__48485\,
            I => \N__48294\
        );

    \I__12326\ : InMux
    port map (
            O => \N__48484\,
            I => \N__48294\
        );

    \I__12325\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48294\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__48472\,
            I => \N__48291\
        );

    \I__12323\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48284\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48284\
        );

    \I__12321\ : LocalMux
    port map (
            O => \N__48461\,
            I => \N__48284\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__48454\,
            I => \N__48275\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__48447\,
            I => \N__48275\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__48444\,
            I => \N__48275\
        );

    \I__12317\ : LocalMux
    port map (
            O => \N__48437\,
            I => \N__48275\
        );

    \I__12316\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48262\
        );

    \I__12315\ : InMux
    port map (
            O => \N__48435\,
            I => \N__48258\
        );

    \I__12314\ : InMux
    port map (
            O => \N__48434\,
            I => \N__48255\
        );

    \I__12313\ : InMux
    port map (
            O => \N__48433\,
            I => \N__48252\
        );

    \I__12312\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48244\
        );

    \I__12311\ : InMux
    port map (
            O => \N__48431\,
            I => \N__48244\
        );

    \I__12310\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48244\
        );

    \I__12309\ : LocalMux
    port map (
            O => \N__48427\,
            I => \N__48241\
        );

    \I__12308\ : InMux
    port map (
            O => \N__48426\,
            I => \N__48238\
        );

    \I__12307\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48227\
        );

    \I__12306\ : InMux
    port map (
            O => \N__48424\,
            I => \N__48227\
        );

    \I__12305\ : InMux
    port map (
            O => \N__48423\,
            I => \N__48227\
        );

    \I__12304\ : InMux
    port map (
            O => \N__48422\,
            I => \N__48227\
        );

    \I__12303\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48227\
        );

    \I__12302\ : InMux
    port map (
            O => \N__48420\,
            I => \N__48222\
        );

    \I__12301\ : InMux
    port map (
            O => \N__48419\,
            I => \N__48222\
        );

    \I__12300\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48215\
        );

    \I__12299\ : InMux
    port map (
            O => \N__48413\,
            I => \N__48215\
        );

    \I__12298\ : InMux
    port map (
            O => \N__48412\,
            I => \N__48215\
        );

    \I__12297\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48208\
        );

    \I__12296\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48208\
        );

    \I__12295\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48208\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__48406\,
            I => \N__48203\
        );

    \I__12293\ : LocalMux
    port map (
            O => \N__48401\,
            I => \N__48203\
        );

    \I__12292\ : LocalMux
    port map (
            O => \N__48396\,
            I => \N__48186\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__48389\,
            I => \N__48186\
        );

    \I__12290\ : LocalMux
    port map (
            O => \N__48384\,
            I => \N__48186\
        );

    \I__12289\ : LocalMux
    port map (
            O => \N__48375\,
            I => \N__48186\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__48366\,
            I => \N__48186\
        );

    \I__12287\ : Span4Mux_v
    port map (
            O => \N__48363\,
            I => \N__48186\
        );

    \I__12286\ : Span4Mux_v
    port map (
            O => \N__48354\,
            I => \N__48186\
        );

    \I__12285\ : Span4Mux_h
    port map (
            O => \N__48349\,
            I => \N__48186\
        );

    \I__12284\ : InMux
    port map (
            O => \N__48348\,
            I => \N__48183\
        );

    \I__12283\ : InMux
    port map (
            O => \N__48347\,
            I => \N__48174\
        );

    \I__12282\ : InMux
    port map (
            O => \N__48346\,
            I => \N__48174\
        );

    \I__12281\ : InMux
    port map (
            O => \N__48345\,
            I => \N__48174\
        );

    \I__12280\ : InMux
    port map (
            O => \N__48344\,
            I => \N__48174\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__48341\,
            I => \N__48171\
        );

    \I__12278\ : InMux
    port map (
            O => \N__48340\,
            I => \N__48166\
        );

    \I__12277\ : InMux
    port map (
            O => \N__48339\,
            I => \N__48166\
        );

    \I__12276\ : Span4Mux_h
    port map (
            O => \N__48334\,
            I => \N__48161\
        );

    \I__12275\ : Span4Mux_v
    port map (
            O => \N__48331\,
            I => \N__48161\
        );

    \I__12274\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48156\
        );

    \I__12273\ : InMux
    port map (
            O => \N__48329\,
            I => \N__48156\
        );

    \I__12272\ : InMux
    port map (
            O => \N__48328\,
            I => \N__48153\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__48317\,
            I => \N__48146\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__48310\,
            I => \N__48146\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__48301\,
            I => \N__48146\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__48294\,
            I => \N__48137\
        );

    \I__12267\ : Span4Mux_h
    port map (
            O => \N__48291\,
            I => \N__48137\
        );

    \I__12266\ : Span4Mux_v
    port map (
            O => \N__48284\,
            I => \N__48137\
        );

    \I__12265\ : Span4Mux_h
    port map (
            O => \N__48275\,
            I => \N__48137\
        );

    \I__12264\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48132\
        );

    \I__12263\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48132\
        );

    \I__12262\ : InMux
    port map (
            O => \N__48272\,
            I => \N__48127\
        );

    \I__12261\ : InMux
    port map (
            O => \N__48271\,
            I => \N__48127\
        );

    \I__12260\ : InMux
    port map (
            O => \N__48270\,
            I => \N__48122\
        );

    \I__12259\ : InMux
    port map (
            O => \N__48269\,
            I => \N__48122\
        );

    \I__12258\ : InMux
    port map (
            O => \N__48268\,
            I => \N__48113\
        );

    \I__12257\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48113\
        );

    \I__12256\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48113\
        );

    \I__12255\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48113\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__48262\,
            I => \N__48110\
        );

    \I__12253\ : InMux
    port map (
            O => \N__48261\,
            I => \N__48106\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__48258\,
            I => \N__48100\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__48255\,
            I => \N__48100\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__48252\,
            I => \N__48097\
        );

    \I__12249\ : InMux
    port map (
            O => \N__48251\,
            I => \N__48089\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__48244\,
            I => \N__48078\
        );

    \I__12247\ : Span4Mux_h
    port map (
            O => \N__48241\,
            I => \N__48078\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__48238\,
            I => \N__48078\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__48227\,
            I => \N__48078\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__48222\,
            I => \N__48078\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__48215\,
            I => \N__48065\
        );

    \I__12242\ : LocalMux
    port map (
            O => \N__48208\,
            I => \N__48065\
        );

    \I__12241\ : Span4Mux_v
    port map (
            O => \N__48203\,
            I => \N__48065\
        );

    \I__12240\ : Span4Mux_v
    port map (
            O => \N__48186\,
            I => \N__48065\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__48183\,
            I => \N__48060\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__48174\,
            I => \N__48060\
        );

    \I__12237\ : Span4Mux_h
    port map (
            O => \N__48171\,
            I => \N__48055\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__48166\,
            I => \N__48055\
        );

    \I__12235\ : Span4Mux_v
    port map (
            O => \N__48161\,
            I => \N__48049\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__48156\,
            I => \N__48049\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__48153\,
            I => \N__48034\
        );

    \I__12232\ : Span4Mux_v
    port map (
            O => \N__48146\,
            I => \N__48034\
        );

    \I__12231\ : Span4Mux_v
    port map (
            O => \N__48137\,
            I => \N__48034\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__48132\,
            I => \N__48034\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__48127\,
            I => \N__48034\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__48122\,
            I => \N__48034\
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__48113\,
            I => \N__48034\
        );

    \I__12226\ : Span4Mux_h
    port map (
            O => \N__48110\,
            I => \N__48031\
        );

    \I__12225\ : InMux
    port map (
            O => \N__48109\,
            I => \N__48026\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__48106\,
            I => \N__48023\
        );

    \I__12223\ : InMux
    port map (
            O => \N__48105\,
            I => \N__48020\
        );

    \I__12222\ : Span4Mux_v
    port map (
            O => \N__48100\,
            I => \N__48017\
        );

    \I__12221\ : Span4Mux_h
    port map (
            O => \N__48097\,
            I => \N__48014\
        );

    \I__12220\ : InMux
    port map (
            O => \N__48096\,
            I => \N__48007\
        );

    \I__12219\ : InMux
    port map (
            O => \N__48095\,
            I => \N__48007\
        );

    \I__12218\ : InMux
    port map (
            O => \N__48094\,
            I => \N__48007\
        );

    \I__12217\ : InMux
    port map (
            O => \N__48093\,
            I => \N__48002\
        );

    \I__12216\ : InMux
    port map (
            O => \N__48092\,
            I => \N__48002\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__48089\,
            I => \N__47997\
        );

    \I__12214\ : Span4Mux_v
    port map (
            O => \N__48078\,
            I => \N__47997\
        );

    \I__12213\ : InMux
    port map (
            O => \N__48077\,
            I => \N__47990\
        );

    \I__12212\ : InMux
    port map (
            O => \N__48076\,
            I => \N__47990\
        );

    \I__12211\ : InMux
    port map (
            O => \N__48075\,
            I => \N__47990\
        );

    \I__12210\ : InMux
    port map (
            O => \N__48074\,
            I => \N__47987\
        );

    \I__12209\ : Span4Mux_v
    port map (
            O => \N__48065\,
            I => \N__47984\
        );

    \I__12208\ : Span4Mux_v
    port map (
            O => \N__48060\,
            I => \N__47979\
        );

    \I__12207\ : Span4Mux_v
    port map (
            O => \N__48055\,
            I => \N__47979\
        );

    \I__12206\ : CascadeMux
    port map (
            O => \N__48054\,
            I => \N__47976\
        );

    \I__12205\ : Span4Mux_v
    port map (
            O => \N__48049\,
            I => \N__47971\
        );

    \I__12204\ : Span4Mux_v
    port map (
            O => \N__48034\,
            I => \N__47971\
        );

    \I__12203\ : Span4Mux_h
    port map (
            O => \N__48031\,
            I => \N__47968\
        );

    \I__12202\ : InMux
    port map (
            O => \N__48030\,
            I => \N__47963\
        );

    \I__12201\ : InMux
    port map (
            O => \N__48029\,
            I => \N__47963\
        );

    \I__12200\ : LocalMux
    port map (
            O => \N__48026\,
            I => \N__47958\
        );

    \I__12199\ : Span4Mux_s1_h
    port map (
            O => \N__48023\,
            I => \N__47958\
        );

    \I__12198\ : LocalMux
    port map (
            O => \N__48020\,
            I => \N__47953\
        );

    \I__12197\ : Span4Mux_v
    port map (
            O => \N__48017\,
            I => \N__47953\
        );

    \I__12196\ : Sp12to4
    port map (
            O => \N__48014\,
            I => \N__47950\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__48007\,
            I => \N__47941\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__48002\,
            I => \N__47941\
        );

    \I__12193\ : Sp12to4
    port map (
            O => \N__47997\,
            I => \N__47941\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__47990\,
            I => \N__47941\
        );

    \I__12191\ : LocalMux
    port map (
            O => \N__47987\,
            I => \N__47934\
        );

    \I__12190\ : Span4Mux_v
    port map (
            O => \N__47984\,
            I => \N__47934\
        );

    \I__12189\ : Span4Mux_v
    port map (
            O => \N__47979\,
            I => \N__47934\
        );

    \I__12188\ : InMux
    port map (
            O => \N__47976\,
            I => \N__47931\
        );

    \I__12187\ : Span4Mux_h
    port map (
            O => \N__47971\,
            I => \N__47928\
        );

    \I__12186\ : Span4Mux_v
    port map (
            O => \N__47968\,
            I => \N__47925\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__47963\,
            I => \N__47918\
        );

    \I__12184\ : Span4Mux_v
    port map (
            O => \N__47958\,
            I => \N__47918\
        );

    \I__12183\ : Span4Mux_h
    port map (
            O => \N__47953\,
            I => \N__47918\
        );

    \I__12182\ : Span12Mux_v
    port map (
            O => \N__47950\,
            I => \N__47913\
        );

    \I__12181\ : Span12Mux_h
    port map (
            O => \N__47941\,
            I => \N__47913\
        );

    \I__12180\ : Span4Mux_h
    port map (
            O => \N__47934\,
            I => \N__47908\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__47931\,
            I => \N__47908\
        );

    \I__12178\ : Span4Mux_h
    port map (
            O => \N__47928\,
            I => \N__47905\
        );

    \I__12177\ : Odrv4
    port map (
            O => \N__47925\,
            I => \aluOperation_0\
        );

    \I__12176\ : Odrv4
    port map (
            O => \N__47918\,
            I => \aluOperation_0\
        );

    \I__12175\ : Odrv12
    port map (
            O => \N__47913\,
            I => \aluOperation_0\
        );

    \I__12174\ : Odrv4
    port map (
            O => \N__47908\,
            I => \aluOperation_0\
        );

    \I__12173\ : Odrv4
    port map (
            O => \N__47905\,
            I => \aluOperation_0\
        );

    \I__12172\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47889\
        );

    \I__12171\ : InMux
    port map (
            O => \N__47893\,
            I => \N__47883\
        );

    \I__12170\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47880\
        );

    \I__12169\ : LocalMux
    port map (
            O => \N__47889\,
            I => \N__47877\
        );

    \I__12168\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47874\
        );

    \I__12167\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47871\
        );

    \I__12166\ : InMux
    port map (
            O => \N__47886\,
            I => \N__47868\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__47883\,
            I => \N__47865\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__47880\,
            I => \N__47861\
        );

    \I__12163\ : Span4Mux_h
    port map (
            O => \N__47877\,
            I => \N__47858\
        );

    \I__12162\ : LocalMux
    port map (
            O => \N__47874\,
            I => \N__47853\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__47871\,
            I => \N__47853\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__47868\,
            I => \N__47850\
        );

    \I__12159\ : Span4Mux_v
    port map (
            O => \N__47865\,
            I => \N__47847\
        );

    \I__12158\ : InMux
    port map (
            O => \N__47864\,
            I => \N__47844\
        );

    \I__12157\ : Span4Mux_v
    port map (
            O => \N__47861\,
            I => \N__47841\
        );

    \I__12156\ : Span4Mux_h
    port map (
            O => \N__47858\,
            I => \N__47836\
        );

    \I__12155\ : Span4Mux_s2_v
    port map (
            O => \N__47853\,
            I => \N__47836\
        );

    \I__12154\ : Span4Mux_v
    port map (
            O => \N__47850\,
            I => \N__47833\
        );

    \I__12153\ : Span4Mux_h
    port map (
            O => \N__47847\,
            I => \N__47828\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__47844\,
            I => \N__47828\
        );

    \I__12151\ : Span4Mux_v
    port map (
            O => \N__47841\,
            I => \N__47818\
        );

    \I__12150\ : Span4Mux_v
    port map (
            O => \N__47836\,
            I => \N__47818\
        );

    \I__12149\ : Span4Mux_v
    port map (
            O => \N__47833\,
            I => \N__47818\
        );

    \I__12148\ : Span4Mux_h
    port map (
            O => \N__47828\,
            I => \N__47818\
        );

    \I__12147\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47815\
        );

    \I__12146\ : Odrv4
    port map (
            O => \N__47818\,
            I => \ALU.un9_addsub_cry_7_c_RNIQIKVOZ0\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__47815\,
            I => \ALU.un9_addsub_cry_7_c_RNIQIKVOZ0\
        );

    \I__12144\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47805\
        );

    \I__12143\ : InMux
    port map (
            O => \N__47809\,
            I => \N__47802\
        );

    \I__12142\ : InMux
    port map (
            O => \N__47808\,
            I => \N__47799\
        );

    \I__12141\ : LocalMux
    port map (
            O => \N__47805\,
            I => \N__47795\
        );

    \I__12140\ : LocalMux
    port map (
            O => \N__47802\,
            I => \N__47791\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__47799\,
            I => \N__47788\
        );

    \I__12138\ : InMux
    port map (
            O => \N__47798\,
            I => \N__47785\
        );

    \I__12137\ : Span4Mux_v
    port map (
            O => \N__47795\,
            I => \N__47782\
        );

    \I__12136\ : InMux
    port map (
            O => \N__47794\,
            I => \N__47779\
        );

    \I__12135\ : Span4Mux_h
    port map (
            O => \N__47791\,
            I => \N__47774\
        );

    \I__12134\ : Span4Mux_h
    port map (
            O => \N__47788\,
            I => \N__47771\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__47785\,
            I => \N__47768\
        );

    \I__12132\ : Span4Mux_h
    port map (
            O => \N__47782\,
            I => \N__47763\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__47779\,
            I => \N__47763\
        );

    \I__12130\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47760\
        );

    \I__12129\ : InMux
    port map (
            O => \N__47777\,
            I => \N__47757\
        );

    \I__12128\ : Span4Mux_h
    port map (
            O => \N__47774\,
            I => \N__47753\
        );

    \I__12127\ : Span4Mux_h
    port map (
            O => \N__47771\,
            I => \N__47750\
        );

    \I__12126\ : Span4Mux_s3_v
    port map (
            O => \N__47768\,
            I => \N__47747\
        );

    \I__12125\ : Span4Mux_v
    port map (
            O => \N__47763\,
            I => \N__47744\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__47760\,
            I => \N__47741\
        );

    \I__12123\ : LocalMux
    port map (
            O => \N__47757\,
            I => \N__47738\
        );

    \I__12122\ : InMux
    port map (
            O => \N__47756\,
            I => \N__47735\
        );

    \I__12121\ : Odrv4
    port map (
            O => \N__47753\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12120\ : Odrv4
    port map (
            O => \N__47750\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12119\ : Odrv4
    port map (
            O => \N__47747\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12118\ : Odrv4
    port map (
            O => \N__47744\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12117\ : Odrv12
    port map (
            O => \N__47741\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12116\ : Odrv12
    port map (
            O => \N__47738\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__47735\,
            I => \ALU.d_RNI7GCMD22Z0Z_8\
        );

    \I__12114\ : InMux
    port map (
            O => \N__47720\,
            I => \N__47716\
        );

    \I__12113\ : InMux
    port map (
            O => \N__47719\,
            I => \N__47713\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__47716\,
            I => \N__47710\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__47713\,
            I => \N__47707\
        );

    \I__12110\ : Span4Mux_v
    port map (
            O => \N__47710\,
            I => \N__47702\
        );

    \I__12109\ : Span4Mux_v
    port map (
            O => \N__47707\,
            I => \N__47702\
        );

    \I__12108\ : Span4Mux_h
    port map (
            O => \N__47702\,
            I => \N__47699\
        );

    \I__12107\ : Span4Mux_h
    port map (
            O => \N__47699\,
            I => \N__47696\
        );

    \I__12106\ : Odrv4
    port map (
            O => \N__47696\,
            I => \ALU.bZ0Z_8\
        );

    \I__12105\ : ClkMux
    port map (
            O => \N__47693\,
            I => \N__47408\
        );

    \I__12104\ : ClkMux
    port map (
            O => \N__47692\,
            I => \N__47408\
        );

    \I__12103\ : ClkMux
    port map (
            O => \N__47691\,
            I => \N__47408\
        );

    \I__12102\ : ClkMux
    port map (
            O => \N__47690\,
            I => \N__47408\
        );

    \I__12101\ : ClkMux
    port map (
            O => \N__47689\,
            I => \N__47408\
        );

    \I__12100\ : ClkMux
    port map (
            O => \N__47688\,
            I => \N__47408\
        );

    \I__12099\ : ClkMux
    port map (
            O => \N__47687\,
            I => \N__47408\
        );

    \I__12098\ : ClkMux
    port map (
            O => \N__47686\,
            I => \N__47408\
        );

    \I__12097\ : ClkMux
    port map (
            O => \N__47685\,
            I => \N__47408\
        );

    \I__12096\ : ClkMux
    port map (
            O => \N__47684\,
            I => \N__47408\
        );

    \I__12095\ : ClkMux
    port map (
            O => \N__47683\,
            I => \N__47408\
        );

    \I__12094\ : ClkMux
    port map (
            O => \N__47682\,
            I => \N__47408\
        );

    \I__12093\ : ClkMux
    port map (
            O => \N__47681\,
            I => \N__47408\
        );

    \I__12092\ : ClkMux
    port map (
            O => \N__47680\,
            I => \N__47408\
        );

    \I__12091\ : ClkMux
    port map (
            O => \N__47679\,
            I => \N__47408\
        );

    \I__12090\ : ClkMux
    port map (
            O => \N__47678\,
            I => \N__47408\
        );

    \I__12089\ : ClkMux
    port map (
            O => \N__47677\,
            I => \N__47408\
        );

    \I__12088\ : ClkMux
    port map (
            O => \N__47676\,
            I => \N__47408\
        );

    \I__12087\ : ClkMux
    port map (
            O => \N__47675\,
            I => \N__47408\
        );

    \I__12086\ : ClkMux
    port map (
            O => \N__47674\,
            I => \N__47408\
        );

    \I__12085\ : ClkMux
    port map (
            O => \N__47673\,
            I => \N__47408\
        );

    \I__12084\ : ClkMux
    port map (
            O => \N__47672\,
            I => \N__47408\
        );

    \I__12083\ : ClkMux
    port map (
            O => \N__47671\,
            I => \N__47408\
        );

    \I__12082\ : ClkMux
    port map (
            O => \N__47670\,
            I => \N__47408\
        );

    \I__12081\ : ClkMux
    port map (
            O => \N__47669\,
            I => \N__47408\
        );

    \I__12080\ : ClkMux
    port map (
            O => \N__47668\,
            I => \N__47408\
        );

    \I__12079\ : ClkMux
    port map (
            O => \N__47667\,
            I => \N__47408\
        );

    \I__12078\ : ClkMux
    port map (
            O => \N__47666\,
            I => \N__47408\
        );

    \I__12077\ : ClkMux
    port map (
            O => \N__47665\,
            I => \N__47408\
        );

    \I__12076\ : ClkMux
    port map (
            O => \N__47664\,
            I => \N__47408\
        );

    \I__12075\ : ClkMux
    port map (
            O => \N__47663\,
            I => \N__47408\
        );

    \I__12074\ : ClkMux
    port map (
            O => \N__47662\,
            I => \N__47408\
        );

    \I__12073\ : ClkMux
    port map (
            O => \N__47661\,
            I => \N__47408\
        );

    \I__12072\ : ClkMux
    port map (
            O => \N__47660\,
            I => \N__47408\
        );

    \I__12071\ : ClkMux
    port map (
            O => \N__47659\,
            I => \N__47408\
        );

    \I__12070\ : ClkMux
    port map (
            O => \N__47658\,
            I => \N__47408\
        );

    \I__12069\ : ClkMux
    port map (
            O => \N__47657\,
            I => \N__47408\
        );

    \I__12068\ : ClkMux
    port map (
            O => \N__47656\,
            I => \N__47408\
        );

    \I__12067\ : ClkMux
    port map (
            O => \N__47655\,
            I => \N__47408\
        );

    \I__12066\ : ClkMux
    port map (
            O => \N__47654\,
            I => \N__47408\
        );

    \I__12065\ : ClkMux
    port map (
            O => \N__47653\,
            I => \N__47408\
        );

    \I__12064\ : ClkMux
    port map (
            O => \N__47652\,
            I => \N__47408\
        );

    \I__12063\ : ClkMux
    port map (
            O => \N__47651\,
            I => \N__47408\
        );

    \I__12062\ : ClkMux
    port map (
            O => \N__47650\,
            I => \N__47408\
        );

    \I__12061\ : ClkMux
    port map (
            O => \N__47649\,
            I => \N__47408\
        );

    \I__12060\ : ClkMux
    port map (
            O => \N__47648\,
            I => \N__47408\
        );

    \I__12059\ : ClkMux
    port map (
            O => \N__47647\,
            I => \N__47408\
        );

    \I__12058\ : ClkMux
    port map (
            O => \N__47646\,
            I => \N__47408\
        );

    \I__12057\ : ClkMux
    port map (
            O => \N__47645\,
            I => \N__47408\
        );

    \I__12056\ : ClkMux
    port map (
            O => \N__47644\,
            I => \N__47408\
        );

    \I__12055\ : ClkMux
    port map (
            O => \N__47643\,
            I => \N__47408\
        );

    \I__12054\ : ClkMux
    port map (
            O => \N__47642\,
            I => \N__47408\
        );

    \I__12053\ : ClkMux
    port map (
            O => \N__47641\,
            I => \N__47408\
        );

    \I__12052\ : ClkMux
    port map (
            O => \N__47640\,
            I => \N__47408\
        );

    \I__12051\ : ClkMux
    port map (
            O => \N__47639\,
            I => \N__47408\
        );

    \I__12050\ : ClkMux
    port map (
            O => \N__47638\,
            I => \N__47408\
        );

    \I__12049\ : ClkMux
    port map (
            O => \N__47637\,
            I => \N__47408\
        );

    \I__12048\ : ClkMux
    port map (
            O => \N__47636\,
            I => \N__47408\
        );

    \I__12047\ : ClkMux
    port map (
            O => \N__47635\,
            I => \N__47408\
        );

    \I__12046\ : ClkMux
    port map (
            O => \N__47634\,
            I => \N__47408\
        );

    \I__12045\ : ClkMux
    port map (
            O => \N__47633\,
            I => \N__47408\
        );

    \I__12044\ : ClkMux
    port map (
            O => \N__47632\,
            I => \N__47408\
        );

    \I__12043\ : ClkMux
    port map (
            O => \N__47631\,
            I => \N__47408\
        );

    \I__12042\ : ClkMux
    port map (
            O => \N__47630\,
            I => \N__47408\
        );

    \I__12041\ : ClkMux
    port map (
            O => \N__47629\,
            I => \N__47408\
        );

    \I__12040\ : ClkMux
    port map (
            O => \N__47628\,
            I => \N__47408\
        );

    \I__12039\ : ClkMux
    port map (
            O => \N__47627\,
            I => \N__47408\
        );

    \I__12038\ : ClkMux
    port map (
            O => \N__47626\,
            I => \N__47408\
        );

    \I__12037\ : ClkMux
    port map (
            O => \N__47625\,
            I => \N__47408\
        );

    \I__12036\ : ClkMux
    port map (
            O => \N__47624\,
            I => \N__47408\
        );

    \I__12035\ : ClkMux
    port map (
            O => \N__47623\,
            I => \N__47408\
        );

    \I__12034\ : ClkMux
    port map (
            O => \N__47622\,
            I => \N__47408\
        );

    \I__12033\ : ClkMux
    port map (
            O => \N__47621\,
            I => \N__47408\
        );

    \I__12032\ : ClkMux
    port map (
            O => \N__47620\,
            I => \N__47408\
        );

    \I__12031\ : ClkMux
    port map (
            O => \N__47619\,
            I => \N__47408\
        );

    \I__12030\ : ClkMux
    port map (
            O => \N__47618\,
            I => \N__47408\
        );

    \I__12029\ : ClkMux
    port map (
            O => \N__47617\,
            I => \N__47408\
        );

    \I__12028\ : ClkMux
    port map (
            O => \N__47616\,
            I => \N__47408\
        );

    \I__12027\ : ClkMux
    port map (
            O => \N__47615\,
            I => \N__47408\
        );

    \I__12026\ : ClkMux
    port map (
            O => \N__47614\,
            I => \N__47408\
        );

    \I__12025\ : ClkMux
    port map (
            O => \N__47613\,
            I => \N__47408\
        );

    \I__12024\ : ClkMux
    port map (
            O => \N__47612\,
            I => \N__47408\
        );

    \I__12023\ : ClkMux
    port map (
            O => \N__47611\,
            I => \N__47408\
        );

    \I__12022\ : ClkMux
    port map (
            O => \N__47610\,
            I => \N__47408\
        );

    \I__12021\ : ClkMux
    port map (
            O => \N__47609\,
            I => \N__47408\
        );

    \I__12020\ : ClkMux
    port map (
            O => \N__47608\,
            I => \N__47408\
        );

    \I__12019\ : ClkMux
    port map (
            O => \N__47607\,
            I => \N__47408\
        );

    \I__12018\ : ClkMux
    port map (
            O => \N__47606\,
            I => \N__47408\
        );

    \I__12017\ : ClkMux
    port map (
            O => \N__47605\,
            I => \N__47408\
        );

    \I__12016\ : ClkMux
    port map (
            O => \N__47604\,
            I => \N__47408\
        );

    \I__12015\ : ClkMux
    port map (
            O => \N__47603\,
            I => \N__47408\
        );

    \I__12014\ : ClkMux
    port map (
            O => \N__47602\,
            I => \N__47408\
        );

    \I__12013\ : ClkMux
    port map (
            O => \N__47601\,
            I => \N__47408\
        );

    \I__12012\ : ClkMux
    port map (
            O => \N__47600\,
            I => \N__47408\
        );

    \I__12011\ : ClkMux
    port map (
            O => \N__47599\,
            I => \N__47408\
        );

    \I__12010\ : GlobalMux
    port map (
            O => \N__47408\,
            I => \N__47405\
        );

    \I__12009\ : gio2CtrlBuf
    port map (
            O => \N__47405\,
            I => \CLK_0_c_g\
        );

    \I__12008\ : CEMux
    port map (
            O => \N__47402\,
            I => \N__47398\
        );

    \I__12007\ : CEMux
    port map (
            O => \N__47401\,
            I => \N__47394\
        );

    \I__12006\ : LocalMux
    port map (
            O => \N__47398\,
            I => \N__47390\
        );

    \I__12005\ : CEMux
    port map (
            O => \N__47397\,
            I => \N__47387\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__47394\,
            I => \N__47384\
        );

    \I__12003\ : CEMux
    port map (
            O => \N__47393\,
            I => \N__47381\
        );

    \I__12002\ : Span4Mux_h
    port map (
            O => \N__47390\,
            I => \N__47378\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__47387\,
            I => \N__47375\
        );

    \I__12000\ : Span4Mux_v
    port map (
            O => \N__47384\,
            I => \N__47372\
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__47381\,
            I => \N__47369\
        );

    \I__11998\ : Span4Mux_h
    port map (
            O => \N__47378\,
            I => \N__47366\
        );

    \I__11997\ : Span4Mux_h
    port map (
            O => \N__47375\,
            I => \N__47363\
        );

    \I__11996\ : Span4Mux_v
    port map (
            O => \N__47372\,
            I => \N__47360\
        );

    \I__11995\ : Span4Mux_h
    port map (
            O => \N__47369\,
            I => \N__47357\
        );

    \I__11994\ : Span4Mux_v
    port map (
            O => \N__47366\,
            I => \N__47354\
        );

    \I__11993\ : Span4Mux_v
    port map (
            O => \N__47363\,
            I => \N__47351\
        );

    \I__11992\ : Span4Mux_v
    port map (
            O => \N__47360\,
            I => \N__47348\
        );

    \I__11991\ : Sp12to4
    port map (
            O => \N__47357\,
            I => \N__47343\
        );

    \I__11990\ : Sp12to4
    port map (
            O => \N__47354\,
            I => \N__47343\
        );

    \I__11989\ : Span4Mux_v
    port map (
            O => \N__47351\,
            I => \N__47340\
        );

    \I__11988\ : Sp12to4
    port map (
            O => \N__47348\,
            I => \N__47337\
        );

    \I__11987\ : Span12Mux_h
    port map (
            O => \N__47343\,
            I => \N__47334\
        );

    \I__11986\ : Span4Mux_h
    port map (
            O => \N__47340\,
            I => \N__47331\
        );

    \I__11985\ : Odrv12
    port map (
            O => \N__47337\,
            I => \ALU.b_cnvZ0Z_0\
        );

    \I__11984\ : Odrv12
    port map (
            O => \N__47334\,
            I => \ALU.b_cnvZ0Z_0\
        );

    \I__11983\ : Odrv4
    port map (
            O => \N__47331\,
            I => \ALU.b_cnvZ0Z_0\
        );

    \I__11982\ : InMux
    port map (
            O => \N__47324\,
            I => \N__47315\
        );

    \I__11981\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47315\
        );

    \I__11980\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47311\
        );

    \I__11979\ : CascadeMux
    port map (
            O => \N__47321\,
            I => \N__47305\
        );

    \I__11978\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47300\
        );

    \I__11977\ : LocalMux
    port map (
            O => \N__47315\,
            I => \N__47297\
        );

    \I__11976\ : InMux
    port map (
            O => \N__47314\,
            I => \N__47294\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__47311\,
            I => \N__47289\
        );

    \I__11974\ : InMux
    port map (
            O => \N__47310\,
            I => \N__47286\
        );

    \I__11973\ : InMux
    port map (
            O => \N__47309\,
            I => \N__47283\
        );

    \I__11972\ : InMux
    port map (
            O => \N__47308\,
            I => \N__47280\
        );

    \I__11971\ : InMux
    port map (
            O => \N__47305\,
            I => \N__47274\
        );

    \I__11970\ : InMux
    port map (
            O => \N__47304\,
            I => \N__47269\
        );

    \I__11969\ : InMux
    port map (
            O => \N__47303\,
            I => \N__47269\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__47300\,
            I => \N__47264\
        );

    \I__11967\ : Span4Mux_v
    port map (
            O => \N__47297\,
            I => \N__47264\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__47294\,
            I => \N__47261\
        );

    \I__11965\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47256\
        );

    \I__11964\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47253\
        );

    \I__11963\ : Span4Mux_v
    port map (
            O => \N__47289\,
            I => \N__47246\
        );

    \I__11962\ : LocalMux
    port map (
            O => \N__47286\,
            I => \N__47246\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__47283\,
            I => \N__47246\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__47280\,
            I => \N__47243\
        );

    \I__11959\ : InMux
    port map (
            O => \N__47279\,
            I => \N__47238\
        );

    \I__11958\ : InMux
    port map (
            O => \N__47278\,
            I => \N__47238\
        );

    \I__11957\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47235\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__47274\,
            I => \N__47224\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__47269\,
            I => \N__47224\
        );

    \I__11954\ : Span4Mux_v
    port map (
            O => \N__47264\,
            I => \N__47221\
        );

    \I__11953\ : Span4Mux_v
    port map (
            O => \N__47261\,
            I => \N__47217\
        );

    \I__11952\ : InMux
    port map (
            O => \N__47260\,
            I => \N__47212\
        );

    \I__11951\ : InMux
    port map (
            O => \N__47259\,
            I => \N__47212\
        );

    \I__11950\ : LocalMux
    port map (
            O => \N__47256\,
            I => \N__47205\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__47253\,
            I => \N__47205\
        );

    \I__11948\ : Span4Mux_v
    port map (
            O => \N__47246\,
            I => \N__47202\
        );

    \I__11947\ : Span4Mux_v
    port map (
            O => \N__47243\,
            I => \N__47199\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__47238\,
            I => \N__47194\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__47235\,
            I => \N__47194\
        );

    \I__11944\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47185\
        );

    \I__11943\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47185\
        );

    \I__11942\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47185\
        );

    \I__11941\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47185\
        );

    \I__11940\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47180\
        );

    \I__11939\ : InMux
    port map (
            O => \N__47229\,
            I => \N__47180\
        );

    \I__11938\ : Span4Mux_v
    port map (
            O => \N__47224\,
            I => \N__47173\
        );

    \I__11937\ : Span4Mux_h
    port map (
            O => \N__47221\,
            I => \N__47173\
        );

    \I__11936\ : InMux
    port map (
            O => \N__47220\,
            I => \N__47170\
        );

    \I__11935\ : Span4Mux_h
    port map (
            O => \N__47217\,
            I => \N__47165\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47165\
        );

    \I__11933\ : InMux
    port map (
            O => \N__47211\,
            I => \N__47160\
        );

    \I__11932\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47160\
        );

    \I__11931\ : Span4Mux_v
    port map (
            O => \N__47205\,
            I => \N__47157\
        );

    \I__11930\ : Span4Mux_v
    port map (
            O => \N__47202\,
            I => \N__47154\
        );

    \I__11929\ : Span4Mux_v
    port map (
            O => \N__47199\,
            I => \N__47151\
        );

    \I__11928\ : Span4Mux_v
    port map (
            O => \N__47194\,
            I => \N__47146\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__47185\,
            I => \N__47146\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__47180\,
            I => \N__47143\
        );

    \I__11925\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47140\
        );

    \I__11924\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47137\
        );

    \I__11923\ : Span4Mux_v
    port map (
            O => \N__47173\,
            I => \N__47134\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__47170\,
            I => \N__47125\
        );

    \I__11921\ : Span4Mux_v
    port map (
            O => \N__47165\,
            I => \N__47125\
        );

    \I__11920\ : LocalMux
    port map (
            O => \N__47160\,
            I => \N__47125\
        );

    \I__11919\ : Span4Mux_h
    port map (
            O => \N__47157\,
            I => \N__47125\
        );

    \I__11918\ : Span4Mux_h
    port map (
            O => \N__47154\,
            I => \N__47116\
        );

    \I__11917\ : Span4Mux_h
    port map (
            O => \N__47151\,
            I => \N__47116\
        );

    \I__11916\ : Span4Mux_v
    port map (
            O => \N__47146\,
            I => \N__47116\
        );

    \I__11915\ : Span4Mux_s2_v
    port map (
            O => \N__47143\,
            I => \N__47116\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__47140\,
            I => \ALU.a_15_sm0\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__47137\,
            I => \ALU.a_15_sm0\
        );

    \I__11912\ : Odrv4
    port map (
            O => \N__47134\,
            I => \ALU.a_15_sm0\
        );

    \I__11911\ : Odrv4
    port map (
            O => \N__47125\,
            I => \ALU.a_15_sm0\
        );

    \I__11910\ : Odrv4
    port map (
            O => \N__47116\,
            I => \ALU.a_15_sm0\
        );

    \I__11909\ : InMux
    port map (
            O => \N__47105\,
            I => \N__47102\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__47102\,
            I => \N__47093\
        );

    \I__11907\ : InMux
    port map (
            O => \N__47101\,
            I => \N__47090\
        );

    \I__11906\ : InMux
    port map (
            O => \N__47100\,
            I => \N__47084\
        );

    \I__11905\ : InMux
    port map (
            O => \N__47099\,
            I => \N__47077\
        );

    \I__11904\ : InMux
    port map (
            O => \N__47098\,
            I => \N__47077\
        );

    \I__11903\ : InMux
    port map (
            O => \N__47097\,
            I => \N__47077\
        );

    \I__11902\ : InMux
    port map (
            O => \N__47096\,
            I => \N__47074\
        );

    \I__11901\ : Span4Mux_v
    port map (
            O => \N__47093\,
            I => \N__47071\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__47090\,
            I => \N__47068\
        );

    \I__11899\ : InMux
    port map (
            O => \N__47089\,
            I => \N__47064\
        );

    \I__11898\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47061\
        );

    \I__11897\ : InMux
    port map (
            O => \N__47087\,
            I => \N__47058\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__47084\,
            I => \N__47055\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__47077\,
            I => \N__47052\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__47074\,
            I => \N__47046\
        );

    \I__11893\ : Span4Mux_h
    port map (
            O => \N__47071\,
            I => \N__47043\
        );

    \I__11892\ : Span4Mux_v
    port map (
            O => \N__47068\,
            I => \N__47040\
        );

    \I__11891\ : InMux
    port map (
            O => \N__47067\,
            I => \N__47037\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__47064\,
            I => \N__47032\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__47061\,
            I => \N__47032\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__47058\,
            I => \N__47025\
        );

    \I__11887\ : Span4Mux_h
    port map (
            O => \N__47055\,
            I => \N__47025\
        );

    \I__11886\ : Span4Mux_v
    port map (
            O => \N__47052\,
            I => \N__47025\
        );

    \I__11885\ : InMux
    port map (
            O => \N__47051\,
            I => \N__47022\
        );

    \I__11884\ : InMux
    port map (
            O => \N__47050\,
            I => \N__47017\
        );

    \I__11883\ : InMux
    port map (
            O => \N__47049\,
            I => \N__47017\
        );

    \I__11882\ : Span4Mux_v
    port map (
            O => \N__47046\,
            I => \N__47014\
        );

    \I__11881\ : Span4Mux_h
    port map (
            O => \N__47043\,
            I => \N__47005\
        );

    \I__11880\ : Span4Mux_v
    port map (
            O => \N__47040\,
            I => \N__47005\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__47037\,
            I => \N__47005\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__47032\,
            I => \N__47005\
        );

    \I__11877\ : Span4Mux_v
    port map (
            O => \N__47025\,
            I => \N__47002\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__47022\,
            I => \ALU.N_213_0\
        );

    \I__11875\ : LocalMux
    port map (
            O => \N__47017\,
            I => \ALU.N_213_0\
        );

    \I__11874\ : Odrv4
    port map (
            O => \N__47014\,
            I => \ALU.N_213_0\
        );

    \I__11873\ : Odrv4
    port map (
            O => \N__47005\,
            I => \ALU.N_213_0\
        );

    \I__11872\ : Odrv4
    port map (
            O => \N__47002\,
            I => \ALU.N_213_0\
        );

    \I__11871\ : CascadeMux
    port map (
            O => \N__46991\,
            I => \N__46988\
        );

    \I__11870\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46985\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__46985\,
            I => \N__46982\
        );

    \I__11868\ : Span4Mux_h
    port map (
            O => \N__46982\,
            I => \N__46979\
        );

    \I__11867\ : Odrv4
    port map (
            O => \N__46979\,
            I => \ALU.a_15_m2_ns_1Z0Z_7\
        );

    \I__11866\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46970\
        );

    \I__11865\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46967\
        );

    \I__11864\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46957\
        );

    \I__11863\ : CascadeMux
    port map (
            O => \N__46973\,
            I => \N__46953\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__46970\,
            I => \N__46950\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__46967\,
            I => \N__46947\
        );

    \I__11860\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46937\
        );

    \I__11859\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46937\
        );

    \I__11858\ : InMux
    port map (
            O => \N__46964\,
            I => \N__46934\
        );

    \I__11857\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46931\
        );

    \I__11856\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46928\
        );

    \I__11855\ : InMux
    port map (
            O => \N__46961\,
            I => \N__46925\
        );

    \I__11854\ : InMux
    port map (
            O => \N__46960\,
            I => \N__46922\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__46957\,
            I => \N__46919\
        );

    \I__11852\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46913\
        );

    \I__11851\ : InMux
    port map (
            O => \N__46953\,
            I => \N__46913\
        );

    \I__11850\ : Span4Mux_h
    port map (
            O => \N__46950\,
            I => \N__46908\
        );

    \I__11849\ : Span4Mux_h
    port map (
            O => \N__46947\,
            I => \N__46904\
        );

    \I__11848\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46899\
        );

    \I__11847\ : InMux
    port map (
            O => \N__46945\,
            I => \N__46899\
        );

    \I__11846\ : InMux
    port map (
            O => \N__46944\,
            I => \N__46896\
        );

    \I__11845\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46893\
        );

    \I__11844\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46890\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__46937\,
            I => \N__46887\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__46934\,
            I => \N__46884\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__46931\,
            I => \N__46877\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__46928\,
            I => \N__46877\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__46925\,
            I => \N__46877\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__46922\,
            I => \N__46873\
        );

    \I__11837\ : Span4Mux_h
    port map (
            O => \N__46919\,
            I => \N__46870\
        );

    \I__11836\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46867\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__46913\,
            I => \N__46864\
        );

    \I__11834\ : InMux
    port map (
            O => \N__46912\,
            I => \N__46861\
        );

    \I__11833\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46858\
        );

    \I__11832\ : Span4Mux_h
    port map (
            O => \N__46908\,
            I => \N__46855\
        );

    \I__11831\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46852\
        );

    \I__11830\ : Span4Mux_h
    port map (
            O => \N__46904\,
            I => \N__46847\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__46899\,
            I => \N__46847\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__46896\,
            I => \N__46840\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__46893\,
            I => \N__46840\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__46890\,
            I => \N__46840\
        );

    \I__11825\ : Span4Mux_h
    port map (
            O => \N__46887\,
            I => \N__46834\
        );

    \I__11824\ : Span4Mux_h
    port map (
            O => \N__46884\,
            I => \N__46831\
        );

    \I__11823\ : Span4Mux_v
    port map (
            O => \N__46877\,
            I => \N__46828\
        );

    \I__11822\ : InMux
    port map (
            O => \N__46876\,
            I => \N__46825\
        );

    \I__11821\ : Span4Mux_v
    port map (
            O => \N__46873\,
            I => \N__46820\
        );

    \I__11820\ : Span4Mux_v
    port map (
            O => \N__46870\,
            I => \N__46820\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__46867\,
            I => \N__46817\
        );

    \I__11818\ : Span4Mux_v
    port map (
            O => \N__46864\,
            I => \N__46814\
        );

    \I__11817\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46808\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__46858\,
            I => \N__46808\
        );

    \I__11815\ : Span4Mux_h
    port map (
            O => \N__46855\,
            I => \N__46799\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__46852\,
            I => \N__46799\
        );

    \I__11813\ : Span4Mux_v
    port map (
            O => \N__46847\,
            I => \N__46799\
        );

    \I__11812\ : Span4Mux_h
    port map (
            O => \N__46840\,
            I => \N__46799\
        );

    \I__11811\ : InMux
    port map (
            O => \N__46839\,
            I => \N__46794\
        );

    \I__11810\ : InMux
    port map (
            O => \N__46838\,
            I => \N__46794\
        );

    \I__11809\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46791\
        );

    \I__11808\ : Span4Mux_v
    port map (
            O => \N__46834\,
            I => \N__46788\
        );

    \I__11807\ : Span4Mux_h
    port map (
            O => \N__46831\,
            I => \N__46783\
        );

    \I__11806\ : Span4Mux_s2_h
    port map (
            O => \N__46828\,
            I => \N__46783\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__46825\,
            I => \N__46780\
        );

    \I__11804\ : Span4Mux_v
    port map (
            O => \N__46820\,
            I => \N__46773\
        );

    \I__11803\ : Span4Mux_h
    port map (
            O => \N__46817\,
            I => \N__46773\
        );

    \I__11802\ : Span4Mux_h
    port map (
            O => \N__46814\,
            I => \N__46773\
        );

    \I__11801\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46770\
        );

    \I__11800\ : Span4Mux_h
    port map (
            O => \N__46808\,
            I => \N__46763\
        );

    \I__11799\ : Span4Mux_v
    port map (
            O => \N__46799\,
            I => \N__46763\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__46794\,
            I => \N__46763\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__46791\,
            I => \ALU.aluOut_7\
        );

    \I__11796\ : Odrv4
    port map (
            O => \N__46788\,
            I => \ALU.aluOut_7\
        );

    \I__11795\ : Odrv4
    port map (
            O => \N__46783\,
            I => \ALU.aluOut_7\
        );

    \I__11794\ : Odrv12
    port map (
            O => \N__46780\,
            I => \ALU.aluOut_7\
        );

    \I__11793\ : Odrv4
    port map (
            O => \N__46773\,
            I => \ALU.aluOut_7\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__46770\,
            I => \ALU.aluOut_7\
        );

    \I__11791\ : Odrv4
    port map (
            O => \N__46763\,
            I => \ALU.aluOut_7\
        );

    \I__11790\ : CascadeMux
    port map (
            O => \N__46748\,
            I => \N__46745\
        );

    \I__11789\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46742\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46739\
        );

    \I__11787\ : Odrv4
    port map (
            O => \N__46739\,
            I => \ALU.a_15_m2_7\
        );

    \I__11786\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46730\
        );

    \I__11785\ : InMux
    port map (
            O => \N__46735\,
            I => \N__46724\
        );

    \I__11784\ : InMux
    port map (
            O => \N__46734\,
            I => \N__46721\
        );

    \I__11783\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46717\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__46730\,
            I => \N__46712\
        );

    \I__11781\ : InMux
    port map (
            O => \N__46729\,
            I => \N__46709\
        );

    \I__11780\ : InMux
    port map (
            O => \N__46728\,
            I => \N__46706\
        );

    \I__11779\ : InMux
    port map (
            O => \N__46727\,
            I => \N__46703\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__46724\,
            I => \N__46700\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__46721\,
            I => \N__46697\
        );

    \I__11776\ : InMux
    port map (
            O => \N__46720\,
            I => \N__46694\
        );

    \I__11775\ : LocalMux
    port map (
            O => \N__46717\,
            I => \N__46690\
        );

    \I__11774\ : InMux
    port map (
            O => \N__46716\,
            I => \N__46687\
        );

    \I__11773\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46683\
        );

    \I__11772\ : Span4Mux_s3_h
    port map (
            O => \N__46712\,
            I => \N__46676\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__46709\,
            I => \N__46676\
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__46706\,
            I => \N__46673\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__46703\,
            I => \N__46666\
        );

    \I__11768\ : Span4Mux_h
    port map (
            O => \N__46700\,
            I => \N__46659\
        );

    \I__11767\ : Span4Mux_s2_v
    port map (
            O => \N__46697\,
            I => \N__46659\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__46694\,
            I => \N__46659\
        );

    \I__11765\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46654\
        );

    \I__11764\ : Span4Mux_v
    port map (
            O => \N__46690\,
            I => \N__46649\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__46687\,
            I => \N__46649\
        );

    \I__11762\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46645\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46642\
        );

    \I__11760\ : CascadeMux
    port map (
            O => \N__46682\,
            I => \N__46639\
        );

    \I__11759\ : InMux
    port map (
            O => \N__46681\,
            I => \N__46635\
        );

    \I__11758\ : Span4Mux_h
    port map (
            O => \N__46676\,
            I => \N__46630\
        );

    \I__11757\ : Span4Mux_s3_h
    port map (
            O => \N__46673\,
            I => \N__46630\
        );

    \I__11756\ : InMux
    port map (
            O => \N__46672\,
            I => \N__46627\
        );

    \I__11755\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46623\
        );

    \I__11754\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46617\
        );

    \I__11753\ : InMux
    port map (
            O => \N__46669\,
            I => \N__46617\
        );

    \I__11752\ : Span4Mux_v
    port map (
            O => \N__46666\,
            I => \N__46612\
        );

    \I__11751\ : Span4Mux_v
    port map (
            O => \N__46659\,
            I => \N__46609\
        );

    \I__11750\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46606\
        );

    \I__11749\ : InMux
    port map (
            O => \N__46657\,
            I => \N__46603\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__46654\,
            I => \N__46600\
        );

    \I__11747\ : Span4Mux_h
    port map (
            O => \N__46649\,
            I => \N__46597\
        );

    \I__11746\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46594\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__46645\,
            I => \N__46589\
        );

    \I__11744\ : Span4Mux_v
    port map (
            O => \N__46642\,
            I => \N__46589\
        );

    \I__11743\ : InMux
    port map (
            O => \N__46639\,
            I => \N__46586\
        );

    \I__11742\ : InMux
    port map (
            O => \N__46638\,
            I => \N__46583\
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__46635\,
            I => \N__46576\
        );

    \I__11740\ : Span4Mux_v
    port map (
            O => \N__46630\,
            I => \N__46576\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__46627\,
            I => \N__46576\
        );

    \I__11738\ : InMux
    port map (
            O => \N__46626\,
            I => \N__46573\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__46623\,
            I => \N__46570\
        );

    \I__11736\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46567\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46564\
        );

    \I__11734\ : InMux
    port map (
            O => \N__46616\,
            I => \N__46559\
        );

    \I__11733\ : InMux
    port map (
            O => \N__46615\,
            I => \N__46559\
        );

    \I__11732\ : Span4Mux_v
    port map (
            O => \N__46612\,
            I => \N__46556\
        );

    \I__11731\ : Span4Mux_v
    port map (
            O => \N__46609\,
            I => \N__46551\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__46606\,
            I => \N__46551\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__46603\,
            I => \N__46546\
        );

    \I__11728\ : Span4Mux_h
    port map (
            O => \N__46600\,
            I => \N__46546\
        );

    \I__11727\ : Span4Mux_v
    port map (
            O => \N__46597\,
            I => \N__46543\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__46594\,
            I => \N__46538\
        );

    \I__11725\ : Span4Mux_h
    port map (
            O => \N__46589\,
            I => \N__46538\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__46586\,
            I => \N__46535\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__46583\,
            I => \N__46530\
        );

    \I__11722\ : Span4Mux_v
    port map (
            O => \N__46576\,
            I => \N__46530\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__46573\,
            I => \N__46525\
        );

    \I__11720\ : Span4Mux_v
    port map (
            O => \N__46570\,
            I => \N__46525\
        );

    \I__11719\ : LocalMux
    port map (
            O => \N__46567\,
            I => \N__46522\
        );

    \I__11718\ : Span12Mux_v
    port map (
            O => \N__46564\,
            I => \N__46517\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__46559\,
            I => \N__46517\
        );

    \I__11716\ : Span4Mux_h
    port map (
            O => \N__46556\,
            I => \N__46512\
        );

    \I__11715\ : Span4Mux_v
    port map (
            O => \N__46551\,
            I => \N__46512\
        );

    \I__11714\ : Span4Mux_h
    port map (
            O => \N__46546\,
            I => \N__46509\
        );

    \I__11713\ : Span4Mux_v
    port map (
            O => \N__46543\,
            I => \N__46504\
        );

    \I__11712\ : Span4Mux_h
    port map (
            O => \N__46538\,
            I => \N__46504\
        );

    \I__11711\ : Span4Mux_v
    port map (
            O => \N__46535\,
            I => \N__46495\
        );

    \I__11710\ : Span4Mux_h
    port map (
            O => \N__46530\,
            I => \N__46495\
        );

    \I__11709\ : Span4Mux_h
    port map (
            O => \N__46525\,
            I => \N__46495\
        );

    \I__11708\ : Span4Mux_v
    port map (
            O => \N__46522\,
            I => \N__46495\
        );

    \I__11707\ : Odrv12
    port map (
            O => \N__46517\,
            I => \ALU.aluOut_6\
        );

    \I__11706\ : Odrv4
    port map (
            O => \N__46512\,
            I => \ALU.aluOut_6\
        );

    \I__11705\ : Odrv4
    port map (
            O => \N__46509\,
            I => \ALU.aluOut_6\
        );

    \I__11704\ : Odrv4
    port map (
            O => \N__46504\,
            I => \ALU.aluOut_6\
        );

    \I__11703\ : Odrv4
    port map (
            O => \N__46495\,
            I => \ALU.aluOut_6\
        );

    \I__11702\ : CascadeMux
    port map (
            O => \N__46484\,
            I => \ALU.a_15_m2_ns_1Z0Z_6_cascade_\
        );

    \I__11701\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46478\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__46478\,
            I => \N__46475\
        );

    \I__11699\ : Span4Mux_v
    port map (
            O => \N__46475\,
            I => \N__46470\
        );

    \I__11698\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46467\
        );

    \I__11697\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46464\
        );

    \I__11696\ : Span4Mux_h
    port map (
            O => \N__46470\,
            I => \N__46459\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__46467\,
            I => \N__46456\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__46464\,
            I => \N__46453\
        );

    \I__11693\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46450\
        );

    \I__11692\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46445\
        );

    \I__11691\ : Span4Mux_h
    port map (
            O => \N__46459\,
            I => \N__46438\
        );

    \I__11690\ : Span4Mux_v
    port map (
            O => \N__46456\,
            I => \N__46438\
        );

    \I__11689\ : Span4Mux_h
    port map (
            O => \N__46453\,
            I => \N__46433\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46433\
        );

    \I__11687\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46430\
        );

    \I__11686\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46427\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__46445\,
            I => \N__46424\
        );

    \I__11684\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46421\
        );

    \I__11683\ : InMux
    port map (
            O => \N__46443\,
            I => \N__46418\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__46438\,
            I => \N__46413\
        );

    \I__11681\ : Span4Mux_v
    port map (
            O => \N__46433\,
            I => \N__46413\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__46430\,
            I => \ALU.N_219_0\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__46427\,
            I => \ALU.N_219_0\
        );

    \I__11678\ : Odrv4
    port map (
            O => \N__46424\,
            I => \ALU.N_219_0\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__46421\,
            I => \ALU.N_219_0\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__46418\,
            I => \ALU.N_219_0\
        );

    \I__11675\ : Odrv4
    port map (
            O => \N__46413\,
            I => \ALU.N_219_0\
        );

    \I__11674\ : InMux
    port map (
            O => \N__46400\,
            I => \N__46397\
        );

    \I__11673\ : LocalMux
    port map (
            O => \N__46397\,
            I => \ALU.a_15_m2_6\
        );

    \I__11672\ : InMux
    port map (
            O => \N__46394\,
            I => \N__46388\
        );

    \I__11671\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46385\
        );

    \I__11670\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46379\
        );

    \I__11669\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46376\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__46388\,
            I => \N__46373\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__46385\,
            I => \N__46370\
        );

    \I__11666\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46367\
        );

    \I__11665\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46364\
        );

    \I__11664\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46359\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__46379\,
            I => \N__46354\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__46376\,
            I => \N__46354\
        );

    \I__11661\ : Span4Mux_v
    port map (
            O => \N__46373\,
            I => \N__46349\
        );

    \I__11660\ : Span4Mux_h
    port map (
            O => \N__46370\,
            I => \N__46346\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__46367\,
            I => \N__46343\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__46364\,
            I => \N__46340\
        );

    \I__11657\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46335\
        );

    \I__11656\ : InMux
    port map (
            O => \N__46362\,
            I => \N__46335\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46332\
        );

    \I__11654\ : Span4Mux_h
    port map (
            O => \N__46354\,
            I => \N__46327\
        );

    \I__11653\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46323\
        );

    \I__11652\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46320\
        );

    \I__11651\ : Span4Mux_v
    port map (
            O => \N__46349\,
            I => \N__46317\
        );

    \I__11650\ : Sp12to4
    port map (
            O => \N__46346\,
            I => \N__46312\
        );

    \I__11649\ : Span12Mux_h
    port map (
            O => \N__46343\,
            I => \N__46312\
        );

    \I__11648\ : Span4Mux_v
    port map (
            O => \N__46340\,
            I => \N__46305\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__46335\,
            I => \N__46305\
        );

    \I__11646\ : Span4Mux_v
    port map (
            O => \N__46332\,
            I => \N__46302\
        );

    \I__11645\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46299\
        );

    \I__11644\ : InMux
    port map (
            O => \N__46330\,
            I => \N__46296\
        );

    \I__11643\ : Span4Mux_h
    port map (
            O => \N__46327\,
            I => \N__46293\
        );

    \I__11642\ : InMux
    port map (
            O => \N__46326\,
            I => \N__46290\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__46323\,
            I => \N__46285\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__46320\,
            I => \N__46285\
        );

    \I__11639\ : Sp12to4
    port map (
            O => \N__46317\,
            I => \N__46280\
        );

    \I__11638\ : Span12Mux_v
    port map (
            O => \N__46312\,
            I => \N__46280\
        );

    \I__11637\ : InMux
    port map (
            O => \N__46311\,
            I => \N__46277\
        );

    \I__11636\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46274\
        );

    \I__11635\ : IoSpan4Mux
    port map (
            O => \N__46305\,
            I => \N__46271\
        );

    \I__11634\ : Span4Mux_h
    port map (
            O => \N__46302\,
            I => \N__46266\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__46299\,
            I => \N__46266\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__46296\,
            I => \N__46259\
        );

    \I__11631\ : Span4Mux_v
    port map (
            O => \N__46293\,
            I => \N__46259\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__46290\,
            I => \N__46259\
        );

    \I__11629\ : Span12Mux_v
    port map (
            O => \N__46285\,
            I => \N__46256\
        );

    \I__11628\ : Span12Mux_h
    port map (
            O => \N__46280\,
            I => \N__46253\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__46277\,
            I => \N__46250\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__46274\,
            I => \N__46245\
        );

    \I__11625\ : IoSpan4Mux
    port map (
            O => \N__46271\,
            I => \N__46245\
        );

    \I__11624\ : Span4Mux_v
    port map (
            O => \N__46266\,
            I => \N__46240\
        );

    \I__11623\ : Span4Mux_v
    port map (
            O => \N__46259\,
            I => \N__46240\
        );

    \I__11622\ : Odrv12
    port map (
            O => \N__46256\,
            I => \ALU.a_15_sm3\
        );

    \I__11621\ : Odrv12
    port map (
            O => \N__46253\,
            I => \ALU.a_15_sm3\
        );

    \I__11620\ : Odrv4
    port map (
            O => \N__46250\,
            I => \ALU.a_15_sm3\
        );

    \I__11619\ : Odrv4
    port map (
            O => \N__46245\,
            I => \ALU.a_15_sm3\
        );

    \I__11618\ : Odrv4
    port map (
            O => \N__46240\,
            I => \ALU.a_15_sm3\
        );

    \I__11617\ : InMux
    port map (
            O => \N__46229\,
            I => \N__46226\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__46226\,
            I => \N__46223\
        );

    \I__11615\ : Span4Mux_h
    port map (
            O => \N__46223\,
            I => \N__46220\
        );

    \I__11614\ : Span4Mux_h
    port map (
            O => \N__46220\,
            I => \N__46217\
        );

    \I__11613\ : Span4Mux_h
    port map (
            O => \N__46217\,
            I => \N__46214\
        );

    \I__11612\ : Span4Mux_v
    port map (
            O => \N__46214\,
            I => \N__46211\
        );

    \I__11611\ : Odrv4
    port map (
            O => \N__46211\,
            I => \ALU.d_RNIL01TD1Z0Z_6\
        );

    \I__11610\ : InMux
    port map (
            O => \N__46208\,
            I => \N__46205\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__46205\,
            I => \ALU.d_RNIJ75U41Z0Z_6\
        );

    \I__11608\ : CascadeMux
    port map (
            O => \N__46202\,
            I => \N__46197\
        );

    \I__11607\ : CascadeMux
    port map (
            O => \N__46201\,
            I => \N__46194\
        );

    \I__11606\ : CascadeMux
    port map (
            O => \N__46200\,
            I => \N__46186\
        );

    \I__11605\ : InMux
    port map (
            O => \N__46197\,
            I => \N__46181\
        );

    \I__11604\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46181\
        );

    \I__11603\ : CascadeMux
    port map (
            O => \N__46193\,
            I => \N__46178\
        );

    \I__11602\ : CascadeMux
    port map (
            O => \N__46192\,
            I => \N__46175\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__46191\,
            I => \N__46172\
        );

    \I__11600\ : CascadeMux
    port map (
            O => \N__46190\,
            I => \N__46169\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__46189\,
            I => \N__46166\
        );

    \I__11598\ : InMux
    port map (
            O => \N__46186\,
            I => \N__46144\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__46181\,
            I => \N__46141\
        );

    \I__11596\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46138\
        );

    \I__11595\ : InMux
    port map (
            O => \N__46175\,
            I => \N__46123\
        );

    \I__11594\ : InMux
    port map (
            O => \N__46172\,
            I => \N__46123\
        );

    \I__11593\ : InMux
    port map (
            O => \N__46169\,
            I => \N__46123\
        );

    \I__11592\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46123\
        );

    \I__11591\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46123\
        );

    \I__11590\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46123\
        );

    \I__11589\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46123\
        );

    \I__11588\ : CascadeMux
    port map (
            O => \N__46162\,
            I => \N__46119\
        );

    \I__11587\ : CascadeMux
    port map (
            O => \N__46161\,
            I => \N__46114\
        );

    \I__11586\ : CascadeMux
    port map (
            O => \N__46160\,
            I => \N__46111\
        );

    \I__11585\ : CascadeMux
    port map (
            O => \N__46159\,
            I => \N__46108\
        );

    \I__11584\ : CascadeMux
    port map (
            O => \N__46158\,
            I => \N__46105\
        );

    \I__11583\ : CascadeMux
    port map (
            O => \N__46157\,
            I => \N__46102\
        );

    \I__11582\ : CascadeMux
    port map (
            O => \N__46156\,
            I => \N__46099\
        );

    \I__11581\ : CascadeMux
    port map (
            O => \N__46155\,
            I => \N__46095\
        );

    \I__11580\ : CascadeMux
    port map (
            O => \N__46154\,
            I => \N__46092\
        );

    \I__11579\ : CascadeMux
    port map (
            O => \N__46153\,
            I => \N__46089\
        );

    \I__11578\ : CascadeMux
    port map (
            O => \N__46152\,
            I => \N__46086\
        );

    \I__11577\ : CascadeMux
    port map (
            O => \N__46151\,
            I => \N__46073\
        );

    \I__11576\ : CascadeMux
    port map (
            O => \N__46150\,
            I => \N__46070\
        );

    \I__11575\ : CascadeMux
    port map (
            O => \N__46149\,
            I => \N__46067\
        );

    \I__11574\ : CascadeMux
    port map (
            O => \N__46148\,
            I => \N__46064\
        );

    \I__11573\ : CascadeMux
    port map (
            O => \N__46147\,
            I => \N__46061\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__46144\,
            I => \N__46057\
        );

    \I__11571\ : Span4Mux_h
    port map (
            O => \N__46141\,
            I => \N__46050\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__46138\,
            I => \N__46050\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__46123\,
            I => \N__46050\
        );

    \I__11568\ : CascadeMux
    port map (
            O => \N__46122\,
            I => \N__46047\
        );

    \I__11567\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46042\
        );

    \I__11566\ : CascadeMux
    port map (
            O => \N__46118\,
            I => \N__46037\
        );

    \I__11565\ : CascadeMux
    port map (
            O => \N__46117\,
            I => \N__46034\
        );

    \I__11564\ : InMux
    port map (
            O => \N__46114\,
            I => \N__46024\
        );

    \I__11563\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46024\
        );

    \I__11562\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46024\
        );

    \I__11561\ : InMux
    port map (
            O => \N__46105\,
            I => \N__46024\
        );

    \I__11560\ : InMux
    port map (
            O => \N__46102\,
            I => \N__46017\
        );

    \I__11559\ : InMux
    port map (
            O => \N__46099\,
            I => \N__46017\
        );

    \I__11558\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46017\
        );

    \I__11557\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46008\
        );

    \I__11556\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46008\
        );

    \I__11555\ : InMux
    port map (
            O => \N__46089\,
            I => \N__46008\
        );

    \I__11554\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46008\
        );

    \I__11553\ : InMux
    port map (
            O => \N__46085\,
            I => \N__46005\
        );

    \I__11552\ : CascadeMux
    port map (
            O => \N__46084\,
            I => \N__45997\
        );

    \I__11551\ : CascadeMux
    port map (
            O => \N__46083\,
            I => \N__45994\
        );

    \I__11550\ : CascadeMux
    port map (
            O => \N__46082\,
            I => \N__45986\
        );

    \I__11549\ : CascadeMux
    port map (
            O => \N__46081\,
            I => \N__45983\
        );

    \I__11548\ : CascadeMux
    port map (
            O => \N__46080\,
            I => \N__45980\
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__46079\,
            I => \N__45977\
        );

    \I__11546\ : CascadeMux
    port map (
            O => \N__46078\,
            I => \N__45974\
        );

    \I__11545\ : CascadeMux
    port map (
            O => \N__46077\,
            I => \N__45971\
        );

    \I__11544\ : CascadeMux
    port map (
            O => \N__46076\,
            I => \N__45968\
        );

    \I__11543\ : InMux
    port map (
            O => \N__46073\,
            I => \N__45962\
        );

    \I__11542\ : InMux
    port map (
            O => \N__46070\,
            I => \N__45962\
        );

    \I__11541\ : InMux
    port map (
            O => \N__46067\,
            I => \N__45953\
        );

    \I__11540\ : InMux
    port map (
            O => \N__46064\,
            I => \N__45953\
        );

    \I__11539\ : InMux
    port map (
            O => \N__46061\,
            I => \N__45953\
        );

    \I__11538\ : InMux
    port map (
            O => \N__46060\,
            I => \N__45953\
        );

    \I__11537\ : Span4Mux_h
    port map (
            O => \N__46057\,
            I => \N__45950\
        );

    \I__11536\ : Span4Mux_v
    port map (
            O => \N__46050\,
            I => \N__45947\
        );

    \I__11535\ : InMux
    port map (
            O => \N__46047\,
            I => \N__45940\
        );

    \I__11534\ : InMux
    port map (
            O => \N__46046\,
            I => \N__45940\
        );

    \I__11533\ : InMux
    port map (
            O => \N__46045\,
            I => \N__45940\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__46042\,
            I => \N__45937\
        );

    \I__11531\ : InMux
    port map (
            O => \N__46041\,
            I => \N__45934\
        );

    \I__11530\ : InMux
    port map (
            O => \N__46040\,
            I => \N__45931\
        );

    \I__11529\ : InMux
    port map (
            O => \N__46037\,
            I => \N__45927\
        );

    \I__11528\ : InMux
    port map (
            O => \N__46034\,
            I => \N__45924\
        );

    \I__11527\ : InMux
    port map (
            O => \N__46033\,
            I => \N__45920\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__46024\,
            I => \N__45913\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__46017\,
            I => \N__45913\
        );

    \I__11524\ : LocalMux
    port map (
            O => \N__46008\,
            I => \N__45913\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__45910\
        );

    \I__11522\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45907\
        );

    \I__11521\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45904\
        );

    \I__11520\ : CascadeMux
    port map (
            O => \N__46002\,
            I => \N__45900\
        );

    \I__11519\ : CascadeMux
    port map (
            O => \N__46001\,
            I => \N__45897\
        );

    \I__11518\ : CascadeMux
    port map (
            O => \N__46000\,
            I => \N__45894\
        );

    \I__11517\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45886\
        );

    \I__11516\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45886\
        );

    \I__11515\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45886\
        );

    \I__11514\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45883\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__45991\,
            I => \N__45880\
        );

    \I__11512\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45877\
        );

    \I__11511\ : CascadeMux
    port map (
            O => \N__45989\,
            I => \N__45874\
        );

    \I__11510\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45866\
        );

    \I__11509\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45866\
        );

    \I__11508\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45866\
        );

    \I__11507\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45857\
        );

    \I__11506\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45857\
        );

    \I__11505\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45857\
        );

    \I__11504\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45857\
        );

    \I__11503\ : InMux
    port map (
            O => \N__45967\,
            I => \N__45854\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__45962\,
            I => \N__45843\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__45953\,
            I => \N__45843\
        );

    \I__11500\ : Span4Mux_h
    port map (
            O => \N__45950\,
            I => \N__45843\
        );

    \I__11499\ : Span4Mux_v
    port map (
            O => \N__45947\,
            I => \N__45843\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__45940\,
            I => \N__45843\
        );

    \I__11497\ : Span4Mux_h
    port map (
            O => \N__45937\,
            I => \N__45837\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__45934\,
            I => \N__45837\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__45931\,
            I => \N__45833\
        );

    \I__11494\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45830\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__45927\,
            I => \N__45825\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__45924\,
            I => \N__45825\
        );

    \I__11491\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45822\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__45920\,
            I => \N__45819\
        );

    \I__11489\ : Span4Mux_h
    port map (
            O => \N__45913\,
            I => \N__45816\
        );

    \I__11488\ : Span4Mux_v
    port map (
            O => \N__45910\,
            I => \N__45813\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__45907\,
            I => \N__45808\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__45904\,
            I => \N__45808\
        );

    \I__11485\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45805\
        );

    \I__11484\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45798\
        );

    \I__11483\ : InMux
    port map (
            O => \N__45897\,
            I => \N__45798\
        );

    \I__11482\ : InMux
    port map (
            O => \N__45894\,
            I => \N__45798\
        );

    \I__11481\ : InMux
    port map (
            O => \N__45893\,
            I => \N__45795\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__45886\,
            I => \N__45790\
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__45883\,
            I => \N__45790\
        );

    \I__11478\ : InMux
    port map (
            O => \N__45880\,
            I => \N__45787\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__45877\,
            I => \N__45784\
        );

    \I__11476\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45781\
        );

    \I__11475\ : CascadeMux
    port map (
            O => \N__45873\,
            I => \N__45778\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__45866\,
            I => \N__45769\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__45857\,
            I => \N__45769\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__45854\,
            I => \N__45769\
        );

    \I__11471\ : Span4Mux_v
    port map (
            O => \N__45843\,
            I => \N__45769\
        );

    \I__11470\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45766\
        );

    \I__11469\ : Span4Mux_v
    port map (
            O => \N__45837\,
            I => \N__45763\
        );

    \I__11468\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45760\
        );

    \I__11467\ : Span4Mux_h
    port map (
            O => \N__45833\,
            I => \N__45751\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45751\
        );

    \I__11465\ : Span4Mux_v
    port map (
            O => \N__45825\,
            I => \N__45751\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__45822\,
            I => \N__45751\
        );

    \I__11463\ : Span4Mux_v
    port map (
            O => \N__45819\,
            I => \N__45748\
        );

    \I__11462\ : Span4Mux_h
    port map (
            O => \N__45816\,
            I => \N__45741\
        );

    \I__11461\ : Span4Mux_h
    port map (
            O => \N__45813\,
            I => \N__45741\
        );

    \I__11460\ : Span4Mux_v
    port map (
            O => \N__45808\,
            I => \N__45741\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__45805\,
            I => \N__45734\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__45798\,
            I => \N__45734\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45734\
        );

    \I__11456\ : Span4Mux_h
    port map (
            O => \N__45790\,
            I => \N__45731\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__45787\,
            I => \N__45724\
        );

    \I__11454\ : Span4Mux_h
    port map (
            O => \N__45784\,
            I => \N__45724\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__45781\,
            I => \N__45724\
        );

    \I__11452\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45721\
        );

    \I__11451\ : Span4Mux_h
    port map (
            O => \N__45769\,
            I => \N__45718\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__45766\,
            I => \N__45713\
        );

    \I__11449\ : Span4Mux_h
    port map (
            O => \N__45763\,
            I => \N__45713\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__45760\,
            I => \N__45710\
        );

    \I__11447\ : Span4Mux_v
    port map (
            O => \N__45751\,
            I => \N__45705\
        );

    \I__11446\ : Span4Mux_v
    port map (
            O => \N__45748\,
            I => \N__45705\
        );

    \I__11445\ : Span4Mux_v
    port map (
            O => \N__45741\,
            I => \N__45700\
        );

    \I__11444\ : Span4Mux_v
    port map (
            O => \N__45734\,
            I => \N__45700\
        );

    \I__11443\ : Span4Mux_v
    port map (
            O => \N__45731\,
            I => \N__45692\
        );

    \I__11442\ : Span4Mux_v
    port map (
            O => \N__45724\,
            I => \N__45692\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__45721\,
            I => \N__45685\
        );

    \I__11440\ : Span4Mux_h
    port map (
            O => \N__45718\,
            I => \N__45685\
        );

    \I__11439\ : Span4Mux_v
    port map (
            O => \N__45713\,
            I => \N__45685\
        );

    \I__11438\ : Span4Mux_v
    port map (
            O => \N__45710\,
            I => \N__45680\
        );

    \I__11437\ : Span4Mux_h
    port map (
            O => \N__45705\,
            I => \N__45680\
        );

    \I__11436\ : Span4Mux_v
    port map (
            O => \N__45700\,
            I => \N__45677\
        );

    \I__11435\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45674\
        );

    \I__11434\ : InMux
    port map (
            O => \N__45698\,
            I => \N__45671\
        );

    \I__11433\ : InMux
    port map (
            O => \N__45697\,
            I => \N__45668\
        );

    \I__11432\ : Span4Mux_h
    port map (
            O => \N__45692\,
            I => \N__45665\
        );

    \I__11431\ : Span4Mux_v
    port map (
            O => \N__45685\,
            I => \N__45662\
        );

    \I__11430\ : Span4Mux_h
    port map (
            O => \N__45680\,
            I => \N__45659\
        );

    \I__11429\ : Span4Mux_h
    port map (
            O => \N__45677\,
            I => \N__45656\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__45674\,
            I => \N__45653\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__45671\,
            I => \aluOperation_1\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__45668\,
            I => \aluOperation_1\
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__45665\,
            I => \aluOperation_1\
        );

    \I__11424\ : Odrv4
    port map (
            O => \N__45662\,
            I => \aluOperation_1\
        );

    \I__11423\ : Odrv4
    port map (
            O => \N__45659\,
            I => \aluOperation_1\
        );

    \I__11422\ : Odrv4
    port map (
            O => \N__45656\,
            I => \aluOperation_1\
        );

    \I__11421\ : Odrv4
    port map (
            O => \N__45653\,
            I => \aluOperation_1\
        );

    \I__11420\ : CascadeMux
    port map (
            O => \N__45638\,
            I => \ALU.a_15_m5_6_cascade_\
        );

    \I__11419\ : InMux
    port map (
            O => \N__45635\,
            I => \N__45632\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__45632\,
            I => \N__45629\
        );

    \I__11417\ : Odrv12
    port map (
            O => \N__45629\,
            I => \ALU.mult_6\
        );

    \I__11416\ : CascadeMux
    port map (
            O => \N__45626\,
            I => \ALU.d_RNILPR7TQZ0Z_6_cascade_\
        );

    \I__11415\ : InMux
    port map (
            O => \N__45623\,
            I => \N__45619\
        );

    \I__11414\ : CascadeMux
    port map (
            O => \N__45622\,
            I => \N__45616\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__45619\,
            I => \N__45613\
        );

    \I__11412\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45610\
        );

    \I__11411\ : Span4Mux_h
    port map (
            O => \N__45613\,
            I => \N__45607\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45604\
        );

    \I__11409\ : Span4Mux_h
    port map (
            O => \N__45607\,
            I => \N__45601\
        );

    \I__11408\ : Span4Mux_v
    port map (
            O => \N__45604\,
            I => \N__45598\
        );

    \I__11407\ : Span4Mux_v
    port map (
            O => \N__45601\,
            I => \N__45595\
        );

    \I__11406\ : Span4Mux_h
    port map (
            O => \N__45598\,
            I => \N__45592\
        );

    \I__11405\ : Odrv4
    port map (
            O => \N__45595\,
            I => \ALU.hZ0Z_6\
        );

    \I__11404\ : Odrv4
    port map (
            O => \N__45592\,
            I => \ALU.hZ0Z_6\
        );

    \I__11403\ : CEMux
    port map (
            O => \N__45587\,
            I => \N__45583\
        );

    \I__11402\ : CEMux
    port map (
            O => \N__45586\,
            I => \N__45580\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__45583\,
            I => \N__45575\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__45580\,
            I => \N__45575\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__45575\,
            I => \N__45569\
        );

    \I__11398\ : CEMux
    port map (
            O => \N__45574\,
            I => \N__45564\
        );

    \I__11397\ : CEMux
    port map (
            O => \N__45573\,
            I => \N__45561\
        );

    \I__11396\ : CEMux
    port map (
            O => \N__45572\,
            I => \N__45558\
        );

    \I__11395\ : Span4Mux_h
    port map (
            O => \N__45569\,
            I => \N__45554\
        );

    \I__11394\ : CEMux
    port map (
            O => \N__45568\,
            I => \N__45551\
        );

    \I__11393\ : CEMux
    port map (
            O => \N__45567\,
            I => \N__45548\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__45564\,
            I => \N__45545\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__45561\,
            I => \N__45542\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__45558\,
            I => \N__45539\
        );

    \I__11389\ : CEMux
    port map (
            O => \N__45557\,
            I => \N__45535\
        );

    \I__11388\ : Span4Mux_v
    port map (
            O => \N__45554\,
            I => \N__45532\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__45551\,
            I => \N__45529\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__45548\,
            I => \N__45526\
        );

    \I__11385\ : Span4Mux_h
    port map (
            O => \N__45545\,
            I => \N__45522\
        );

    \I__11384\ : Span4Mux_v
    port map (
            O => \N__45542\,
            I => \N__45517\
        );

    \I__11383\ : Span4Mux_h
    port map (
            O => \N__45539\,
            I => \N__45517\
        );

    \I__11382\ : CEMux
    port map (
            O => \N__45538\,
            I => \N__45514\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45511\
        );

    \I__11380\ : Span4Mux_v
    port map (
            O => \N__45532\,
            I => \N__45508\
        );

    \I__11379\ : Span4Mux_h
    port map (
            O => \N__45529\,
            I => \N__45505\
        );

    \I__11378\ : Span4Mux_v
    port map (
            O => \N__45526\,
            I => \N__45502\
        );

    \I__11377\ : CEMux
    port map (
            O => \N__45525\,
            I => \N__45499\
        );

    \I__11376\ : Span4Mux_v
    port map (
            O => \N__45522\,
            I => \N__45495\
        );

    \I__11375\ : Span4Mux_v
    port map (
            O => \N__45517\,
            I => \N__45490\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__45514\,
            I => \N__45490\
        );

    \I__11373\ : Span4Mux_v
    port map (
            O => \N__45511\,
            I => \N__45486\
        );

    \I__11372\ : IoSpan4Mux
    port map (
            O => \N__45508\,
            I => \N__45483\
        );

    \I__11371\ : Span4Mux_v
    port map (
            O => \N__45505\,
            I => \N__45476\
        );

    \I__11370\ : Span4Mux_h
    port map (
            O => \N__45502\,
            I => \N__45476\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__45499\,
            I => \N__45476\
        );

    \I__11368\ : CEMux
    port map (
            O => \N__45498\,
            I => \N__45473\
        );

    \I__11367\ : Span4Mux_v
    port map (
            O => \N__45495\,
            I => \N__45468\
        );

    \I__11366\ : Span4Mux_h
    port map (
            O => \N__45490\,
            I => \N__45468\
        );

    \I__11365\ : CEMux
    port map (
            O => \N__45489\,
            I => \N__45465\
        );

    \I__11364\ : Span4Mux_v
    port map (
            O => \N__45486\,
            I => \N__45462\
        );

    \I__11363\ : Span4Mux_s2_v
    port map (
            O => \N__45483\,
            I => \N__45459\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__45476\,
            I => \N__45456\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__45473\,
            I => \N__45453\
        );

    \I__11360\ : Span4Mux_h
    port map (
            O => \N__45468\,
            I => \N__45450\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__45465\,
            I => \N__45447\
        );

    \I__11358\ : Span4Mux_h
    port map (
            O => \N__45462\,
            I => \N__45444\
        );

    \I__11357\ : Span4Mux_s2_h
    port map (
            O => \N__45459\,
            I => \N__45439\
        );

    \I__11356\ : Span4Mux_v
    port map (
            O => \N__45456\,
            I => \N__45439\
        );

    \I__11355\ : Span4Mux_v
    port map (
            O => \N__45453\,
            I => \N__45436\
        );

    \I__11354\ : Span4Mux_s3_h
    port map (
            O => \N__45450\,
            I => \N__45431\
        );

    \I__11353\ : Span4Mux_h
    port map (
            O => \N__45447\,
            I => \N__45431\
        );

    \I__11352\ : Span4Mux_h
    port map (
            O => \N__45444\,
            I => \N__45428\
        );

    \I__11351\ : Span4Mux_h
    port map (
            O => \N__45439\,
            I => \N__45425\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__45436\,
            I => \N__45422\
        );

    \I__11349\ : Span4Mux_v
    port map (
            O => \N__45431\,
            I => \N__45419\
        );

    \I__11348\ : Odrv4
    port map (
            O => \N__45428\,
            I => \ALU.h_cnvZ0Z_0\
        );

    \I__11347\ : Odrv4
    port map (
            O => \N__45425\,
            I => \ALU.h_cnvZ0Z_0\
        );

    \I__11346\ : Odrv4
    port map (
            O => \N__45422\,
            I => \ALU.h_cnvZ0Z_0\
        );

    \I__11345\ : Odrv4
    port map (
            O => \N__45419\,
            I => \ALU.h_cnvZ0Z_0\
        );

    \I__11344\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45406\
        );

    \I__11343\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45403\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__45406\,
            I => \N__45400\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__45403\,
            I => \N__45397\
        );

    \I__11340\ : Span4Mux_h
    port map (
            O => \N__45400\,
            I => \N__45392\
        );

    \I__11339\ : Span4Mux_h
    port map (
            O => \N__45397\,
            I => \N__45392\
        );

    \I__11338\ : Odrv4
    port map (
            O => \N__45392\,
            I => \ALU.fZ0Z_4\
        );

    \I__11337\ : InMux
    port map (
            O => \N__45389\,
            I => \N__45386\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__45386\,
            I => \N__45383\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__45383\,
            I => \N__45380\
        );

    \I__11334\ : Span4Mux_h
    port map (
            O => \N__45380\,
            I => \N__45377\
        );

    \I__11333\ : Odrv4
    port map (
            O => \N__45377\,
            I => \ALU.f_RNIJ0FJZ0Z_4\
        );

    \I__11332\ : InMux
    port map (
            O => \N__45374\,
            I => \N__45370\
        );

    \I__11331\ : InMux
    port map (
            O => \N__45373\,
            I => \N__45367\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__45370\,
            I => \N__45364\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__45367\,
            I => \N__45359\
        );

    \I__11328\ : Span12Mux_v
    port map (
            O => \N__45364\,
            I => \N__45359\
        );

    \I__11327\ : Odrv12
    port map (
            O => \N__45359\,
            I => \ALU.hZ0Z_7\
        );

    \I__11326\ : InMux
    port map (
            O => \N__45356\,
            I => \N__45353\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__45353\,
            I => \N__45350\
        );

    \I__11324\ : Span12Mux_s9_h
    port map (
            O => \N__45350\,
            I => \N__45346\
        );

    \I__11323\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45343\
        );

    \I__11322\ : Odrv12
    port map (
            O => \N__45346\,
            I => \ALU.dZ0Z_7\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__45343\,
            I => \ALU.dZ0Z_7\
        );

    \I__11320\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45330\
        );

    \I__11319\ : InMux
    port map (
            O => \N__45337\,
            I => \N__45323\
        );

    \I__11318\ : InMux
    port map (
            O => \N__45336\,
            I => \N__45323\
        );

    \I__11317\ : InMux
    port map (
            O => \N__45335\,
            I => \N__45323\
        );

    \I__11316\ : InMux
    port map (
            O => \N__45334\,
            I => \N__45318\
        );

    \I__11315\ : InMux
    port map (
            O => \N__45333\,
            I => \N__45315\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__45330\,
            I => \N__45309\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__45323\,
            I => \N__45306\
        );

    \I__11312\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45303\
        );

    \I__11311\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45300\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__45318\,
            I => \N__45296\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__45315\,
            I => \N__45293\
        );

    \I__11308\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45288\
        );

    \I__11307\ : InMux
    port map (
            O => \N__45313\,
            I => \N__45288\
        );

    \I__11306\ : InMux
    port map (
            O => \N__45312\,
            I => \N__45285\
        );

    \I__11305\ : Span4Mux_v
    port map (
            O => \N__45309\,
            I => \N__45270\
        );

    \I__11304\ : Span4Mux_v
    port map (
            O => \N__45306\,
            I => \N__45270\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__45303\,
            I => \N__45265\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__45300\,
            I => \N__45265\
        );

    \I__11301\ : InMux
    port map (
            O => \N__45299\,
            I => \N__45262\
        );

    \I__11300\ : Span4Mux_h
    port map (
            O => \N__45296\,
            I => \N__45255\
        );

    \I__11299\ : Span4Mux_v
    port map (
            O => \N__45293\,
            I => \N__45255\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__45288\,
            I => \N__45255\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__45285\,
            I => \N__45252\
        );

    \I__11296\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45247\
        );

    \I__11295\ : InMux
    port map (
            O => \N__45283\,
            I => \N__45247\
        );

    \I__11294\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45242\
        );

    \I__11293\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45242\
        );

    \I__11292\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45231\
        );

    \I__11291\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45231\
        );

    \I__11290\ : InMux
    port map (
            O => \N__45278\,
            I => \N__45231\
        );

    \I__11289\ : InMux
    port map (
            O => \N__45277\,
            I => \N__45231\
        );

    \I__11288\ : InMux
    port map (
            O => \N__45276\,
            I => \N__45231\
        );

    \I__11287\ : InMux
    port map (
            O => \N__45275\,
            I => \N__45228\
        );

    \I__11286\ : Span4Mux_v
    port map (
            O => \N__45270\,
            I => \N__45223\
        );

    \I__11285\ : Span4Mux_v
    port map (
            O => \N__45265\,
            I => \N__45223\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__45262\,
            I => \N__45216\
        );

    \I__11283\ : Span4Mux_v
    port map (
            O => \N__45255\,
            I => \N__45216\
        );

    \I__11282\ : Span4Mux_v
    port map (
            O => \N__45252\,
            I => \N__45216\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__45247\,
            I => \aluOperand2_2\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__45242\,
            I => \aluOperand2_2\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__45231\,
            I => \aluOperand2_2\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__45228\,
            I => \aluOperand2_2\
        );

    \I__11277\ : Odrv4
    port map (
            O => \N__45223\,
            I => \aluOperand2_2\
        );

    \I__11276\ : Odrv4
    port map (
            O => \N__45216\,
            I => \aluOperand2_2\
        );

    \I__11275\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45200\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__45200\,
            I => \N__45197\
        );

    \I__11273\ : Span4Mux_h
    port map (
            O => \N__45197\,
            I => \N__45194\
        );

    \I__11272\ : Span4Mux_h
    port map (
            O => \N__45194\,
            I => \N__45191\
        );

    \I__11271\ : Span4Mux_h
    port map (
            O => \N__45191\,
            I => \N__45188\
        );

    \I__11270\ : Odrv4
    port map (
            O => \N__45188\,
            I => \ALU.d_RNIU60LZ0Z_7\
        );

    \I__11269\ : CascadeMux
    port map (
            O => \N__45185\,
            I => \N__45182\
        );

    \I__11268\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45179\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__45179\,
            I => \N__45176\
        );

    \I__11266\ : Span4Mux_h
    port map (
            O => \N__45176\,
            I => \N__45172\
        );

    \I__11265\ : InMux
    port map (
            O => \N__45175\,
            I => \N__45169\
        );

    \I__11264\ : Span4Mux_h
    port map (
            O => \N__45172\,
            I => \N__45166\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__45169\,
            I => \N__45163\
        );

    \I__11262\ : Odrv4
    port map (
            O => \N__45166\,
            I => \ALU.hZ0Z_3\
        );

    \I__11261\ : Odrv4
    port map (
            O => \N__45163\,
            I => \ALU.hZ0Z_3\
        );

    \I__11260\ : InMux
    port map (
            O => \N__45158\,
            I => \N__45155\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__45155\,
            I => \N__45152\
        );

    \I__11258\ : Span4Mux_v
    port map (
            O => \N__45152\,
            I => \N__45149\
        );

    \I__11257\ : Span4Mux_h
    port map (
            O => \N__45149\,
            I => \N__45145\
        );

    \I__11256\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45142\
        );

    \I__11255\ : Odrv4
    port map (
            O => \N__45145\,
            I => \ALU.dZ0Z_3\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__45142\,
            I => \ALU.dZ0Z_3\
        );

    \I__11253\ : InMux
    port map (
            O => \N__45137\,
            I => \N__45130\
        );

    \I__11252\ : InMux
    port map (
            O => \N__45136\,
            I => \N__45130\
        );

    \I__11251\ : CascadeMux
    port map (
            O => \N__45135\,
            I => \N__45123\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__45130\,
            I => \N__45116\
        );

    \I__11249\ : InMux
    port map (
            O => \N__45129\,
            I => \N__45113\
        );

    \I__11248\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45109\
        );

    \I__11247\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45104\
        );

    \I__11246\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45104\
        );

    \I__11245\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45100\
        );

    \I__11244\ : InMux
    port map (
            O => \N__45122\,
            I => \N__45097\
        );

    \I__11243\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45094\
        );

    \I__11242\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45091\
        );

    \I__11241\ : InMux
    port map (
            O => \N__45119\,
            I => \N__45088\
        );

    \I__11240\ : Span4Mux_v
    port map (
            O => \N__45116\,
            I => \N__45085\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45082\
        );

    \I__11238\ : InMux
    port map (
            O => \N__45112\,
            I => \N__45073\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__45109\,
            I => \N__45070\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__45104\,
            I => \N__45067\
        );

    \I__11235\ : InMux
    port map (
            O => \N__45103\,
            I => \N__45064\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__45100\,
            I => \N__45060\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__45097\,
            I => \N__45057\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__45094\,
            I => \N__45050\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__45091\,
            I => \N__45050\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__45088\,
            I => \N__45050\
        );

    \I__11229\ : Span4Mux_s3_h
    port map (
            O => \N__45085\,
            I => \N__45047\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__45082\,
            I => \N__45044\
        );

    \I__11227\ : InMux
    port map (
            O => \N__45081\,
            I => \N__45041\
        );

    \I__11226\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45030\
        );

    \I__11225\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45030\
        );

    \I__11224\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45030\
        );

    \I__11223\ : InMux
    port map (
            O => \N__45077\,
            I => \N__45030\
        );

    \I__11222\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45030\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__45073\,
            I => \N__45027\
        );

    \I__11220\ : Span4Mux_v
    port map (
            O => \N__45070\,
            I => \N__45022\
        );

    \I__11219\ : Span4Mux_h
    port map (
            O => \N__45067\,
            I => \N__45022\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__45064\,
            I => \N__45019\
        );

    \I__11217\ : InMux
    port map (
            O => \N__45063\,
            I => \N__45016\
        );

    \I__11216\ : Span4Mux_v
    port map (
            O => \N__45060\,
            I => \N__45009\
        );

    \I__11215\ : Span4Mux_v
    port map (
            O => \N__45057\,
            I => \N__45009\
        );

    \I__11214\ : Span4Mux_v
    port map (
            O => \N__45050\,
            I => \N__45009\
        );

    \I__11213\ : Span4Mux_h
    port map (
            O => \N__45047\,
            I => \N__45004\
        );

    \I__11212\ : Span4Mux_v
    port map (
            O => \N__45044\,
            I => \N__45004\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__45041\,
            I => \aluOperand2_2_rep2\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__45030\,
            I => \aluOperand2_2_rep2\
        );

    \I__11209\ : Odrv4
    port map (
            O => \N__45027\,
            I => \aluOperand2_2_rep2\
        );

    \I__11208\ : Odrv4
    port map (
            O => \N__45022\,
            I => \aluOperand2_2_rep2\
        );

    \I__11207\ : Odrv4
    port map (
            O => \N__45019\,
            I => \aluOperand2_2_rep2\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__45016\,
            I => \aluOperand2_2_rep2\
        );

    \I__11205\ : Odrv4
    port map (
            O => \N__45009\,
            I => \aluOperand2_2_rep2\
        );

    \I__11204\ : Odrv4
    port map (
            O => \N__45004\,
            I => \aluOperand2_2_rep2\
        );

    \I__11203\ : InMux
    port map (
            O => \N__44987\,
            I => \N__44984\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__44984\,
            I => \N__44981\
        );

    \I__11201\ : Span4Mux_h
    port map (
            O => \N__44981\,
            I => \N__44978\
        );

    \I__11200\ : Span4Mux_h
    port map (
            O => \N__44978\,
            I => \N__44975\
        );

    \I__11199\ : Odrv4
    port map (
            O => \N__44975\,
            I => \ALU.d_RNILAR7Z0Z_3\
        );

    \I__11198\ : CascadeMux
    port map (
            O => \N__44972\,
            I => \ALU.a_15_m2_4_cascade_\
        );

    \I__11197\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44966\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__44966\,
            I => \N__44963\
        );

    \I__11195\ : Span4Mux_v
    port map (
            O => \N__44963\,
            I => \N__44960\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__44960\,
            I => \N__44956\
        );

    \I__11193\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44953\
        );

    \I__11192\ : Span4Mux_h
    port map (
            O => \N__44956\,
            I => \N__44950\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44947\
        );

    \I__11190\ : Odrv4
    port map (
            O => \N__44950\,
            I => \ALU.N_419\
        );

    \I__11189\ : Odrv4
    port map (
            O => \N__44947\,
            I => \ALU.N_419\
        );

    \I__11188\ : InMux
    port map (
            O => \N__44942\,
            I => \N__44939\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__44939\,
            I => \ALU.a_15_m4_4\
        );

    \I__11186\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44933\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__44933\,
            I => \N__44930\
        );

    \I__11184\ : Sp12to4
    port map (
            O => \N__44930\,
            I => \N__44927\
        );

    \I__11183\ : Span12Mux_v
    port map (
            O => \N__44927\,
            I => \N__44924\
        );

    \I__11182\ : Odrv12
    port map (
            O => \N__44924\,
            I => \ALU.mult_4\
        );

    \I__11181\ : InMux
    port map (
            O => \N__44921\,
            I => \N__44918\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__44918\,
            I => \ALU.a_15_m5_4\
        );

    \I__11179\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44912\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__44912\,
            I => \N__44909\
        );

    \I__11177\ : Span4Mux_h
    port map (
            O => \N__44909\,
            I => \N__44904\
        );

    \I__11176\ : InMux
    port map (
            O => \N__44908\,
            I => \N__44899\
        );

    \I__11175\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44899\
        );

    \I__11174\ : Sp12to4
    port map (
            O => \N__44904\,
            I => \N__44896\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44893\
        );

    \I__11172\ : Odrv12
    port map (
            O => \N__44896\,
            I => a_3
        );

    \I__11171\ : Odrv12
    port map (
            O => \N__44893\,
            I => a_3
        );

    \I__11170\ : CEMux
    port map (
            O => \N__44888\,
            I => \N__44885\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__44885\,
            I => \N__44881\
        );

    \I__11168\ : CEMux
    port map (
            O => \N__44884\,
            I => \N__44878\
        );

    \I__11167\ : Span4Mux_h
    port map (
            O => \N__44881\,
            I => \N__44873\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__44878\,
            I => \N__44873\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__44873\,
            I => \N__44867\
        );

    \I__11164\ : CEMux
    port map (
            O => \N__44872\,
            I => \N__44864\
        );

    \I__11163\ : CEMux
    port map (
            O => \N__44871\,
            I => \N__44861\
        );

    \I__11162\ : CEMux
    port map (
            O => \N__44870\,
            I => \N__44858\
        );

    \I__11161\ : Span4Mux_v
    port map (
            O => \N__44867\,
            I => \N__44853\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__44864\,
            I => \N__44853\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__44861\,
            I => \N__44850\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__44858\,
            I => \N__44846\
        );

    \I__11157\ : Span4Mux_v
    port map (
            O => \N__44853\,
            I => \N__44841\
        );

    \I__11156\ : Span4Mux_v
    port map (
            O => \N__44850\,
            I => \N__44841\
        );

    \I__11155\ : CEMux
    port map (
            O => \N__44849\,
            I => \N__44838\
        );

    \I__11154\ : Span4Mux_h
    port map (
            O => \N__44846\,
            I => \N__44834\
        );

    \I__11153\ : IoSpan4Mux
    port map (
            O => \N__44841\,
            I => \N__44831\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__44838\,
            I => \N__44828\
        );

    \I__11151\ : CEMux
    port map (
            O => \N__44837\,
            I => \N__44825\
        );

    \I__11150\ : Sp12to4
    port map (
            O => \N__44834\,
            I => \N__44822\
        );

    \I__11149\ : IoSpan4Mux
    port map (
            O => \N__44831\,
            I => \N__44819\
        );

    \I__11148\ : Span4Mux_h
    port map (
            O => \N__44828\,
            I => \N__44816\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__44825\,
            I => \N__44813\
        );

    \I__11146\ : Span12Mux_s8_h
    port map (
            O => \N__44822\,
            I => \N__44810\
        );

    \I__11145\ : Span4Mux_s0_v
    port map (
            O => \N__44819\,
            I => \N__44807\
        );

    \I__11144\ : Span4Mux_h
    port map (
            O => \N__44816\,
            I => \N__44804\
        );

    \I__11143\ : Span4Mux_v
    port map (
            O => \N__44813\,
            I => \N__44801\
        );

    \I__11142\ : Span12Mux_v
    port map (
            O => \N__44810\,
            I => \N__44798\
        );

    \I__11141\ : Span4Mux_h
    port map (
            O => \N__44807\,
            I => \N__44795\
        );

    \I__11140\ : Span4Mux_v
    port map (
            O => \N__44804\,
            I => \N__44792\
        );

    \I__11139\ : Span4Mux_v
    port map (
            O => \N__44801\,
            I => \N__44789\
        );

    \I__11138\ : Odrv12
    port map (
            O => \N__44798\,
            I => \ALU.a_cnvZ0Z_0\
        );

    \I__11137\ : Odrv4
    port map (
            O => \N__44795\,
            I => \ALU.a_cnvZ0Z_0\
        );

    \I__11136\ : Odrv4
    port map (
            O => \N__44792\,
            I => \ALU.a_cnvZ0Z_0\
        );

    \I__11135\ : Odrv4
    port map (
            O => \N__44789\,
            I => \ALU.a_cnvZ0Z_0\
        );

    \I__11134\ : InMux
    port map (
            O => \N__44780\,
            I => \N__44777\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__44777\,
            I => \N__44774\
        );

    \I__11132\ : Odrv4
    port map (
            O => \N__44774\,
            I => \FTDI.TXshiftZ0Z_2\
        );

    \I__11131\ : InMux
    port map (
            O => \N__44771\,
            I => \N__44763\
        );

    \I__11130\ : InMux
    port map (
            O => \N__44770\,
            I => \N__44763\
        );

    \I__11129\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44760\
        );

    \I__11128\ : CascadeMux
    port map (
            O => \N__44768\,
            I => \N__44750\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__44763\,
            I => \N__44745\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44741\
        );

    \I__11125\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44726\
        );

    \I__11124\ : InMux
    port map (
            O => \N__44758\,
            I => \N__44726\
        );

    \I__11123\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44726\
        );

    \I__11122\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44726\
        );

    \I__11121\ : InMux
    port map (
            O => \N__44755\,
            I => \N__44726\
        );

    \I__11120\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44726\
        );

    \I__11119\ : InMux
    port map (
            O => \N__44753\,
            I => \N__44726\
        );

    \I__11118\ : InMux
    port map (
            O => \N__44750\,
            I => \N__44723\
        );

    \I__11117\ : CascadeMux
    port map (
            O => \N__44749\,
            I => \N__44720\
        );

    \I__11116\ : CascadeMux
    port map (
            O => \N__44748\,
            I => \N__44714\
        );

    \I__11115\ : Span4Mux_s2_v
    port map (
            O => \N__44745\,
            I => \N__44711\
        );

    \I__11114\ : InMux
    port map (
            O => \N__44744\,
            I => \N__44708\
        );

    \I__11113\ : Span4Mux_h
    port map (
            O => \N__44741\,
            I => \N__44701\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__44726\,
            I => \N__44701\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__44723\,
            I => \N__44701\
        );

    \I__11110\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44698\
        );

    \I__11109\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44693\
        );

    \I__11108\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44693\
        );

    \I__11107\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44688\
        );

    \I__11106\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44688\
        );

    \I__11105\ : Odrv4
    port map (
            O => \N__44711\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__44708\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__11103\ : Odrv4
    port map (
            O => \N__44701\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__44698\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__44693\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__44688\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__11099\ : InMux
    port map (
            O => \N__44675\,
            I => \N__44672\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__44672\,
            I => \N__44669\
        );

    \I__11097\ : Odrv4
    port map (
            O => \N__44669\,
            I => \FTDI.TXshiftZ0Z_1\
        );

    \I__11096\ : CEMux
    port map (
            O => \N__44666\,
            I => \N__44663\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__44663\,
            I => \N__44660\
        );

    \I__11094\ : Span4Mux_h
    port map (
            O => \N__44660\,
            I => \N__44656\
        );

    \I__11093\ : CEMux
    port map (
            O => \N__44659\,
            I => \N__44653\
        );

    \I__11092\ : Sp12to4
    port map (
            O => \N__44656\,
            I => \N__44648\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__44653\,
            I => \N__44648\
        );

    \I__11090\ : Odrv12
    port map (
            O => \N__44648\,
            I => \FTDI.un1_TXstate_0_sqmuxa_0_i\
        );

    \I__11089\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44642\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__44642\,
            I => \N__44638\
        );

    \I__11087\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44635\
        );

    \I__11086\ : Span4Mux_v
    port map (
            O => \N__44638\,
            I => \N__44632\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__44635\,
            I => \N__44629\
        );

    \I__11084\ : Span4Mux_h
    port map (
            O => \N__44632\,
            I => \N__44625\
        );

    \I__11083\ : Span4Mux_h
    port map (
            O => \N__44629\,
            I => \N__44622\
        );

    \I__11082\ : InMux
    port map (
            O => \N__44628\,
            I => \N__44619\
        );

    \I__11081\ : Odrv4
    port map (
            O => \N__44625\,
            I => a_5
        );

    \I__11080\ : Odrv4
    port map (
            O => \N__44622\,
            I => a_5
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__44619\,
            I => a_5
        );

    \I__11078\ : InMux
    port map (
            O => \N__44612\,
            I => \N__44609\
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__44609\,
            I => \N__44606\
        );

    \I__11076\ : Span4Mux_h
    port map (
            O => \N__44606\,
            I => \N__44603\
        );

    \I__11075\ : Odrv4
    port map (
            O => \N__44603\,
            I => \TXbufferZ0Z_5\
        );

    \I__11074\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44597\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__44597\,
            I => \N__44593\
        );

    \I__11072\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44590\
        );

    \I__11071\ : Span4Mux_v
    port map (
            O => \N__44593\,
            I => \N__44587\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__44590\,
            I => \N__44583\
        );

    \I__11069\ : Span4Mux_h
    port map (
            O => \N__44587\,
            I => \N__44580\
        );

    \I__11068\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44577\
        );

    \I__11067\ : Span4Mux_h
    port map (
            O => \N__44583\,
            I => \N__44574\
        );

    \I__11066\ : Odrv4
    port map (
            O => \N__44580\,
            I => a_1
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__44577\,
            I => a_1
        );

    \I__11064\ : Odrv4
    port map (
            O => \N__44574\,
            I => a_1
        );

    \I__11063\ : InMux
    port map (
            O => \N__44567\,
            I => \N__44564\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44561\
        );

    \I__11061\ : Odrv4
    port map (
            O => \N__44561\,
            I => \TXbufferZ0Z_1\
        );

    \I__11060\ : CEMux
    port map (
            O => \N__44558\,
            I => \N__44555\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__44555\,
            I => \N__44552\
        );

    \I__11058\ : Span4Mux_v
    port map (
            O => \N__44552\,
            I => \N__44548\
        );

    \I__11057\ : CEMux
    port map (
            O => \N__44551\,
            I => \N__44545\
        );

    \I__11056\ : Odrv4
    port map (
            O => \N__44548\,
            I => m326dup
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__44545\,
            I => m326dup
        );

    \I__11054\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44534\
        );

    \I__11053\ : InMux
    port map (
            O => \N__44539\,
            I => \N__44531\
        );

    \I__11052\ : CascadeMux
    port map (
            O => \N__44538\,
            I => \N__44528\
        );

    \I__11051\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44515\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__44534\,
            I => \N__44512\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__44531\,
            I => \N__44509\
        );

    \I__11048\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44506\
        );

    \I__11047\ : InMux
    port map (
            O => \N__44527\,
            I => \N__44501\
        );

    \I__11046\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44501\
        );

    \I__11045\ : CascadeMux
    port map (
            O => \N__44525\,
            I => \N__44496\
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__44524\,
            I => \N__44493\
        );

    \I__11043\ : CascadeMux
    port map (
            O => \N__44523\,
            I => \N__44488\
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__44522\,
            I => \N__44484\
        );

    \I__11041\ : CascadeMux
    port map (
            O => \N__44521\,
            I => \N__44481\
        );

    \I__11040\ : InMux
    port map (
            O => \N__44520\,
            I => \N__44476\
        );

    \I__11039\ : InMux
    port map (
            O => \N__44519\,
            I => \N__44471\
        );

    \I__11038\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44471\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__44515\,
            I => \N__44466\
        );

    \I__11036\ : Span4Mux_v
    port map (
            O => \N__44512\,
            I => \N__44466\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__44509\,
            I => \N__44459\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__44506\,
            I => \N__44459\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__44501\,
            I => \N__44459\
        );

    \I__11032\ : InMux
    port map (
            O => \N__44500\,
            I => \N__44456\
        );

    \I__11031\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44453\
        );

    \I__11030\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44450\
        );

    \I__11029\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44445\
        );

    \I__11028\ : CascadeMux
    port map (
            O => \N__44492\,
            I => \N__44439\
        );

    \I__11027\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44434\
        );

    \I__11026\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44431\
        );

    \I__11025\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44426\
        );

    \I__11024\ : InMux
    port map (
            O => \N__44484\,
            I => \N__44426\
        );

    \I__11023\ : InMux
    port map (
            O => \N__44481\,
            I => \N__44423\
        );

    \I__11022\ : InMux
    port map (
            O => \N__44480\,
            I => \N__44417\
        );

    \I__11021\ : InMux
    port map (
            O => \N__44479\,
            I => \N__44414\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__44476\,
            I => \N__44409\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__44471\,
            I => \N__44409\
        );

    \I__11018\ : Span4Mux_v
    port map (
            O => \N__44466\,
            I => \N__44404\
        );

    \I__11017\ : Span4Mux_v
    port map (
            O => \N__44459\,
            I => \N__44404\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__44456\,
            I => \N__44396\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__44453\,
            I => \N__44396\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__44450\,
            I => \N__44396\
        );

    \I__11013\ : CascadeMux
    port map (
            O => \N__44449\,
            I => \N__44390\
        );

    \I__11012\ : InMux
    port map (
            O => \N__44448\,
            I => \N__44387\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__44445\,
            I => \N__44384\
        );

    \I__11010\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44381\
        );

    \I__11009\ : InMux
    port map (
            O => \N__44443\,
            I => \N__44374\
        );

    \I__11008\ : InMux
    port map (
            O => \N__44442\,
            I => \N__44374\
        );

    \I__11007\ : InMux
    port map (
            O => \N__44439\,
            I => \N__44374\
        );

    \I__11006\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44371\
        );

    \I__11005\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44368\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__44434\,
            I => \N__44363\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__44431\,
            I => \N__44363\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__44426\,
            I => \N__44358\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__44423\,
            I => \N__44358\
        );

    \I__11000\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44355\
        );

    \I__10999\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44352\
        );

    \I__10998\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44349\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__44417\,
            I => \N__44346\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__44414\,
            I => \N__44341\
        );

    \I__10995\ : Span4Mux_v
    port map (
            O => \N__44409\,
            I => \N__44341\
        );

    \I__10994\ : Span4Mux_v
    port map (
            O => \N__44404\,
            I => \N__44338\
        );

    \I__10993\ : CascadeMux
    port map (
            O => \N__44403\,
            I => \N__44335\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__44396\,
            I => \N__44331\
        );

    \I__10991\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44326\
        );

    \I__10990\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44326\
        );

    \I__10989\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44318\
        );

    \I__10988\ : InMux
    port map (
            O => \N__44390\,
            I => \N__44318\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__44387\,
            I => \N__44315\
        );

    \I__10986\ : Span4Mux_s2_v
    port map (
            O => \N__44384\,
            I => \N__44306\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__44381\,
            I => \N__44306\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__44374\,
            I => \N__44306\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__44371\,
            I => \N__44306\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44303\
        );

    \I__10981\ : Span4Mux_v
    port map (
            O => \N__44363\,
            I => \N__44292\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__44358\,
            I => \N__44292\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__44355\,
            I => \N__44292\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__44352\,
            I => \N__44292\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__44349\,
            I => \N__44292\
        );

    \I__10976\ : Span4Mux_s2_v
    port map (
            O => \N__44346\,
            I => \N__44285\
        );

    \I__10975\ : Span4Mux_s2_v
    port map (
            O => \N__44341\,
            I => \N__44285\
        );

    \I__10974\ : Span4Mux_h
    port map (
            O => \N__44338\,
            I => \N__44285\
        );

    \I__10973\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44280\
        );

    \I__10972\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44280\
        );

    \I__10971\ : Sp12to4
    port map (
            O => \N__44331\,
            I => \N__44275\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__44326\,
            I => \N__44275\
        );

    \I__10969\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44270\
        );

    \I__10968\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44270\
        );

    \I__10967\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44267\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__44318\,
            I => \N__44260\
        );

    \I__10965\ : Span4Mux_v
    port map (
            O => \N__44315\,
            I => \N__44260\
        );

    \I__10964\ : Span4Mux_v
    port map (
            O => \N__44306\,
            I => \N__44260\
        );

    \I__10963\ : Span12Mux_v
    port map (
            O => \N__44303\,
            I => \N__44249\
        );

    \I__10962\ : Sp12to4
    port map (
            O => \N__44292\,
            I => \N__44249\
        );

    \I__10961\ : Sp12to4
    port map (
            O => \N__44285\,
            I => \N__44249\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__44280\,
            I => \N__44249\
        );

    \I__10959\ : Span12Mux_s2_v
    port map (
            O => \N__44275\,
            I => \N__44249\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__44270\,
            I => \aluParams_3\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__44267\,
            I => \aluParams_3\
        );

    \I__10956\ : Odrv4
    port map (
            O => \N__44260\,
            I => \aluParams_3\
        );

    \I__10955\ : Odrv12
    port map (
            O => \N__44249\,
            I => \aluParams_3\
        );

    \I__10954\ : InMux
    port map (
            O => \N__44240\,
            I => \N__44237\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__44237\,
            I => \N__44234\
        );

    \I__10952\ : Span4Mux_v
    port map (
            O => \N__44234\,
            I => \N__44231\
        );

    \I__10951\ : Odrv4
    port map (
            O => \N__44231\,
            I => \ALU.N_308\
        );

    \I__10950\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44220\
        );

    \I__10949\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44215\
        );

    \I__10948\ : InMux
    port map (
            O => \N__44226\,
            I => \N__44212\
        );

    \I__10947\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44207\
        );

    \I__10946\ : InMux
    port map (
            O => \N__44224\,
            I => \N__44207\
        );

    \I__10945\ : InMux
    port map (
            O => \N__44223\,
            I => \N__44199\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__44220\,
            I => \N__44195\
        );

    \I__10943\ : InMux
    port map (
            O => \N__44219\,
            I => \N__44192\
        );

    \I__10942\ : CascadeMux
    port map (
            O => \N__44218\,
            I => \N__44189\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__44215\,
            I => \N__44182\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__44212\,
            I => \N__44182\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__44207\,
            I => \N__44179\
        );

    \I__10938\ : InMux
    port map (
            O => \N__44206\,
            I => \N__44174\
        );

    \I__10937\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44174\
        );

    \I__10936\ : InMux
    port map (
            O => \N__44204\,
            I => \N__44169\
        );

    \I__10935\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44169\
        );

    \I__10934\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44166\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__44199\,
            I => \N__44163\
        );

    \I__10932\ : InMux
    port map (
            O => \N__44198\,
            I => \N__44160\
        );

    \I__10931\ : Span4Mux_v
    port map (
            O => \N__44195\,
            I => \N__44156\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__44192\,
            I => \N__44153\
        );

    \I__10929\ : InMux
    port map (
            O => \N__44189\,
            I => \N__44143\
        );

    \I__10928\ : InMux
    port map (
            O => \N__44188\,
            I => \N__44143\
        );

    \I__10927\ : InMux
    port map (
            O => \N__44187\,
            I => \N__44140\
        );

    \I__10926\ : Span4Mux_h
    port map (
            O => \N__44182\,
            I => \N__44134\
        );

    \I__10925\ : Span4Mux_v
    port map (
            O => \N__44179\,
            I => \N__44134\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__44174\,
            I => \N__44122\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__44169\,
            I => \N__44122\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__44166\,
            I => \N__44122\
        );

    \I__10921\ : Span4Mux_h
    port map (
            O => \N__44163\,
            I => \N__44122\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__44160\,
            I => \N__44122\
        );

    \I__10919\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44118\
        );

    \I__10918\ : Span4Mux_h
    port map (
            O => \N__44156\,
            I => \N__44113\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__44153\,
            I => \N__44113\
        );

    \I__10916\ : InMux
    port map (
            O => \N__44152\,
            I => \N__44108\
        );

    \I__10915\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44108\
        );

    \I__10914\ : InMux
    port map (
            O => \N__44150\,
            I => \N__44105\
        );

    \I__10913\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44100\
        );

    \I__10912\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44100\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__44143\,
            I => \N__44097\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__44140\,
            I => \N__44094\
        );

    \I__10909\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44091\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__44134\,
            I => \N__44086\
        );

    \I__10907\ : InMux
    port map (
            O => \N__44133\,
            I => \N__44083\
        );

    \I__10906\ : Span4Mux_v
    port map (
            O => \N__44122\,
            I => \N__44080\
        );

    \I__10905\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44077\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__44118\,
            I => \N__44074\
        );

    \I__10903\ : Span4Mux_v
    port map (
            O => \N__44113\,
            I => \N__44071\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44068\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__44105\,
            I => \N__44061\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__44100\,
            I => \N__44061\
        );

    \I__10899\ : Span4Mux_v
    port map (
            O => \N__44097\,
            I => \N__44061\
        );

    \I__10898\ : Span4Mux_v
    port map (
            O => \N__44094\,
            I => \N__44055\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44055\
        );

    \I__10896\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44050\
        );

    \I__10895\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44050\
        );

    \I__10894\ : Span4Mux_v
    port map (
            O => \N__44086\,
            I => \N__44047\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__44083\,
            I => \N__44044\
        );

    \I__10892\ : Span4Mux_h
    port map (
            O => \N__44080\,
            I => \N__44039\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__44077\,
            I => \N__44039\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__44074\,
            I => \N__44030\
        );

    \I__10889\ : Span4Mux_h
    port map (
            O => \N__44071\,
            I => \N__44030\
        );

    \I__10888\ : Span4Mux_v
    port map (
            O => \N__44068\,
            I => \N__44030\
        );

    \I__10887\ : Span4Mux_v
    port map (
            O => \N__44061\,
            I => \N__44025\
        );

    \I__10886\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44022\
        );

    \I__10885\ : Span4Mux_h
    port map (
            O => \N__44055\,
            I => \N__44013\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__44050\,
            I => \N__44013\
        );

    \I__10883\ : Span4Mux_h
    port map (
            O => \N__44047\,
            I => \N__44013\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__44044\,
            I => \N__44013\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__44039\,
            I => \N__44010\
        );

    \I__10880\ : InMux
    port map (
            O => \N__44038\,
            I => \N__44007\
        );

    \I__10879\ : InMux
    port map (
            O => \N__44037\,
            I => \N__44004\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__44030\,
            I => \N__44001\
        );

    \I__10877\ : InMux
    port map (
            O => \N__44029\,
            I => \N__43998\
        );

    \I__10876\ : InMux
    port map (
            O => \N__44028\,
            I => \N__43995\
        );

    \I__10875\ : Sp12to4
    port map (
            O => \N__44025\,
            I => \N__43992\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__44022\,
            I => \N__43987\
        );

    \I__10873\ : Span4Mux_v
    port map (
            O => \N__44013\,
            I => \N__43987\
        );

    \I__10872\ : Span4Mux_s0_v
    port map (
            O => \N__44010\,
            I => \N__43984\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__44007\,
            I => \aluOperation_2\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__44004\,
            I => \aluOperation_2\
        );

    \I__10869\ : Odrv4
    port map (
            O => \N__44001\,
            I => \aluOperation_2\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__43998\,
            I => \aluOperation_2\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__43995\,
            I => \aluOperation_2\
        );

    \I__10866\ : Odrv12
    port map (
            O => \N__43992\,
            I => \aluOperation_2\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__43987\,
            I => \aluOperation_2\
        );

    \I__10864\ : Odrv4
    port map (
            O => \N__43984\,
            I => \aluOperation_2\
        );

    \I__10863\ : CascadeMux
    port map (
            O => \N__43967\,
            I => \N__43964\
        );

    \I__10862\ : InMux
    port map (
            O => \N__43964\,
            I => \N__43959\
        );

    \I__10861\ : CascadeMux
    port map (
            O => \N__43963\,
            I => \N__43956\
        );

    \I__10860\ : CascadeMux
    port map (
            O => \N__43962\,
            I => \N__43953\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__43959\,
            I => \N__43949\
        );

    \I__10858\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43946\
        );

    \I__10857\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43943\
        );

    \I__10856\ : CascadeMux
    port map (
            O => \N__43952\,
            I => \N__43940\
        );

    \I__10855\ : Span4Mux_h
    port map (
            O => \N__43949\,
            I => \N__43934\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__43946\,
            I => \N__43930\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__43943\,
            I => \N__43926\
        );

    \I__10852\ : InMux
    port map (
            O => \N__43940\,
            I => \N__43923\
        );

    \I__10851\ : CascadeMux
    port map (
            O => \N__43939\,
            I => \N__43920\
        );

    \I__10850\ : CascadeMux
    port map (
            O => \N__43938\,
            I => \N__43916\
        );

    \I__10849\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43913\
        );

    \I__10848\ : Span4Mux_h
    port map (
            O => \N__43934\,
            I => \N__43910\
        );

    \I__10847\ : InMux
    port map (
            O => \N__43933\,
            I => \N__43907\
        );

    \I__10846\ : Span4Mux_v
    port map (
            O => \N__43930\,
            I => \N__43904\
        );

    \I__10845\ : CascadeMux
    port map (
            O => \N__43929\,
            I => \N__43901\
        );

    \I__10844\ : Span4Mux_h
    port map (
            O => \N__43926\,
            I => \N__43894\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__43923\,
            I => \N__43894\
        );

    \I__10842\ : InMux
    port map (
            O => \N__43920\,
            I => \N__43891\
        );

    \I__10841\ : CascadeMux
    port map (
            O => \N__43919\,
            I => \N__43888\
        );

    \I__10840\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43885\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__43913\,
            I => \N__43882\
        );

    \I__10838\ : Span4Mux_v
    port map (
            O => \N__43910\,
            I => \N__43876\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__43907\,
            I => \N__43876\
        );

    \I__10836\ : Span4Mux_v
    port map (
            O => \N__43904\,
            I => \N__43873\
        );

    \I__10835\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43870\
        );

    \I__10834\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43865\
        );

    \I__10833\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43865\
        );

    \I__10832\ : Span4Mux_h
    port map (
            O => \N__43894\,
            I => \N__43862\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__43891\,
            I => \N__43856\
        );

    \I__10830\ : InMux
    port map (
            O => \N__43888\,
            I => \N__43853\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__43885\,
            I => \N__43850\
        );

    \I__10828\ : Span4Mux_v
    port map (
            O => \N__43882\,
            I => \N__43847\
        );

    \I__10827\ : CascadeMux
    port map (
            O => \N__43881\,
            I => \N__43844\
        );

    \I__10826\ : Span4Mux_v
    port map (
            O => \N__43876\,
            I => \N__43841\
        );

    \I__10825\ : Span4Mux_v
    port map (
            O => \N__43873\,
            I => \N__43838\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43833\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__43865\,
            I => \N__43833\
        );

    \I__10822\ : Span4Mux_h
    port map (
            O => \N__43862\,
            I => \N__43830\
        );

    \I__10821\ : InMux
    port map (
            O => \N__43861\,
            I => \N__43825\
        );

    \I__10820\ : InMux
    port map (
            O => \N__43860\,
            I => \N__43825\
        );

    \I__10819\ : InMux
    port map (
            O => \N__43859\,
            I => \N__43822\
        );

    \I__10818\ : Span4Mux_v
    port map (
            O => \N__43856\,
            I => \N__43819\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__43853\,
            I => \N__43816\
        );

    \I__10816\ : Span4Mux_v
    port map (
            O => \N__43850\,
            I => \N__43811\
        );

    \I__10815\ : Span4Mux_h
    port map (
            O => \N__43847\,
            I => \N__43811\
        );

    \I__10814\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43808\
        );

    \I__10813\ : Span4Mux_v
    port map (
            O => \N__43841\,
            I => \N__43805\
        );

    \I__10812\ : Span4Mux_h
    port map (
            O => \N__43838\,
            I => \N__43800\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__43833\,
            I => \N__43800\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__43830\,
            I => \N__43795\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__43825\,
            I => \N__43795\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43792\
        );

    \I__10807\ : Span4Mux_h
    port map (
            O => \N__43819\,
            I => \N__43781\
        );

    \I__10806\ : Span4Mux_v
    port map (
            O => \N__43816\,
            I => \N__43781\
        );

    \I__10805\ : Span4Mux_v
    port map (
            O => \N__43811\,
            I => \N__43781\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__43808\,
            I => \N__43781\
        );

    \I__10803\ : Span4Mux_s1_v
    port map (
            O => \N__43805\,
            I => \N__43781\
        );

    \I__10802\ : Span4Mux_h
    port map (
            O => \N__43800\,
            I => \N__43776\
        );

    \I__10801\ : Span4Mux_v
    port map (
            O => \N__43795\,
            I => \N__43776\
        );

    \I__10800\ : Odrv4
    port map (
            O => \N__43792\,
            I => \ALU.log_0_sqmuxa\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__43781\,
            I => \ALU.log_0_sqmuxa\
        );

    \I__10798\ : Odrv4
    port map (
            O => \N__43776\,
            I => \ALU.log_0_sqmuxa\
        );

    \I__10797\ : CascadeMux
    port map (
            O => \N__43769\,
            I => \N__43764\
        );

    \I__10796\ : InMux
    port map (
            O => \N__43768\,
            I => \N__43758\
        );

    \I__10795\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43755\
        );

    \I__10794\ : InMux
    port map (
            O => \N__43764\,
            I => \N__43751\
        );

    \I__10793\ : InMux
    port map (
            O => \N__43763\,
            I => \N__43748\
        );

    \I__10792\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43744\
        );

    \I__10791\ : InMux
    port map (
            O => \N__43761\,
            I => \N__43741\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__43758\,
            I => \N__43736\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__43755\,
            I => \N__43736\
        );

    \I__10788\ : InMux
    port map (
            O => \N__43754\,
            I => \N__43733\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__43751\,
            I => \N__43730\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__43748\,
            I => \N__43723\
        );

    \I__10785\ : CascadeMux
    port map (
            O => \N__43747\,
            I => \N__43720\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__43744\,
            I => \N__43716\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__43741\,
            I => \N__43708\
        );

    \I__10782\ : Span4Mux_v
    port map (
            O => \N__43736\,
            I => \N__43708\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__43733\,
            I => \N__43704\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__43730\,
            I => \N__43701\
        );

    \I__10779\ : InMux
    port map (
            O => \N__43729\,
            I => \N__43698\
        );

    \I__10778\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43694\
        );

    \I__10777\ : CascadeMux
    port map (
            O => \N__43727\,
            I => \N__43691\
        );

    \I__10776\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43685\
        );

    \I__10775\ : Span4Mux_v
    port map (
            O => \N__43723\,
            I => \N__43680\
        );

    \I__10774\ : InMux
    port map (
            O => \N__43720\,
            I => \N__43677\
        );

    \I__10773\ : CascadeMux
    port map (
            O => \N__43719\,
            I => \N__43670\
        );

    \I__10772\ : Span4Mux_v
    port map (
            O => \N__43716\,
            I => \N__43661\
        );

    \I__10771\ : InMux
    port map (
            O => \N__43715\,
            I => \N__43654\
        );

    \I__10770\ : InMux
    port map (
            O => \N__43714\,
            I => \N__43654\
        );

    \I__10769\ : InMux
    port map (
            O => \N__43713\,
            I => \N__43654\
        );

    \I__10768\ : Span4Mux_v
    port map (
            O => \N__43708\,
            I => \N__43650\
        );

    \I__10767\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43647\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__43704\,
            I => \N__43642\
        );

    \I__10765\ : Span4Mux_v
    port map (
            O => \N__43701\,
            I => \N__43642\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__43698\,
            I => \N__43639\
        );

    \I__10763\ : InMux
    port map (
            O => \N__43697\,
            I => \N__43635\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__43694\,
            I => \N__43632\
        );

    \I__10761\ : InMux
    port map (
            O => \N__43691\,
            I => \N__43629\
        );

    \I__10760\ : InMux
    port map (
            O => \N__43690\,
            I => \N__43626\
        );

    \I__10759\ : InMux
    port map (
            O => \N__43689\,
            I => \N__43623\
        );

    \I__10758\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43617\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__43685\,
            I => \N__43614\
        );

    \I__10756\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43609\
        );

    \I__10755\ : InMux
    port map (
            O => \N__43683\,
            I => \N__43609\
        );

    \I__10754\ : Span4Mux_v
    port map (
            O => \N__43680\,
            I => \N__43604\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__43677\,
            I => \N__43604\
        );

    \I__10752\ : InMux
    port map (
            O => \N__43676\,
            I => \N__43601\
        );

    \I__10751\ : InMux
    port map (
            O => \N__43675\,
            I => \N__43598\
        );

    \I__10750\ : InMux
    port map (
            O => \N__43674\,
            I => \N__43595\
        );

    \I__10749\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43588\
        );

    \I__10748\ : InMux
    port map (
            O => \N__43670\,
            I => \N__43588\
        );

    \I__10747\ : InMux
    port map (
            O => \N__43669\,
            I => \N__43588\
        );

    \I__10746\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43579\
        );

    \I__10745\ : InMux
    port map (
            O => \N__43667\,
            I => \N__43576\
        );

    \I__10744\ : InMux
    port map (
            O => \N__43666\,
            I => \N__43573\
        );

    \I__10743\ : InMux
    port map (
            O => \N__43665\,
            I => \N__43568\
        );

    \I__10742\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43568\
        );

    \I__10741\ : Span4Mux_v
    port map (
            O => \N__43661\,
            I => \N__43565\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__43654\,
            I => \N__43562\
        );

    \I__10739\ : InMux
    port map (
            O => \N__43653\,
            I => \N__43559\
        );

    \I__10738\ : Span4Mux_h
    port map (
            O => \N__43650\,
            I => \N__43552\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__43647\,
            I => \N__43552\
        );

    \I__10736\ : Span4Mux_v
    port map (
            O => \N__43642\,
            I => \N__43552\
        );

    \I__10735\ : Sp12to4
    port map (
            O => \N__43639\,
            I => \N__43549\
        );

    \I__10734\ : CascadeMux
    port map (
            O => \N__43638\,
            I => \N__43546\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__43635\,
            I => \N__43542\
        );

    \I__10732\ : Span4Mux_v
    port map (
            O => \N__43632\,
            I => \N__43533\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__43629\,
            I => \N__43533\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__43626\,
            I => \N__43533\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__43623\,
            I => \N__43533\
        );

    \I__10728\ : InMux
    port map (
            O => \N__43622\,
            I => \N__43528\
        );

    \I__10727\ : InMux
    port map (
            O => \N__43621\,
            I => \N__43528\
        );

    \I__10726\ : InMux
    port map (
            O => \N__43620\,
            I => \N__43525\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__43617\,
            I => \N__43522\
        );

    \I__10724\ : Span4Mux_h
    port map (
            O => \N__43614\,
            I => \N__43517\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__43609\,
            I => \N__43517\
        );

    \I__10722\ : Span4Mux_h
    port map (
            O => \N__43604\,
            I => \N__43512\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__43601\,
            I => \N__43512\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__43598\,
            I => \N__43507\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__43595\,
            I => \N__43502\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__43588\,
            I => \N__43502\
        );

    \I__10717\ : InMux
    port map (
            O => \N__43587\,
            I => \N__43495\
        );

    \I__10716\ : InMux
    port map (
            O => \N__43586\,
            I => \N__43495\
        );

    \I__10715\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43495\
        );

    \I__10714\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43492\
        );

    \I__10713\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43486\
        );

    \I__10712\ : InMux
    port map (
            O => \N__43582\,
            I => \N__43486\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__43579\,
            I => \N__43471\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__43576\,
            I => \N__43471\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__43573\,
            I => \N__43471\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__43568\,
            I => \N__43471\
        );

    \I__10707\ : Span4Mux_h
    port map (
            O => \N__43565\,
            I => \N__43471\
        );

    \I__10706\ : Span4Mux_h
    port map (
            O => \N__43562\,
            I => \N__43471\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__43559\,
            I => \N__43471\
        );

    \I__10704\ : Span4Mux_v
    port map (
            O => \N__43552\,
            I => \N__43468\
        );

    \I__10703\ : Span12Mux_v
    port map (
            O => \N__43549\,
            I => \N__43465\
        );

    \I__10702\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43460\
        );

    \I__10701\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43460\
        );

    \I__10700\ : Span4Mux_h
    port map (
            O => \N__43542\,
            I => \N__43455\
        );

    \I__10699\ : Span4Mux_h
    port map (
            O => \N__43533\,
            I => \N__43455\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__43528\,
            I => \N__43448\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__43525\,
            I => \N__43448\
        );

    \I__10696\ : Span4Mux_h
    port map (
            O => \N__43522\,
            I => \N__43448\
        );

    \I__10695\ : Span4Mux_v
    port map (
            O => \N__43517\,
            I => \N__43443\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__43512\,
            I => \N__43443\
        );

    \I__10693\ : InMux
    port map (
            O => \N__43511\,
            I => \N__43438\
        );

    \I__10692\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43438\
        );

    \I__10691\ : Span12Mux_h
    port map (
            O => \N__43507\,
            I => \N__43429\
        );

    \I__10690\ : Sp12to4
    port map (
            O => \N__43502\,
            I => \N__43429\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__43495\,
            I => \N__43429\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__43492\,
            I => \N__43429\
        );

    \I__10687\ : InMux
    port map (
            O => \N__43491\,
            I => \N__43426\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__43486\,
            I => \N__43419\
        );

    \I__10685\ : Span4Mux_v
    port map (
            O => \N__43471\,
            I => \N__43419\
        );

    \I__10684\ : Span4Mux_s1_v
    port map (
            O => \N__43468\,
            I => \N__43419\
        );

    \I__10683\ : Odrv12
    port map (
            O => \N__43465\,
            I => \aluParams_0\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__43460\,
            I => \aluParams_0\
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__43455\,
            I => \aluParams_0\
        );

    \I__10680\ : Odrv4
    port map (
            O => \N__43448\,
            I => \aluParams_0\
        );

    \I__10679\ : Odrv4
    port map (
            O => \N__43443\,
            I => \aluParams_0\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__43438\,
            I => \aluParams_0\
        );

    \I__10677\ : Odrv12
    port map (
            O => \N__43429\,
            I => \aluParams_0\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__43426\,
            I => \aluParams_0\
        );

    \I__10675\ : Odrv4
    port map (
            O => \N__43419\,
            I => \aluParams_0\
        );

    \I__10674\ : InMux
    port map (
            O => \N__43400\,
            I => \N__43397\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__43397\,
            I => \N__43393\
        );

    \I__10672\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43390\
        );

    \I__10671\ : Span4Mux_h
    port map (
            O => \N__43393\,
            I => \N__43387\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__43390\,
            I => \N__43384\
        );

    \I__10669\ : Span4Mux_h
    port map (
            O => \N__43387\,
            I => \N__43381\
        );

    \I__10668\ : Span4Mux_h
    port map (
            O => \N__43384\,
            I => \N__43378\
        );

    \I__10667\ : Odrv4
    port map (
            O => \N__43381\,
            I => \ALU.dZ0Z_5\
        );

    \I__10666\ : Odrv4
    port map (
            O => \N__43378\,
            I => \ALU.dZ0Z_5\
        );

    \I__10665\ : InMux
    port map (
            O => \N__43373\,
            I => \N__43369\
        );

    \I__10664\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43366\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__43369\,
            I => \N__43363\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__43366\,
            I => \N__43360\
        );

    \I__10661\ : Span4Mux_h
    port map (
            O => \N__43363\,
            I => \N__43357\
        );

    \I__10660\ : Span4Mux_h
    port map (
            O => \N__43360\,
            I => \N__43354\
        );

    \I__10659\ : Span4Mux_h
    port map (
            O => \N__43357\,
            I => \N__43351\
        );

    \I__10658\ : Odrv4
    port map (
            O => \N__43354\,
            I => \ALU.dZ0Z_6\
        );

    \I__10657\ : Odrv4
    port map (
            O => \N__43351\,
            I => \ALU.dZ0Z_6\
        );

    \I__10656\ : CEMux
    port map (
            O => \N__43346\,
            I => \N__43341\
        );

    \I__10655\ : CEMux
    port map (
            O => \N__43345\,
            I => \N__43337\
        );

    \I__10654\ : CEMux
    port map (
            O => \N__43344\,
            I => \N__43334\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__43341\,
            I => \N__43331\
        );

    \I__10652\ : CEMux
    port map (
            O => \N__43340\,
            I => \N__43328\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__43337\,
            I => \N__43325\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__43334\,
            I => \N__43321\
        );

    \I__10649\ : Span4Mux_h
    port map (
            O => \N__43331\,
            I => \N__43318\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__43328\,
            I => \N__43315\
        );

    \I__10647\ : Span4Mux_v
    port map (
            O => \N__43325\,
            I => \N__43312\
        );

    \I__10646\ : CEMux
    port map (
            O => \N__43324\,
            I => \N__43309\
        );

    \I__10645\ : Sp12to4
    port map (
            O => \N__43321\,
            I => \N__43306\
        );

    \I__10644\ : Span4Mux_v
    port map (
            O => \N__43318\,
            I => \N__43301\
        );

    \I__10643\ : Span4Mux_h
    port map (
            O => \N__43315\,
            I => \N__43301\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__43312\,
            I => \N__43298\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__43309\,
            I => \N__43295\
        );

    \I__10640\ : Span12Mux_h
    port map (
            O => \N__43306\,
            I => \N__43292\
        );

    \I__10639\ : Sp12to4
    port map (
            O => \N__43301\,
            I => \N__43287\
        );

    \I__10638\ : Sp12to4
    port map (
            O => \N__43298\,
            I => \N__43287\
        );

    \I__10637\ : Span4Mux_s1_v
    port map (
            O => \N__43295\,
            I => \N__43284\
        );

    \I__10636\ : Span12Mux_v
    port map (
            O => \N__43292\,
            I => \N__43281\
        );

    \I__10635\ : Span12Mux_v
    port map (
            O => \N__43287\,
            I => \N__43278\
        );

    \I__10634\ : Span4Mux_h
    port map (
            O => \N__43284\,
            I => \N__43275\
        );

    \I__10633\ : Odrv12
    port map (
            O => \N__43281\,
            I => \ALU.d_cnvZ0Z_0\
        );

    \I__10632\ : Odrv12
    port map (
            O => \N__43278\,
            I => \ALU.d_cnvZ0Z_0\
        );

    \I__10631\ : Odrv4
    port map (
            O => \N__43275\,
            I => \ALU.d_cnvZ0Z_0\
        );

    \I__10630\ : CascadeMux
    port map (
            O => \N__43268\,
            I => \N__43265\
        );

    \I__10629\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43262\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__43262\,
            I => \N__43258\
        );

    \I__10627\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43255\
        );

    \I__10626\ : Span4Mux_v
    port map (
            O => \N__43258\,
            I => \N__43252\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__43255\,
            I => \ALU.fZ0Z_3\
        );

    \I__10624\ : Odrv4
    port map (
            O => \N__43252\,
            I => \ALU.fZ0Z_3\
        );

    \I__10623\ : InMux
    port map (
            O => \N__43247\,
            I => \N__43244\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__43244\,
            I => \N__43241\
        );

    \I__10621\ : Span4Mux_v
    port map (
            O => \N__43241\,
            I => \N__43238\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__43238\,
            I => \N__43235\
        );

    \I__10619\ : Odrv4
    port map (
            O => \N__43235\,
            I => \ALU.f_RNIHUEJZ0Z_3\
        );

    \I__10618\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43228\
        );

    \I__10617\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43225\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__43228\,
            I => \N__43222\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__43225\,
            I => \N__43219\
        );

    \I__10614\ : Span12Mux_v
    port map (
            O => \N__43222\,
            I => \N__43216\
        );

    \I__10613\ : Odrv12
    port map (
            O => \N__43219\,
            I => \ALU.rshift_1_12\
        );

    \I__10612\ : Odrv12
    port map (
            O => \N__43216\,
            I => \ALU.rshift_1_12\
        );

    \I__10611\ : InMux
    port map (
            O => \N__43211\,
            I => \N__43208\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__43208\,
            I => \N__43205\
        );

    \I__10609\ : Span4Mux_v
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__10608\ : Sp12to4
    port map (
            O => \N__43202\,
            I => \N__43199\
        );

    \I__10607\ : Span12Mux_h
    port map (
            O => \N__43199\,
            I => \N__43196\
        );

    \I__10606\ : Odrv12
    port map (
            O => \N__43196\,
            I => \ALU.N_532\
        );

    \I__10605\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43190\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__43190\,
            I => \N__43186\
        );

    \I__10603\ : CascadeMux
    port map (
            O => \N__43189\,
            I => \N__43181\
        );

    \I__10602\ : Span4Mux_v
    port map (
            O => \N__43186\,
            I => \N__43176\
        );

    \I__10601\ : InMux
    port map (
            O => \N__43185\,
            I => \N__43173\
        );

    \I__10600\ : CascadeMux
    port map (
            O => \N__43184\,
            I => \N__43169\
        );

    \I__10599\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43166\
        );

    \I__10598\ : CascadeMux
    port map (
            O => \N__43180\,
            I => \N__43162\
        );

    \I__10597\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43159\
        );

    \I__10596\ : Span4Mux_v
    port map (
            O => \N__43176\,
            I => \N__43156\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__43173\,
            I => \N__43153\
        );

    \I__10594\ : InMux
    port map (
            O => \N__43172\,
            I => \N__43144\
        );

    \I__10593\ : InMux
    port map (
            O => \N__43169\,
            I => \N__43144\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__43166\,
            I => \N__43141\
        );

    \I__10591\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43136\
        );

    \I__10590\ : InMux
    port map (
            O => \N__43162\,
            I => \N__43133\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__43159\,
            I => \N__43130\
        );

    \I__10588\ : Span4Mux_v
    port map (
            O => \N__43156\,
            I => \N__43125\
        );

    \I__10587\ : Span4Mux_v
    port map (
            O => \N__43153\,
            I => \N__43125\
        );

    \I__10586\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43120\
        );

    \I__10585\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43120\
        );

    \I__10584\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43117\
        );

    \I__10583\ : InMux
    port map (
            O => \N__43149\,
            I => \N__43114\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__43144\,
            I => \N__43111\
        );

    \I__10581\ : Span4Mux_v
    port map (
            O => \N__43141\,
            I => \N__43106\
        );

    \I__10580\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43101\
        );

    \I__10579\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43101\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__43136\,
            I => \N__43098\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__43133\,
            I => \N__43094\
        );

    \I__10576\ : Span4Mux_v
    port map (
            O => \N__43130\,
            I => \N__43091\
        );

    \I__10575\ : Span4Mux_v
    port map (
            O => \N__43125\,
            I => \N__43087\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__43120\,
            I => \N__43082\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__43117\,
            I => \N__43082\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__43114\,
            I => \N__43077\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__43111\,
            I => \N__43077\
        );

    \I__10570\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43072\
        );

    \I__10569\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43072\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__43106\,
            I => \N__43067\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__43101\,
            I => \N__43067\
        );

    \I__10566\ : Span4Mux_v
    port map (
            O => \N__43098\,
            I => \N__43064\
        );

    \I__10565\ : InMux
    port map (
            O => \N__43097\,
            I => \N__43061\
        );

    \I__10564\ : Span4Mux_s3_h
    port map (
            O => \N__43094\,
            I => \N__43056\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__43091\,
            I => \N__43056\
        );

    \I__10562\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43053\
        );

    \I__10561\ : Span4Mux_h
    port map (
            O => \N__43087\,
            I => \N__43048\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__43082\,
            I => \N__43048\
        );

    \I__10559\ : Span4Mux_h
    port map (
            O => \N__43077\,
            I => \N__43043\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__43072\,
            I => \N__43043\
        );

    \I__10557\ : Span4Mux_v
    port map (
            O => \N__43067\,
            I => \N__43038\
        );

    \I__10556\ : Span4Mux_h
    port map (
            O => \N__43064\,
            I => \N__43038\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__43061\,
            I => \aluOperation_4\
        );

    \I__10554\ : Odrv4
    port map (
            O => \N__43056\,
            I => \aluOperation_4\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__43053\,
            I => \aluOperation_4\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__43048\,
            I => \aluOperation_4\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__43043\,
            I => \aluOperation_4\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__43038\,
            I => \aluOperation_4\
        );

    \I__10549\ : CascadeMux
    port map (
            O => \N__43025\,
            I => \ALU.rshift_4_cascade_\
        );

    \I__10548\ : InMux
    port map (
            O => \N__43022\,
            I => \N__43019\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__43019\,
            I => \N__43016\
        );

    \I__10546\ : Span4Mux_v
    port map (
            O => \N__43016\,
            I => \N__43013\
        );

    \I__10545\ : Span4Mux_v
    port map (
            O => \N__43013\,
            I => \N__43010\
        );

    \I__10544\ : Span4Mux_h
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__43007\,
            I => \N__43004\
        );

    \I__10542\ : Odrv4
    port map (
            O => \N__43004\,
            I => \ALU.N_289_0\
        );

    \I__10541\ : CascadeMux
    port map (
            O => \N__43001\,
            I => \ALU.a_15_m3_4_cascade_\
        );

    \I__10540\ : InMux
    port map (
            O => \N__42998\,
            I => \N__42987\
        );

    \I__10539\ : CascadeMux
    port map (
            O => \N__42997\,
            I => \N__42984\
        );

    \I__10538\ : InMux
    port map (
            O => \N__42996\,
            I => \N__42981\
        );

    \I__10537\ : InMux
    port map (
            O => \N__42995\,
            I => \N__42977\
        );

    \I__10536\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42974\
        );

    \I__10535\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42966\
        );

    \I__10534\ : InMux
    port map (
            O => \N__42992\,
            I => \N__42963\
        );

    \I__10533\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42960\
        );

    \I__10532\ : CascadeMux
    port map (
            O => \N__42990\,
            I => \N__42954\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__42987\,
            I => \N__42951\
        );

    \I__10530\ : InMux
    port map (
            O => \N__42984\,
            I => \N__42948\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__42981\,
            I => \N__42942\
        );

    \I__10528\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42939\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__42977\,
            I => \N__42934\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__42974\,
            I => \N__42934\
        );

    \I__10525\ : InMux
    port map (
            O => \N__42973\,
            I => \N__42928\
        );

    \I__10524\ : InMux
    port map (
            O => \N__42972\,
            I => \N__42928\
        );

    \I__10523\ : CascadeMux
    port map (
            O => \N__42971\,
            I => \N__42923\
        );

    \I__10522\ : CascadeMux
    port map (
            O => \N__42970\,
            I => \N__42920\
        );

    \I__10521\ : CascadeMux
    port map (
            O => \N__42969\,
            I => \N__42917\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__42966\,
            I => \N__42913\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__42963\,
            I => \N__42910\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__42960\,
            I => \N__42907\
        );

    \I__10517\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42900\
        );

    \I__10516\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42897\
        );

    \I__10515\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42892\
        );

    \I__10514\ : InMux
    port map (
            O => \N__42954\,
            I => \N__42892\
        );

    \I__10513\ : Span4Mux_s3_v
    port map (
            O => \N__42951\,
            I => \N__42886\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__42948\,
            I => \N__42886\
        );

    \I__10511\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42879\
        );

    \I__10510\ : InMux
    port map (
            O => \N__42946\,
            I => \N__42879\
        );

    \I__10509\ : InMux
    port map (
            O => \N__42945\,
            I => \N__42879\
        );

    \I__10508\ : Span4Mux_s3_v
    port map (
            O => \N__42942\,
            I => \N__42874\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__42939\,
            I => \N__42874\
        );

    \I__10506\ : Span4Mux_h
    port map (
            O => \N__42934\,
            I => \N__42871\
        );

    \I__10505\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42868\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__42928\,
            I => \N__42865\
        );

    \I__10503\ : InMux
    port map (
            O => \N__42927\,
            I => \N__42862\
        );

    \I__10502\ : InMux
    port map (
            O => \N__42926\,
            I => \N__42859\
        );

    \I__10501\ : InMux
    port map (
            O => \N__42923\,
            I => \N__42856\
        );

    \I__10500\ : InMux
    port map (
            O => \N__42920\,
            I => \N__42849\
        );

    \I__10499\ : InMux
    port map (
            O => \N__42917\,
            I => \N__42849\
        );

    \I__10498\ : InMux
    port map (
            O => \N__42916\,
            I => \N__42849\
        );

    \I__10497\ : Span4Mux_v
    port map (
            O => \N__42913\,
            I => \N__42844\
        );

    \I__10496\ : Span4Mux_v
    port map (
            O => \N__42910\,
            I => \N__42844\
        );

    \I__10495\ : Span4Mux_v
    port map (
            O => \N__42907\,
            I => \N__42841\
        );

    \I__10494\ : InMux
    port map (
            O => \N__42906\,
            I => \N__42838\
        );

    \I__10493\ : InMux
    port map (
            O => \N__42905\,
            I => \N__42835\
        );

    \I__10492\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42830\
        );

    \I__10491\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42830\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__42900\,
            I => \N__42827\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__42897\,
            I => \N__42824\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__42892\,
            I => \N__42818\
        );

    \I__10487\ : InMux
    port map (
            O => \N__42891\,
            I => \N__42815\
        );

    \I__10486\ : Span4Mux_h
    port map (
            O => \N__42886\,
            I => \N__42810\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__42879\,
            I => \N__42810\
        );

    \I__10484\ : Span4Mux_v
    port map (
            O => \N__42874\,
            I => \N__42807\
        );

    \I__10483\ : Span4Mux_v
    port map (
            O => \N__42871\,
            I => \N__42800\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__42868\,
            I => \N__42800\
        );

    \I__10481\ : Span4Mux_s2_h
    port map (
            O => \N__42865\,
            I => \N__42800\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__42862\,
            I => \N__42797\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__42859\,
            I => \N__42790\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__42856\,
            I => \N__42790\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__42849\,
            I => \N__42790\
        );

    \I__10476\ : Span4Mux_h
    port map (
            O => \N__42844\,
            I => \N__42782\
        );

    \I__10475\ : Span4Mux_v
    port map (
            O => \N__42841\,
            I => \N__42782\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__42838\,
            I => \N__42777\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__42835\,
            I => \N__42777\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__42830\,
            I => \N__42774\
        );

    \I__10471\ : Span4Mux_v
    port map (
            O => \N__42827\,
            I => \N__42769\
        );

    \I__10470\ : Span4Mux_s1_h
    port map (
            O => \N__42824\,
            I => \N__42769\
        );

    \I__10469\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42764\
        );

    \I__10468\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42764\
        );

    \I__10467\ : InMux
    port map (
            O => \N__42821\,
            I => \N__42761\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__42818\,
            I => \N__42758\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__42815\,
            I => \N__42753\
        );

    \I__10464\ : Span4Mux_v
    port map (
            O => \N__42810\,
            I => \N__42753\
        );

    \I__10463\ : Span4Mux_v
    port map (
            O => \N__42807\,
            I => \N__42748\
        );

    \I__10462\ : Span4Mux_v
    port map (
            O => \N__42800\,
            I => \N__42748\
        );

    \I__10461\ : Span4Mux_h
    port map (
            O => \N__42797\,
            I => \N__42743\
        );

    \I__10460\ : Span4Mux_v
    port map (
            O => \N__42790\,
            I => \N__42743\
        );

    \I__10459\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42738\
        );

    \I__10458\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42738\
        );

    \I__10457\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42735\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__42782\,
            I => \N__42724\
        );

    \I__10455\ : Span4Mux_h
    port map (
            O => \N__42777\,
            I => \N__42724\
        );

    \I__10454\ : Span4Mux_v
    port map (
            O => \N__42774\,
            I => \N__42724\
        );

    \I__10453\ : Span4Mux_h
    port map (
            O => \N__42769\,
            I => \N__42724\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__42764\,
            I => \N__42724\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__42761\,
            I => \ALU.aluOut_4\
        );

    \I__10450\ : Odrv4
    port map (
            O => \N__42758\,
            I => \ALU.aluOut_4\
        );

    \I__10449\ : Odrv4
    port map (
            O => \N__42753\,
            I => \ALU.aluOut_4\
        );

    \I__10448\ : Odrv4
    port map (
            O => \N__42748\,
            I => \ALU.aluOut_4\
        );

    \I__10447\ : Odrv4
    port map (
            O => \N__42743\,
            I => \ALU.aluOut_4\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__42738\,
            I => \ALU.aluOut_4\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__42735\,
            I => \ALU.aluOut_4\
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__42724\,
            I => \ALU.aluOut_4\
        );

    \I__10443\ : CascadeMux
    port map (
            O => \N__42707\,
            I => \N__42704\
        );

    \I__10442\ : InMux
    port map (
            O => \N__42704\,
            I => \N__42701\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__42701\,
            I => \ALU.a_15_m2_ns_1Z0Z_4\
        );

    \I__10440\ : CascadeMux
    port map (
            O => \N__42698\,
            I => \N__42693\
        );

    \I__10439\ : InMux
    port map (
            O => \N__42697\,
            I => \N__42684\
        );

    \I__10438\ : InMux
    port map (
            O => \N__42696\,
            I => \N__42680\
        );

    \I__10437\ : InMux
    port map (
            O => \N__42693\,
            I => \N__42677\
        );

    \I__10436\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42668\
        );

    \I__10435\ : InMux
    port map (
            O => \N__42691\,
            I => \N__42668\
        );

    \I__10434\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42668\
        );

    \I__10433\ : InMux
    port map (
            O => \N__42689\,
            I => \N__42663\
        );

    \I__10432\ : InMux
    port map (
            O => \N__42688\,
            I => \N__42657\
        );

    \I__10431\ : InMux
    port map (
            O => \N__42687\,
            I => \N__42657\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__42684\,
            I => \N__42654\
        );

    \I__10429\ : InMux
    port map (
            O => \N__42683\,
            I => \N__42651\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__42680\,
            I => \N__42648\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__42677\,
            I => \N__42645\
        );

    \I__10426\ : InMux
    port map (
            O => \N__42676\,
            I => \N__42639\
        );

    \I__10425\ : InMux
    port map (
            O => \N__42675\,
            I => \N__42639\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__42668\,
            I => \N__42636\
        );

    \I__10423\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42631\
        );

    \I__10422\ : InMux
    port map (
            O => \N__42666\,
            I => \N__42631\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__42663\,
            I => \N__42628\
        );

    \I__10420\ : InMux
    port map (
            O => \N__42662\,
            I => \N__42625\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__42657\,
            I => \N__42622\
        );

    \I__10418\ : Span4Mux_v
    port map (
            O => \N__42654\,
            I => \N__42619\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__42651\,
            I => \N__42616\
        );

    \I__10416\ : Span4Mux_h
    port map (
            O => \N__42648\,
            I => \N__42611\
        );

    \I__10415\ : Span4Mux_h
    port map (
            O => \N__42645\,
            I => \N__42611\
        );

    \I__10414\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42608\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__42639\,
            I => \N__42603\
        );

    \I__10412\ : Span4Mux_s2_h
    port map (
            O => \N__42636\,
            I => \N__42603\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__42631\,
            I => \N__42598\
        );

    \I__10410\ : Span4Mux_s2_h
    port map (
            O => \N__42628\,
            I => \N__42598\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__42625\,
            I => \N__42595\
        );

    \I__10408\ : Span4Mux_s3_h
    port map (
            O => \N__42622\,
            I => \N__42592\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__42619\,
            I => \N__42587\
        );

    \I__10406\ : Span4Mux_v
    port map (
            O => \N__42616\,
            I => \N__42587\
        );

    \I__10405\ : Span4Mux_v
    port map (
            O => \N__42611\,
            I => \N__42584\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__42608\,
            I => \N__42577\
        );

    \I__10403\ : Span4Mux_h
    port map (
            O => \N__42603\,
            I => \N__42577\
        );

    \I__10402\ : Span4Mux_h
    port map (
            O => \N__42598\,
            I => \N__42577\
        );

    \I__10401\ : Span4Mux_s3_h
    port map (
            O => \N__42595\,
            I => \N__42572\
        );

    \I__10400\ : Span4Mux_v
    port map (
            O => \N__42592\,
            I => \N__42572\
        );

    \I__10399\ : Odrv4
    port map (
            O => \N__42587\,
            I => \ALU.N_231_0\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__42584\,
            I => \ALU.N_231_0\
        );

    \I__10397\ : Odrv4
    port map (
            O => \N__42577\,
            I => \ALU.N_231_0\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__42572\,
            I => \ALU.N_231_0\
        );

    \I__10395\ : InMux
    port map (
            O => \N__42563\,
            I => \N__42560\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__42560\,
            I => \N__42557\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__42557\,
            I => \ALU.un9_addsub_cry_4_c_RNIL4NZ0Z97\
        );

    \I__10392\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42551\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__42551\,
            I => \N__42548\
        );

    \I__10390\ : Span4Mux_v
    port map (
            O => \N__42548\,
            I => \N__42545\
        );

    \I__10389\ : Span4Mux_h
    port map (
            O => \N__42545\,
            I => \N__42542\
        );

    \I__10388\ : Odrv4
    port map (
            O => \N__42542\,
            I => \ALU.un2_addsub_cry_4_c_RNI284VEZ0\
        );

    \I__10387\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42536\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__42536\,
            I => \N__42533\
        );

    \I__10385\ : Odrv4
    port map (
            O => \N__42533\,
            I => \ALU.un9_addsub_cry_5_c_RNI6SCFZ0Z7\
        );

    \I__10384\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42527\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__42527\,
            I => \N__42523\
        );

    \I__10382\ : CascadeMux
    port map (
            O => \N__42526\,
            I => \N__42519\
        );

    \I__10381\ : Span4Mux_v
    port map (
            O => \N__42523\,
            I => \N__42514\
        );

    \I__10380\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42511\
        );

    \I__10379\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42508\
        );

    \I__10378\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42499\
        );

    \I__10377\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42496\
        );

    \I__10376\ : Span4Mux_h
    port map (
            O => \N__42514\,
            I => \N__42490\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__42511\,
            I => \N__42490\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__42508\,
            I => \N__42487\
        );

    \I__10373\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42482\
        );

    \I__10372\ : InMux
    port map (
            O => \N__42506\,
            I => \N__42482\
        );

    \I__10371\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42473\
        );

    \I__10370\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42473\
        );

    \I__10369\ : InMux
    port map (
            O => \N__42503\,
            I => \N__42473\
        );

    \I__10368\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42473\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__42499\,
            I => \N__42470\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__42496\,
            I => \N__42467\
        );

    \I__10365\ : InMux
    port map (
            O => \N__42495\,
            I => \N__42464\
        );

    \I__10364\ : Span4Mux_v
    port map (
            O => \N__42490\,
            I => \N__42460\
        );

    \I__10363\ : Span4Mux_v
    port map (
            O => \N__42487\,
            I => \N__42445\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__42482\,
            I => \N__42445\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__42473\,
            I => \N__42445\
        );

    \I__10360\ : Span4Mux_h
    port map (
            O => \N__42470\,
            I => \N__42445\
        );

    \I__10359\ : Span4Mux_v
    port map (
            O => \N__42467\,
            I => \N__42445\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__42464\,
            I => \N__42445\
        );

    \I__10357\ : InMux
    port map (
            O => \N__42463\,
            I => \N__42442\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__42460\,
            I => \N__42439\
        );

    \I__10355\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42436\
        );

    \I__10354\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42433\
        );

    \I__10353\ : Span4Mux_v
    port map (
            O => \N__42445\,
            I => \N__42430\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__42442\,
            I => \ALU.addsub_0_sqmuxa\
        );

    \I__10351\ : Odrv4
    port map (
            O => \N__42439\,
            I => \ALU.addsub_0_sqmuxa\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__42436\,
            I => \ALU.addsub_0_sqmuxa\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__42433\,
            I => \ALU.addsub_0_sqmuxa\
        );

    \I__10348\ : Odrv4
    port map (
            O => \N__42430\,
            I => \ALU.addsub_0_sqmuxa\
        );

    \I__10347\ : InMux
    port map (
            O => \N__42419\,
            I => \N__42416\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__42416\,
            I => \N__42413\
        );

    \I__10345\ : Span4Mux_h
    port map (
            O => \N__42413\,
            I => \N__42410\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__42410\,
            I => \N__42407\
        );

    \I__10343\ : Odrv4
    port map (
            O => \N__42407\,
            I => \ALU.un2_addsub_cry_5_c_RNIL7IGFZ0\
        );

    \I__10342\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42401\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__42401\,
            I => \N__42398\
        );

    \I__10340\ : Span4Mux_v
    port map (
            O => \N__42398\,
            I => \N__42395\
        );

    \I__10339\ : Span4Mux_h
    port map (
            O => \N__42395\,
            I => \N__42392\
        );

    \I__10338\ : Odrv4
    port map (
            O => \N__42392\,
            I => \ALU.N_422\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__42389\,
            I => \ALU.d_RNIP43E91Z0Z_7_cascade_\
        );

    \I__10336\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42383\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__42383\,
            I => \N__42380\
        );

    \I__10334\ : Span4Mux_v
    port map (
            O => \N__42380\,
            I => \N__42377\
        );

    \I__10333\ : Span4Mux_h
    port map (
            O => \N__42377\,
            I => \N__42374\
        );

    \I__10332\ : Odrv4
    port map (
            O => \N__42374\,
            I => \ALU.d_RNIT87FA1Z0Z_7\
        );

    \I__10331\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42368\
        );

    \I__10330\ : LocalMux
    port map (
            O => \N__42368\,
            I => \N__42365\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__42365\,
            I => \N__42362\
        );

    \I__10328\ : Span4Mux_h
    port map (
            O => \N__42362\,
            I => \N__42359\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__42359\,
            I => \ALU.madd_cry_5_THRU_CO\
        );

    \I__10326\ : CascadeMux
    port map (
            O => \N__42356\,
            I => \ALU.a_15_m5_7_cascade_\
        );

    \I__10325\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42350\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__42350\,
            I => \N__42346\
        );

    \I__10323\ : InMux
    port map (
            O => \N__42349\,
            I => \N__42343\
        );

    \I__10322\ : Span4Mux_v
    port map (
            O => \N__42346\,
            I => \N__42340\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__42343\,
            I => \N__42337\
        );

    \I__10320\ : Span4Mux_h
    port map (
            O => \N__42340\,
            I => \N__42332\
        );

    \I__10319\ : Span4Mux_v
    port map (
            O => \N__42337\,
            I => \N__42332\
        );

    \I__10318\ : Span4Mux_h
    port map (
            O => \N__42332\,
            I => \N__42329\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__42329\,
            I => \ALU.madd_axb_6\
        );

    \I__10316\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42323\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__42323\,
            I => \N__42318\
        );

    \I__10314\ : InMux
    port map (
            O => \N__42322\,
            I => \N__42315\
        );

    \I__10313\ : InMux
    port map (
            O => \N__42321\,
            I => \N__42312\
        );

    \I__10312\ : Span4Mux_h
    port map (
            O => \N__42318\,
            I => \N__42308\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__42315\,
            I => \N__42305\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__42312\,
            I => \N__42302\
        );

    \I__10309\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42299\
        );

    \I__10308\ : Span4Mux_h
    port map (
            O => \N__42308\,
            I => \N__42289\
        );

    \I__10307\ : Span4Mux_v
    port map (
            O => \N__42305\,
            I => \N__42289\
        );

    \I__10306\ : Span4Mux_v
    port map (
            O => \N__42302\,
            I => \N__42289\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__42299\,
            I => \N__42286\
        );

    \I__10304\ : InMux
    port map (
            O => \N__42298\,
            I => \N__42283\
        );

    \I__10303\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42280\
        );

    \I__10302\ : InMux
    port map (
            O => \N__42296\,
            I => \N__42277\
        );

    \I__10301\ : Odrv4
    port map (
            O => \N__42289\,
            I => \ALU.d_RNIO75MAZ0Z_0\
        );

    \I__10300\ : Odrv12
    port map (
            O => \N__42286\,
            I => \ALU.d_RNIO75MAZ0Z_0\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__42283\,
            I => \ALU.d_RNIO75MAZ0Z_0\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__42280\,
            I => \ALU.d_RNIO75MAZ0Z_0\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__42277\,
            I => \ALU.d_RNIO75MAZ0Z_0\
        );

    \I__10296\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42261\
        );

    \I__10295\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42258\
        );

    \I__10294\ : InMux
    port map (
            O => \N__42264\,
            I => \N__42255\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__42261\,
            I => \N__42249\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__42258\,
            I => \N__42246\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__42255\,
            I => \N__42243\
        );

    \I__10290\ : InMux
    port map (
            O => \N__42254\,
            I => \N__42240\
        );

    \I__10289\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42237\
        );

    \I__10288\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42234\
        );

    \I__10287\ : Span4Mux_v
    port map (
            O => \N__42249\,
            I => \N__42228\
        );

    \I__10286\ : Span4Mux_v
    port map (
            O => \N__42246\,
            I => \N__42228\
        );

    \I__10285\ : Span4Mux_v
    port map (
            O => \N__42243\,
            I => \N__42225\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__42240\,
            I => \N__42222\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__42237\,
            I => \N__42219\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__42234\,
            I => \N__42216\
        );

    \I__10281\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42213\
        );

    \I__10280\ : Span4Mux_h
    port map (
            O => \N__42228\,
            I => \N__42210\
        );

    \I__10279\ : Span4Mux_h
    port map (
            O => \N__42225\,
            I => \N__42199\
        );

    \I__10278\ : Span4Mux_v
    port map (
            O => \N__42222\,
            I => \N__42199\
        );

    \I__10277\ : Span4Mux_h
    port map (
            O => \N__42219\,
            I => \N__42199\
        );

    \I__10276\ : Span4Mux_v
    port map (
            O => \N__42216\,
            I => \N__42199\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__42213\,
            I => \N__42199\
        );

    \I__10274\ : Odrv4
    port map (
            O => \N__42210\,
            I => \ALU.d_RNI9BO713Z0Z_0\
        );

    \I__10273\ : Odrv4
    port map (
            O => \N__42199\,
            I => \ALU.d_RNI9BO713Z0Z_0\
        );

    \I__10272\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42190\
        );

    \I__10271\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42187\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__42190\,
            I => \N__42184\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__42187\,
            I => \N__42181\
        );

    \I__10268\ : Span4Mux_h
    port map (
            O => \N__42184\,
            I => \N__42178\
        );

    \I__10267\ : Span4Mux_h
    port map (
            O => \N__42181\,
            I => \N__42175\
        );

    \I__10266\ : Span4Mux_h
    port map (
            O => \N__42178\,
            I => \N__42172\
        );

    \I__10265\ : Span4Mux_h
    port map (
            O => \N__42175\,
            I => \N__42169\
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__42172\,
            I => \ALU.dZ0Z_0\
        );

    \I__10263\ : Odrv4
    port map (
            O => \N__42169\,
            I => \ALU.dZ0Z_0\
        );

    \I__10262\ : InMux
    port map (
            O => \N__42164\,
            I => \N__42158\
        );

    \I__10261\ : InMux
    port map (
            O => \N__42163\,
            I => \N__42155\
        );

    \I__10260\ : InMux
    port map (
            O => \N__42162\,
            I => \N__42152\
        );

    \I__10259\ : InMux
    port map (
            O => \N__42161\,
            I => \N__42147\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__42158\,
            I => \N__42139\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__42155\,
            I => \N__42139\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__42152\,
            I => \N__42139\
        );

    \I__10255\ : InMux
    port map (
            O => \N__42151\,
            I => \N__42136\
        );

    \I__10254\ : InMux
    port map (
            O => \N__42150\,
            I => \N__42133\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__42147\,
            I => \N__42130\
        );

    \I__10252\ : InMux
    port map (
            O => \N__42146\,
            I => \N__42127\
        );

    \I__10251\ : Span4Mux_v
    port map (
            O => \N__42139\,
            I => \N__42119\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__42136\,
            I => \N__42119\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__42133\,
            I => \N__42119\
        );

    \I__10248\ : Span4Mux_h
    port map (
            O => \N__42130\,
            I => \N__42114\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__42127\,
            I => \N__42114\
        );

    \I__10246\ : InMux
    port map (
            O => \N__42126\,
            I => \N__42111\
        );

    \I__10245\ : Span4Mux_h
    port map (
            O => \N__42119\,
            I => \N__42108\
        );

    \I__10244\ : Sp12to4
    port map (
            O => \N__42114\,
            I => \N__42103\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__42111\,
            I => \N__42103\
        );

    \I__10242\ : Odrv4
    port map (
            O => \N__42108\,
            I => \ALU.un9_addsub_cry_1_c_RNIM56ULZ0\
        );

    \I__10241\ : Odrv12
    port map (
            O => \N__42103\,
            I => \ALU.un9_addsub_cry_1_c_RNIM56ULZ0\
        );

    \I__10240\ : InMux
    port map (
            O => \N__42098\,
            I => \N__42093\
        );

    \I__10239\ : InMux
    port map (
            O => \N__42097\,
            I => \N__42089\
        );

    \I__10238\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42086\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__42093\,
            I => \N__42083\
        );

    \I__10236\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42080\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__42089\,
            I => \N__42073\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__42086\,
            I => \N__42073\
        );

    \I__10233\ : Span4Mux_v
    port map (
            O => \N__42083\,
            I => \N__42069\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__42080\,
            I => \N__42066\
        );

    \I__10231\ : InMux
    port map (
            O => \N__42079\,
            I => \N__42063\
        );

    \I__10230\ : InMux
    port map (
            O => \N__42078\,
            I => \N__42060\
        );

    \I__10229\ : Span4Mux_v
    port map (
            O => \N__42073\,
            I => \N__42057\
        );

    \I__10228\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42054\
        );

    \I__10227\ : Span4Mux_h
    port map (
            O => \N__42069\,
            I => \N__42045\
        );

    \I__10226\ : Span4Mux_v
    port map (
            O => \N__42066\,
            I => \N__42045\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__42063\,
            I => \N__42045\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__42060\,
            I => \N__42045\
        );

    \I__10223\ : Odrv4
    port map (
            O => \N__42057\,
            I => \ALU.d_RNIIFMN04Z0Z_2\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__42054\,
            I => \ALU.d_RNIIFMN04Z0Z_2\
        );

    \I__10221\ : Odrv4
    port map (
            O => \N__42045\,
            I => \ALU.d_RNIIFMN04Z0Z_2\
        );

    \I__10220\ : InMux
    port map (
            O => \N__42038\,
            I => \N__42035\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__42035\,
            I => \N__42031\
        );

    \I__10218\ : InMux
    port map (
            O => \N__42034\,
            I => \N__42028\
        );

    \I__10217\ : Span4Mux_v
    port map (
            O => \N__42031\,
            I => \N__42023\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__42028\,
            I => \N__42023\
        );

    \I__10215\ : Span4Mux_v
    port map (
            O => \N__42023\,
            I => \N__42020\
        );

    \I__10214\ : Odrv4
    port map (
            O => \N__42020\,
            I => \ALU.dZ0Z_2\
        );

    \I__10213\ : InMux
    port map (
            O => \N__42017\,
            I => \N__42006\
        );

    \I__10212\ : InMux
    port map (
            O => \N__42016\,
            I => \N__42006\
        );

    \I__10211\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42002\
        );

    \I__10210\ : InMux
    port map (
            O => \N__42014\,
            I => \N__41999\
        );

    \I__10209\ : InMux
    port map (
            O => \N__42013\,
            I => \N__41996\
        );

    \I__10208\ : InMux
    port map (
            O => \N__42012\,
            I => \N__41989\
        );

    \I__10207\ : InMux
    port map (
            O => \N__42011\,
            I => \N__41986\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__42006\,
            I => \N__41983\
        );

    \I__10205\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41980\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__42002\,
            I => \N__41966\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__41999\,
            I => \N__41966\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__41996\,
            I => \N__41966\
        );

    \I__10201\ : InMux
    port map (
            O => \N__41995\,
            I => \N__41963\
        );

    \I__10200\ : InMux
    port map (
            O => \N__41994\,
            I => \N__41960\
        );

    \I__10199\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41956\
        );

    \I__10198\ : InMux
    port map (
            O => \N__41992\,
            I => \N__41952\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__41989\,
            I => \N__41947\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__41986\,
            I => \N__41947\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__41983\,
            I => \N__41944\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__41980\,
            I => \N__41938\
        );

    \I__10193\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41931\
        );

    \I__10192\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41931\
        );

    \I__10191\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41931\
        );

    \I__10190\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41928\
        );

    \I__10189\ : CascadeMux
    port map (
            O => \N__41975\,
            I => \N__41923\
        );

    \I__10188\ : InMux
    port map (
            O => \N__41974\,
            I => \N__41920\
        );

    \I__10187\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41916\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__41966\,
            I => \N__41911\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__41963\,
            I => \N__41911\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__41960\,
            I => \N__41908\
        );

    \I__10183\ : InMux
    port map (
            O => \N__41959\,
            I => \N__41905\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__41956\,
            I => \N__41902\
        );

    \I__10181\ : InMux
    port map (
            O => \N__41955\,
            I => \N__41899\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__41952\,
            I => \N__41892\
        );

    \I__10179\ : Span4Mux_v
    port map (
            O => \N__41947\,
            I => \N__41892\
        );

    \I__10178\ : Span4Mux_v
    port map (
            O => \N__41944\,
            I => \N__41892\
        );

    \I__10177\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41887\
        );

    \I__10176\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41887\
        );

    \I__10175\ : InMux
    port map (
            O => \N__41941\,
            I => \N__41884\
        );

    \I__10174\ : Span4Mux_h
    port map (
            O => \N__41938\,
            I => \N__41879\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__41931\,
            I => \N__41874\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41874\
        );

    \I__10171\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41871\
        );

    \I__10170\ : InMux
    port map (
            O => \N__41926\,
            I => \N__41868\
        );

    \I__10169\ : InMux
    port map (
            O => \N__41923\,
            I => \N__41865\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__41920\,
            I => \N__41857\
        );

    \I__10167\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41854\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41851\
        );

    \I__10165\ : Span4Mux_v
    port map (
            O => \N__41911\,
            I => \N__41848\
        );

    \I__10164\ : Span4Mux_s2_h
    port map (
            O => \N__41908\,
            I => \N__41843\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__41905\,
            I => \N__41843\
        );

    \I__10162\ : Span4Mux_h
    port map (
            O => \N__41902\,
            I => \N__41840\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__41899\,
            I => \N__41833\
        );

    \I__10160\ : Sp12to4
    port map (
            O => \N__41892\,
            I => \N__41833\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__41887\,
            I => \N__41833\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__41884\,
            I => \N__41830\
        );

    \I__10157\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41825\
        );

    \I__10156\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41825\
        );

    \I__10155\ : Span4Mux_h
    port map (
            O => \N__41879\,
            I => \N__41820\
        );

    \I__10154\ : Span4Mux_v
    port map (
            O => \N__41874\,
            I => \N__41820\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__41871\,
            I => \N__41813\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41813\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__41865\,
            I => \N__41813\
        );

    \I__10150\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41810\
        );

    \I__10149\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41804\
        );

    \I__10148\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41804\
        );

    \I__10147\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41799\
        );

    \I__10146\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41799\
        );

    \I__10145\ : Span12Mux_v
    port map (
            O => \N__41857\,
            I => \N__41794\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__41854\,
            I => \N__41794\
        );

    \I__10143\ : Span4Mux_h
    port map (
            O => \N__41851\,
            I => \N__41787\
        );

    \I__10142\ : Span4Mux_v
    port map (
            O => \N__41848\,
            I => \N__41787\
        );

    \I__10141\ : Span4Mux_h
    port map (
            O => \N__41843\,
            I => \N__41787\
        );

    \I__10140\ : Sp12to4
    port map (
            O => \N__41840\,
            I => \N__41782\
        );

    \I__10139\ : Span12Mux_s6_h
    port map (
            O => \N__41833\,
            I => \N__41782\
        );

    \I__10138\ : Span4Mux_h
    port map (
            O => \N__41830\,
            I => \N__41779\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__41825\,
            I => \N__41776\
        );

    \I__10136\ : Span4Mux_v
    port map (
            O => \N__41820\,
            I => \N__41769\
        );

    \I__10135\ : Span4Mux_h
    port map (
            O => \N__41813\,
            I => \N__41769\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__41810\,
            I => \N__41769\
        );

    \I__10133\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41766\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__41804\,
            I => \ALU.aluOut_3\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__41799\,
            I => \ALU.aluOut_3\
        );

    \I__10130\ : Odrv12
    port map (
            O => \N__41794\,
            I => \ALU.aluOut_3\
        );

    \I__10129\ : Odrv4
    port map (
            O => \N__41787\,
            I => \ALU.aluOut_3\
        );

    \I__10128\ : Odrv12
    port map (
            O => \N__41782\,
            I => \ALU.aluOut_3\
        );

    \I__10127\ : Odrv4
    port map (
            O => \N__41779\,
            I => \ALU.aluOut_3\
        );

    \I__10126\ : Odrv4
    port map (
            O => \N__41776\,
            I => \ALU.aluOut_3\
        );

    \I__10125\ : Odrv4
    port map (
            O => \N__41769\,
            I => \ALU.aluOut_3\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__41766\,
            I => \ALU.aluOut_3\
        );

    \I__10123\ : CascadeMux
    port map (
            O => \N__41747\,
            I => \N__41744\
        );

    \I__10122\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41741\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__41741\,
            I => \ALU.a_15_m2_ns_1Z0Z_3\
        );

    \I__10120\ : InMux
    port map (
            O => \N__41738\,
            I => \N__41730\
        );

    \I__10119\ : InMux
    port map (
            O => \N__41737\,
            I => \N__41730\
        );

    \I__10118\ : InMux
    port map (
            O => \N__41736\,
            I => \N__41727\
        );

    \I__10117\ : InMux
    port map (
            O => \N__41735\,
            I => \N__41723\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__41730\,
            I => \N__41716\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__41727\,
            I => \N__41713\
        );

    \I__10114\ : InMux
    port map (
            O => \N__41726\,
            I => \N__41710\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__41723\,
            I => \N__41707\
        );

    \I__10112\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41701\
        );

    \I__10111\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41696\
        );

    \I__10110\ : InMux
    port map (
            O => \N__41720\,
            I => \N__41696\
        );

    \I__10109\ : InMux
    port map (
            O => \N__41719\,
            I => \N__41691\
        );

    \I__10108\ : Span4Mux_s2_h
    port map (
            O => \N__41716\,
            I => \N__41688\
        );

    \I__10107\ : Span4Mux_v
    port map (
            O => \N__41713\,
            I => \N__41685\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__41710\,
            I => \N__41682\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__41707\,
            I => \N__41679\
        );

    \I__10104\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41676\
        );

    \I__10103\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41671\
        );

    \I__10102\ : InMux
    port map (
            O => \N__41704\,
            I => \N__41671\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__41701\,
            I => \N__41668\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__41696\,
            I => \N__41664\
        );

    \I__10099\ : InMux
    port map (
            O => \N__41695\,
            I => \N__41659\
        );

    \I__10098\ : InMux
    port map (
            O => \N__41694\,
            I => \N__41659\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__41691\,
            I => \N__41654\
        );

    \I__10096\ : Span4Mux_h
    port map (
            O => \N__41688\,
            I => \N__41654\
        );

    \I__10095\ : Span4Mux_v
    port map (
            O => \N__41685\,
            I => \N__41649\
        );

    \I__10094\ : Span4Mux_v
    port map (
            O => \N__41682\,
            I => \N__41649\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__41679\,
            I => \N__41646\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__41676\,
            I => \N__41641\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__41671\,
            I => \N__41641\
        );

    \I__10090\ : Span12Mux_s6_h
    port map (
            O => \N__41668\,
            I => \N__41638\
        );

    \I__10089\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41635\
        );

    \I__10088\ : Span4Mux_h
    port map (
            O => \N__41664\,
            I => \N__41628\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__41659\,
            I => \N__41628\
        );

    \I__10086\ : Span4Mux_v
    port map (
            O => \N__41654\,
            I => \N__41628\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__41649\,
            I => \N__41625\
        );

    \I__10084\ : Span4Mux_h
    port map (
            O => \N__41646\,
            I => \N__41620\
        );

    \I__10083\ : Span4Mux_v
    port map (
            O => \N__41641\,
            I => \N__41620\
        );

    \I__10082\ : Odrv12
    port map (
            O => \N__41638\,
            I => \ALU.N_237_0\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__41635\,
            I => \ALU.N_237_0\
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__41628\,
            I => \ALU.N_237_0\
        );

    \I__10079\ : Odrv4
    port map (
            O => \N__41625\,
            I => \ALU.N_237_0\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__41620\,
            I => \ALU.N_237_0\
        );

    \I__10077\ : CascadeMux
    port map (
            O => \N__41609\,
            I => \ALU.a_15_m2_3_cascade_\
        );

    \I__10076\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41603\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__41603\,
            I => \N__41600\
        );

    \I__10074\ : Span4Mux_h
    port map (
            O => \N__41600\,
            I => \N__41597\
        );

    \I__10073\ : Span4Mux_h
    port map (
            O => \N__41597\,
            I => \N__41594\
        );

    \I__10072\ : Span4Mux_v
    port map (
            O => \N__41594\,
            I => \N__41591\
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__41591\,
            I => \ALU.lshift_1_3\
        );

    \I__10070\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41585\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__41585\,
            I => \ALU.d_RNI95MLPZ0Z_3\
        );

    \I__10068\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41579\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41576\
        );

    \I__10066\ : Odrv12
    port map (
            O => \N__41576\,
            I => \ALU.mult_3\
        );

    \I__10065\ : InMux
    port map (
            O => \N__41573\,
            I => \N__41570\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__41570\,
            I => \ALU.a_15_m5_3\
        );

    \I__10063\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41564\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__41564\,
            I => \N__41560\
        );

    \I__10061\ : CascadeMux
    port map (
            O => \N__41563\,
            I => \N__41557\
        );

    \I__10060\ : Span4Mux_v
    port map (
            O => \N__41560\,
            I => \N__41554\
        );

    \I__10059\ : InMux
    port map (
            O => \N__41557\,
            I => \N__41551\
        );

    \I__10058\ : Span4Mux_h
    port map (
            O => \N__41554\,
            I => \N__41548\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__41551\,
            I => \N__41545\
        );

    \I__10056\ : Span4Mux_h
    port map (
            O => \N__41548\,
            I => \N__41539\
        );

    \I__10055\ : Span4Mux_v
    port map (
            O => \N__41545\,
            I => \N__41539\
        );

    \I__10054\ : CascadeMux
    port map (
            O => \N__41544\,
            I => \N__41535\
        );

    \I__10053\ : Span4Mux_h
    port map (
            O => \N__41539\,
            I => \N__41531\
        );

    \I__10052\ : InMux
    port map (
            O => \N__41538\,
            I => \N__41526\
        );

    \I__10051\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41526\
        );

    \I__10050\ : InMux
    port map (
            O => \N__41534\,
            I => \N__41523\
        );

    \I__10049\ : Span4Mux_v
    port map (
            O => \N__41531\,
            I => \N__41520\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__41526\,
            I => \N__41517\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__41523\,
            I => \RXbuffer_2\
        );

    \I__10046\ : Odrv4
    port map (
            O => \N__41520\,
            I => \RXbuffer_2\
        );

    \I__10045\ : Odrv4
    port map (
            O => \N__41517\,
            I => \RXbuffer_2\
        );

    \I__10044\ : CascadeMux
    port map (
            O => \N__41510\,
            I => \N__41503\
        );

    \I__10043\ : CascadeMux
    port map (
            O => \N__41509\,
            I => \N__41497\
        );

    \I__10042\ : CascadeMux
    port map (
            O => \N__41508\,
            I => \N__41494\
        );

    \I__10041\ : CascadeMux
    port map (
            O => \N__41507\,
            I => \N__41491\
        );

    \I__10040\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41479\
        );

    \I__10039\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41479\
        );

    \I__10038\ : InMux
    port map (
            O => \N__41502\,
            I => \N__41479\
        );

    \I__10037\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41471\
        );

    \I__10036\ : InMux
    port map (
            O => \N__41500\,
            I => \N__41468\
        );

    \I__10035\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41458\
        );

    \I__10034\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41458\
        );

    \I__10033\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41458\
        );

    \I__10032\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41458\
        );

    \I__10031\ : InMux
    port map (
            O => \N__41489\,
            I => \N__41455\
        );

    \I__10030\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41448\
        );

    \I__10029\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41448\
        );

    \I__10028\ : InMux
    port map (
            O => \N__41486\,
            I => \N__41448\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__41479\,
            I => \N__41445\
        );

    \I__10026\ : CascadeMux
    port map (
            O => \N__41478\,
            I => \N__41442\
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__41477\,
            I => \N__41439\
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__41476\,
            I => \N__41435\
        );

    \I__10023\ : CascadeMux
    port map (
            O => \N__41475\,
            I => \N__41432\
        );

    \I__10022\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41420\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__41471\,
            I => \N__41417\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__41468\,
            I => \N__41414\
        );

    \I__10019\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41410\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__41458\,
            I => \N__41400\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__41455\,
            I => \N__41400\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41400\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__41445\,
            I => \N__41400\
        );

    \I__10014\ : InMux
    port map (
            O => \N__41442\,
            I => \N__41396\
        );

    \I__10013\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41391\
        );

    \I__10012\ : InMux
    port map (
            O => \N__41438\,
            I => \N__41391\
        );

    \I__10011\ : InMux
    port map (
            O => \N__41435\,
            I => \N__41382\
        );

    \I__10010\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41382\
        );

    \I__10009\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41382\
        );

    \I__10008\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41382\
        );

    \I__10007\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41375\
        );

    \I__10006\ : InMux
    port map (
            O => \N__41428\,
            I => \N__41375\
        );

    \I__10005\ : InMux
    port map (
            O => \N__41427\,
            I => \N__41375\
        );

    \I__10004\ : InMux
    port map (
            O => \N__41426\,
            I => \N__41366\
        );

    \I__10003\ : InMux
    port map (
            O => \N__41425\,
            I => \N__41366\
        );

    \I__10002\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41366\
        );

    \I__10001\ : InMux
    port map (
            O => \N__41423\,
            I => \N__41366\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__41420\,
            I => \N__41363\
        );

    \I__9999\ : Span4Mux_h
    port map (
            O => \N__41417\,
            I => \N__41360\
        );

    \I__9998\ : Span4Mux_v
    port map (
            O => \N__41414\,
            I => \N__41356\
        );

    \I__9997\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41353\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__41410\,
            I => \N__41350\
        );

    \I__9995\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41347\
        );

    \I__9994\ : Span4Mux_v
    port map (
            O => \N__41400\,
            I => \N__41344\
        );

    \I__9993\ : InMux
    port map (
            O => \N__41399\,
            I => \N__41341\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__41396\,
            I => \N__41335\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__41391\,
            I => \N__41332\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__41382\,
            I => \N__41329\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__41375\,
            I => \N__41324\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__41366\,
            I => \N__41324\
        );

    \I__9987\ : Span4Mux_h
    port map (
            O => \N__41363\,
            I => \N__41319\
        );

    \I__9986\ : Span4Mux_h
    port map (
            O => \N__41360\,
            I => \N__41319\
        );

    \I__9985\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41316\
        );

    \I__9984\ : Span4Mux_h
    port map (
            O => \N__41356\,
            I => \N__41313\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__41353\,
            I => \N__41306\
        );

    \I__9982\ : Span4Mux_v
    port map (
            O => \N__41350\,
            I => \N__41306\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__41347\,
            I => \N__41306\
        );

    \I__9980\ : Span4Mux_h
    port map (
            O => \N__41344\,
            I => \N__41301\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41301\
        );

    \I__9978\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41294\
        );

    \I__9977\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41294\
        );

    \I__9976\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41294\
        );

    \I__9975\ : Span4Mux_h
    port map (
            O => \N__41335\,
            I => \N__41289\
        );

    \I__9974\ : Span4Mux_h
    port map (
            O => \N__41332\,
            I => \N__41286\
        );

    \I__9973\ : Span4Mux_s3_v
    port map (
            O => \N__41329\,
            I => \N__41281\
        );

    \I__9972\ : Span4Mux_s2_h
    port map (
            O => \N__41324\,
            I => \N__41281\
        );

    \I__9971\ : Span4Mux_v
    port map (
            O => \N__41319\,
            I => \N__41278\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__41316\,
            I => \N__41271\
        );

    \I__9969\ : Span4Mux_v
    port map (
            O => \N__41313\,
            I => \N__41271\
        );

    \I__9968\ : Span4Mux_h
    port map (
            O => \N__41306\,
            I => \N__41271\
        );

    \I__9967\ : Span4Mux_v
    port map (
            O => \N__41301\,
            I => \N__41266\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__41294\,
            I => \N__41266\
        );

    \I__9965\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41261\
        );

    \I__9964\ : InMux
    port map (
            O => \N__41292\,
            I => \N__41261\
        );

    \I__9963\ : Span4Mux_v
    port map (
            O => \N__41289\,
            I => \N__41258\
        );

    \I__9962\ : Span4Mux_v
    port map (
            O => \N__41286\,
            I => \N__41255\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__41281\,
            I => \N__41252\
        );

    \I__9960\ : Span4Mux_v
    port map (
            O => \N__41278\,
            I => \N__41249\
        );

    \I__9959\ : Span4Mux_v
    port map (
            O => \N__41271\,
            I => \N__41244\
        );

    \I__9958\ : Span4Mux_s0_v
    port map (
            O => \N__41266\,
            I => \N__41244\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__41261\,
            I => \testStateZ0Z_1\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__41258\,
            I => \testStateZ0Z_1\
        );

    \I__9955\ : Odrv4
    port map (
            O => \N__41255\,
            I => \testStateZ0Z_1\
        );

    \I__9954\ : Odrv4
    port map (
            O => \N__41252\,
            I => \testStateZ0Z_1\
        );

    \I__9953\ : Odrv4
    port map (
            O => \N__41249\,
            I => \testStateZ0Z_1\
        );

    \I__9952\ : Odrv4
    port map (
            O => \N__41244\,
            I => \testStateZ0Z_1\
        );

    \I__9951\ : InMux
    port map (
            O => \N__41231\,
            I => \N__41227\
        );

    \I__9950\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41224\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41221\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41215\
        );

    \I__9947\ : Span4Mux_v
    port map (
            O => \N__41221\,
            I => \N__41211\
        );

    \I__9946\ : InMux
    port map (
            O => \N__41220\,
            I => \N__41208\
        );

    \I__9945\ : InMux
    port map (
            O => \N__41219\,
            I => \N__41194\
        );

    \I__9944\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41194\
        );

    \I__9943\ : Span4Mux_v
    port map (
            O => \N__41215\,
            I => \N__41191\
        );

    \I__9942\ : InMux
    port map (
            O => \N__41214\,
            I => \N__41188\
        );

    \I__9941\ : Span4Mux_v
    port map (
            O => \N__41211\,
            I => \N__41183\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__41208\,
            I => \N__41183\
        );

    \I__9939\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41178\
        );

    \I__9938\ : InMux
    port map (
            O => \N__41206\,
            I => \N__41178\
        );

    \I__9937\ : InMux
    port map (
            O => \N__41205\,
            I => \N__41163\
        );

    \I__9936\ : InMux
    port map (
            O => \N__41204\,
            I => \N__41163\
        );

    \I__9935\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41163\
        );

    \I__9934\ : InMux
    port map (
            O => \N__41202\,
            I => \N__41163\
        );

    \I__9933\ : InMux
    port map (
            O => \N__41201\,
            I => \N__41163\
        );

    \I__9932\ : InMux
    port map (
            O => \N__41200\,
            I => \N__41163\
        );

    \I__9931\ : InMux
    port map (
            O => \N__41199\,
            I => \N__41163\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__41194\,
            I => \N__41160\
        );

    \I__9929\ : Sp12to4
    port map (
            O => \N__41191\,
            I => \N__41156\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41153\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__41183\,
            I => \N__41150\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__41178\,
            I => \N__41147\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__41163\,
            I => \N__41142\
        );

    \I__9924\ : Sp12to4
    port map (
            O => \N__41160\,
            I => \N__41142\
        );

    \I__9923\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41139\
        );

    \I__9922\ : Span12Mux_v
    port map (
            O => \N__41156\,
            I => \N__41136\
        );

    \I__9921\ : Span4Mux_v
    port map (
            O => \N__41153\,
            I => \N__41133\
        );

    \I__9920\ : Span4Mux_h
    port map (
            O => \N__41150\,
            I => \N__41128\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__41147\,
            I => \N__41128\
        );

    \I__9918\ : Span12Mux_s5_h
    port map (
            O => \N__41142\,
            I => \N__41123\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__41139\,
            I => \N__41123\
        );

    \I__9916\ : Odrv12
    port map (
            O => \N__41136\,
            I => \ALU.N_58_0\
        );

    \I__9915\ : Odrv4
    port map (
            O => \N__41133\,
            I => \ALU.N_58_0\
        );

    \I__9914\ : Odrv4
    port map (
            O => \N__41128\,
            I => \ALU.N_58_0\
        );

    \I__9913\ : Odrv12
    port map (
            O => \N__41123\,
            I => \ALU.N_58_0\
        );

    \I__9912\ : InMux
    port map (
            O => \N__41114\,
            I => \N__41109\
        );

    \I__9911\ : CascadeMux
    port map (
            O => \N__41113\,
            I => \N__41104\
        );

    \I__9910\ : InMux
    port map (
            O => \N__41112\,
            I => \N__41101\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__41109\,
            I => \N__41098\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__41108\,
            I => \N__41095\
        );

    \I__9907\ : InMux
    port map (
            O => \N__41107\,
            I => \N__41090\
        );

    \I__9906\ : InMux
    port map (
            O => \N__41104\,
            I => \N__41090\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__41101\,
            I => \N__41087\
        );

    \I__9904\ : Span4Mux_v
    port map (
            O => \N__41098\,
            I => \N__41084\
        );

    \I__9903\ : InMux
    port map (
            O => \N__41095\,
            I => \N__41081\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__41090\,
            I => \N__41078\
        );

    \I__9901\ : Span12Mux_s8_h
    port map (
            O => \N__41087\,
            I => \N__41075\
        );

    \I__9900\ : Span4Mux_h
    port map (
            O => \N__41084\,
            I => \N__41072\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__41081\,
            I => \testWordZ0Z_10\
        );

    \I__9898\ : Odrv4
    port map (
            O => \N__41078\,
            I => \testWordZ0Z_10\
        );

    \I__9897\ : Odrv12
    port map (
            O => \N__41075\,
            I => \testWordZ0Z_10\
        );

    \I__9896\ : Odrv4
    port map (
            O => \N__41072\,
            I => \testWordZ0Z_10\
        );

    \I__9895\ : CEMux
    port map (
            O => \N__41063\,
            I => \N__41027\
        );

    \I__9894\ : CEMux
    port map (
            O => \N__41062\,
            I => \N__41027\
        );

    \I__9893\ : CEMux
    port map (
            O => \N__41061\,
            I => \N__41027\
        );

    \I__9892\ : CEMux
    port map (
            O => \N__41060\,
            I => \N__41027\
        );

    \I__9891\ : CEMux
    port map (
            O => \N__41059\,
            I => \N__41027\
        );

    \I__9890\ : CEMux
    port map (
            O => \N__41058\,
            I => \N__41027\
        );

    \I__9889\ : CEMux
    port map (
            O => \N__41057\,
            I => \N__41027\
        );

    \I__9888\ : CEMux
    port map (
            O => \N__41056\,
            I => \N__41027\
        );

    \I__9887\ : CEMux
    port map (
            O => \N__41055\,
            I => \N__41027\
        );

    \I__9886\ : CEMux
    port map (
            O => \N__41054\,
            I => \N__41027\
        );

    \I__9885\ : CEMux
    port map (
            O => \N__41053\,
            I => \N__41027\
        );

    \I__9884\ : CEMux
    port map (
            O => \N__41052\,
            I => \N__41027\
        );

    \I__9883\ : GlobalMux
    port map (
            O => \N__41027\,
            I => \N__41024\
        );

    \I__9882\ : gio2CtrlBuf
    port map (
            O => \N__41024\,
            I => \testState_i_g_2\
        );

    \I__9881\ : InMux
    port map (
            O => \N__41021\,
            I => \N__41018\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__9879\ : Odrv12
    port map (
            O => \N__41015\,
            I => \ALU.un9_addsub_cry_0_c_RNI2UZ0Z096\
        );

    \I__9878\ : InMux
    port map (
            O => \N__41012\,
            I => \N__41009\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__41009\,
            I => \N__41006\
        );

    \I__9876\ : Span12Mux_h
    port map (
            O => \N__41006\,
            I => \N__41003\
        );

    \I__9875\ : Odrv12
    port map (
            O => \N__41003\,
            I => \ALU.un2_addsub_cry_0_c_RNI5MA0EZ0\
        );

    \I__9874\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40995\
        );

    \I__9873\ : InMux
    port map (
            O => \N__40999\,
            I => \N__40991\
        );

    \I__9872\ : InMux
    port map (
            O => \N__40998\,
            I => \N__40988\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__40995\,
            I => \N__40985\
        );

    \I__9870\ : InMux
    port map (
            O => \N__40994\,
            I => \N__40982\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__40991\,
            I => \N__40976\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__40988\,
            I => \N__40969\
        );

    \I__9867\ : Span4Mux_h
    port map (
            O => \N__40985\,
            I => \N__40969\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__40982\,
            I => \N__40969\
        );

    \I__9865\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40966\
        );

    \I__9864\ : InMux
    port map (
            O => \N__40980\,
            I => \N__40963\
        );

    \I__9863\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40960\
        );

    \I__9862\ : Span4Mux_h
    port map (
            O => \N__40976\,
            I => \N__40956\
        );

    \I__9861\ : Span4Mux_v
    port map (
            O => \N__40969\,
            I => \N__40951\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__40966\,
            I => \N__40951\
        );

    \I__9859\ : LocalMux
    port map (
            O => \N__40963\,
            I => \N__40946\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__40960\,
            I => \N__40946\
        );

    \I__9857\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40943\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__40956\,
            I => \N__40940\
        );

    \I__9855\ : Span4Mux_h
    port map (
            O => \N__40951\,
            I => \N__40937\
        );

    \I__9854\ : Span4Mux_v
    port map (
            O => \N__40946\,
            I => \N__40932\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__40943\,
            I => \N__40932\
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__40940\,
            I => \ALU.un9_addsub_cry_0_c_RNIEMTLKZ0\
        );

    \I__9851\ : Odrv4
    port map (
            O => \N__40937\,
            I => \ALU.un9_addsub_cry_0_c_RNIEMTLKZ0\
        );

    \I__9850\ : Odrv4
    port map (
            O => \N__40932\,
            I => \ALU.un9_addsub_cry_0_c_RNIEMTLKZ0\
        );

    \I__9849\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40922\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__40922\,
            I => \N__40919\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__40919\,
            I => \ALU.un9_addsub_cry_1_c_RNI6TDZ0Z17\
        );

    \I__9846\ : InMux
    port map (
            O => \N__40916\,
            I => \N__40913\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__40913\,
            I => \N__40910\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__40910\,
            I => \N__40907\
        );

    \I__9843\ : Sp12to4
    port map (
            O => \N__40907\,
            I => \N__40904\
        );

    \I__9842\ : Odrv12
    port map (
            O => \N__40904\,
            I => \ALU.un2_addsub_cry_1_c_RNI966GEZ0\
        );

    \I__9841\ : InMux
    port map (
            O => \N__40901\,
            I => \N__40898\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__40898\,
            I => \N__40895\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__40895\,
            I => \ALU.un9_addsub_cry_2_c_RNIA3LGZ0Z7\
        );

    \I__9838\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40889\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__40889\,
            I => \N__40886\
        );

    \I__9836\ : Span4Mux_h
    port map (
            O => \N__40886\,
            I => \N__40883\
        );

    \I__9835\ : Span4Mux_h
    port map (
            O => \N__40883\,
            I => \N__40880\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__40880\,
            I => \ALU.un2_addsub_cry_2_c_RNI5IV5FZ0\
        );

    \I__9833\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40874\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__40874\,
            I => \N__40871\
        );

    \I__9831\ : Span4Mux_v
    port map (
            O => \N__40871\,
            I => \N__40868\
        );

    \I__9830\ : Span4Mux_h
    port map (
            O => \N__40868\,
            I => \N__40865\
        );

    \I__9829\ : Odrv4
    port map (
            O => \N__40865\,
            I => \ALU.un2_addsub_cry_3_c_RNIOGGJGZ0\
        );

    \I__9828\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40859\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__40859\,
            I => \N__40856\
        );

    \I__9826\ : Odrv4
    port map (
            O => \N__40856\,
            I => \ALU.un9_addsub_cry_3_c_RNI525RZ0Z7\
        );

    \I__9825\ : InMux
    port map (
            O => \N__40853\,
            I => \N__40850\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__40850\,
            I => \N__40844\
        );

    \I__9823\ : InMux
    port map (
            O => \N__40849\,
            I => \N__40841\
        );

    \I__9822\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40836\
        );

    \I__9821\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40836\
        );

    \I__9820\ : Span4Mux_h
    port map (
            O => \N__40844\,
            I => \N__40833\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__40841\,
            I => \N__40830\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__40836\,
            I => \N__40827\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__40833\,
            I => \N__40823\
        );

    \I__9816\ : Span4Mux_h
    port map (
            O => \N__40830\,
            I => \N__40820\
        );

    \I__9815\ : Span4Mux_h
    port map (
            O => \N__40827\,
            I => \N__40817\
        );

    \I__9814\ : InMux
    port map (
            O => \N__40826\,
            I => \N__40814\
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__40823\,
            I => \ALU.N_180_0\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__40820\,
            I => \ALU.N_180_0\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__40817\,
            I => \ALU.N_180_0\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__40814\,
            I => \ALU.N_180_0\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__40805\,
            I => \N__40802\
        );

    \I__9808\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40799\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__40799\,
            I => \N__40796\
        );

    \I__9806\ : Span4Mux_v
    port map (
            O => \N__40796\,
            I => \N__40793\
        );

    \I__9805\ : Sp12to4
    port map (
            O => \N__40793\,
            I => \N__40790\
        );

    \I__9804\ : Odrv12
    port map (
            O => \N__40790\,
            I => \ALU.d_RNIFKNTEZ0Z_12\
        );

    \I__9803\ : InMux
    port map (
            O => \N__40787\,
            I => \N__40784\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__40784\,
            I => \N__40781\
        );

    \I__9801\ : Span4Mux_h
    port map (
            O => \N__40781\,
            I => \N__40778\
        );

    \I__9800\ : Odrv4
    port map (
            O => \N__40778\,
            I => \ALU.un9_addsub_cry_11_c_RNI10BQKZ0\
        );

    \I__9799\ : InMux
    port map (
            O => \N__40775\,
            I => \ALU.un9_addsub_cry_11\
        );

    \I__9798\ : CascadeMux
    port map (
            O => \N__40772\,
            I => \N__40769\
        );

    \I__9797\ : InMux
    port map (
            O => \N__40769\,
            I => \N__40760\
        );

    \I__9796\ : InMux
    port map (
            O => \N__40768\,
            I => \N__40753\
        );

    \I__9795\ : InMux
    port map (
            O => \N__40767\,
            I => \N__40753\
        );

    \I__9794\ : InMux
    port map (
            O => \N__40766\,
            I => \N__40753\
        );

    \I__9793\ : InMux
    port map (
            O => \N__40765\,
            I => \N__40748\
        );

    \I__9792\ : CascadeMux
    port map (
            O => \N__40764\,
            I => \N__40743\
        );

    \I__9791\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40740\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__40760\,
            I => \N__40737\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__40753\,
            I => \N__40734\
        );

    \I__9788\ : InMux
    port map (
            O => \N__40752\,
            I => \N__40729\
        );

    \I__9787\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40729\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__40748\,
            I => \N__40726\
        );

    \I__9785\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40723\
        );

    \I__9784\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40718\
        );

    \I__9783\ : InMux
    port map (
            O => \N__40743\,
            I => \N__40718\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__40740\,
            I => \N__40715\
        );

    \I__9781\ : Span4Mux_s3_h
    port map (
            O => \N__40737\,
            I => \N__40712\
        );

    \I__9780\ : Span4Mux_v
    port map (
            O => \N__40734\,
            I => \N__40708\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__40729\,
            I => \N__40701\
        );

    \I__9778\ : Span4Mux_h
    port map (
            O => \N__40726\,
            I => \N__40701\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__40723\,
            I => \N__40701\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__40718\,
            I => \N__40696\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__40715\,
            I => \N__40696\
        );

    \I__9774\ : Span4Mux_h
    port map (
            O => \N__40712\,
            I => \N__40693\
        );

    \I__9773\ : InMux
    port map (
            O => \N__40711\,
            I => \N__40690\
        );

    \I__9772\ : Span4Mux_h
    port map (
            O => \N__40708\,
            I => \N__40685\
        );

    \I__9771\ : Span4Mux_v
    port map (
            O => \N__40701\,
            I => \N__40685\
        );

    \I__9770\ : Span4Mux_h
    port map (
            O => \N__40696\,
            I => \N__40682\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__40693\,
            I => \N__40679\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__40690\,
            I => \N__40674\
        );

    \I__9767\ : Span4Mux_h
    port map (
            O => \N__40685\,
            I => \N__40674\
        );

    \I__9766\ : Span4Mux_h
    port map (
            O => \N__40682\,
            I => \N__40671\
        );

    \I__9765\ : Odrv4
    port map (
            O => \N__40679\,
            I => \ALU.aluOut_13\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__40674\,
            I => \ALU.aluOut_13\
        );

    \I__9763\ : Odrv4
    port map (
            O => \N__40671\,
            I => \ALU.aluOut_13\
        );

    \I__9762\ : CascadeMux
    port map (
            O => \N__40664\,
            I => \N__40661\
        );

    \I__9761\ : InMux
    port map (
            O => \N__40661\,
            I => \N__40658\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40655\
        );

    \I__9759\ : Span4Mux_v
    port map (
            O => \N__40655\,
            I => \N__40652\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__40652\,
            I => \ALU.N_177_0_i\
        );

    \I__9757\ : InMux
    port map (
            O => \N__40649\,
            I => \N__40646\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__40646\,
            I => \N__40643\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__40643\,
            I => \N__40640\
        );

    \I__9754\ : Odrv4
    port map (
            O => \N__40640\,
            I => \ALU.un9_addsub_cry_12_c_RNIBB5QZ0Z9\
        );

    \I__9753\ : InMux
    port map (
            O => \N__40637\,
            I => \ALU.un9_addsub_cry_12\
        );

    \I__9752\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40631\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__40631\,
            I => \N__40628\
        );

    \I__9750\ : Span4Mux_h
    port map (
            O => \N__40628\,
            I => \N__40623\
        );

    \I__9749\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40620\
        );

    \I__9748\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40611\
        );

    \I__9747\ : Span4Mux_v
    port map (
            O => \N__40623\,
            I => \N__40606\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__40620\,
            I => \N__40606\
        );

    \I__9745\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40601\
        );

    \I__9744\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40601\
        );

    \I__9743\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40596\
        );

    \I__9742\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40593\
        );

    \I__9741\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40590\
        );

    \I__9740\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40587\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__40611\,
            I => \N__40584\
        );

    \I__9738\ : Span4Mux_h
    port map (
            O => \N__40606\,
            I => \N__40579\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__40601\,
            I => \N__40579\
        );

    \I__9736\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40574\
        );

    \I__9735\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40574\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__40596\,
            I => \ALU.aluOut_14\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__40593\,
            I => \ALU.aluOut_14\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__40590\,
            I => \ALU.aluOut_14\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__40587\,
            I => \ALU.aluOut_14\
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__40584\,
            I => \ALU.aluOut_14\
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__40579\,
            I => \ALU.aluOut_14\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__40574\,
            I => \ALU.aluOut_14\
        );

    \I__9727\ : CascadeMux
    port map (
            O => \N__40559\,
            I => \N__40556\
        );

    \I__9726\ : InMux
    port map (
            O => \N__40556\,
            I => \N__40553\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__40553\,
            I => \N__40550\
        );

    \I__9724\ : Span4Mux_v
    port map (
            O => \N__40550\,
            I => \N__40547\
        );

    \I__9723\ : Span4Mux_h
    port map (
            O => \N__40547\,
            I => \N__40544\
        );

    \I__9722\ : Span4Mux_h
    port map (
            O => \N__40544\,
            I => \N__40541\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__40541\,
            I => \ALU.N_171_0_i\
        );

    \I__9720\ : InMux
    port map (
            O => \N__40538\,
            I => \N__40535\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__40535\,
            I => \N__40532\
        );

    \I__9718\ : Span4Mux_h
    port map (
            O => \N__40532\,
            I => \N__40529\
        );

    \I__9717\ : Odrv4
    port map (
            O => \N__40529\,
            I => \ALU.un9_addsub_cry_13_c_RNI4JGFZ0Z9\
        );

    \I__9716\ : InMux
    port map (
            O => \N__40526\,
            I => \ALU.un9_addsub_cry_13\
        );

    \I__9715\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40520\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__40520\,
            I => \N__40517\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__40517\,
            I => \N__40514\
        );

    \I__9712\ : Sp12to4
    port map (
            O => \N__40514\,
            I => \N__40511\
        );

    \I__9711\ : Odrv12
    port map (
            O => \N__40511\,
            I => \ALU.un9_addsub_axb_15\
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__40508\,
            I => \N__40505\
        );

    \I__9709\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40502\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__40502\,
            I => \N__40499\
        );

    \I__9707\ : Span4Mux_v
    port map (
            O => \N__40499\,
            I => \N__40496\
        );

    \I__9706\ : Sp12to4
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__9705\ : Odrv12
    port map (
            O => \N__40493\,
            I => \ALU.un2_addsub_cry_14_c_RNINOKZ0Z69\
        );

    \I__9704\ : InMux
    port map (
            O => \N__40490\,
            I => \ALU.un9_addsub_cry_14\
        );

    \I__9703\ : InMux
    port map (
            O => \N__40487\,
            I => \N__40484\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__40484\,
            I => \ALU.un9_addsub_cry_14_c_RNIS374JZ0\
        );

    \I__9701\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40478\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__40478\,
            I => \N__40475\
        );

    \I__9699\ : Span4Mux_v
    port map (
            O => \N__40475\,
            I => \N__40472\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__40472\,
            I => \N__40469\
        );

    \I__9697\ : Odrv4
    port map (
            O => \N__40469\,
            I => \ALU.c_RNIA9V4LZ0Z_15\
        );

    \I__9696\ : InMux
    port map (
            O => \N__40466\,
            I => \N__40463\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__40463\,
            I => \N__40460\
        );

    \I__9694\ : Span12Mux_v
    port map (
            O => \N__40460\,
            I => \N__40457\
        );

    \I__9693\ : Odrv12
    port map (
            O => \N__40457\,
            I => \ALU.d_RNI9DPVUZ0Z_6\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__40454\,
            I => \ALU.rshift_3_cascade_\
        );

    \I__9691\ : InMux
    port map (
            O => \N__40451\,
            I => \N__40448\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__40448\,
            I => \N__40445\
        );

    \I__9689\ : Span12Mux_s9_v
    port map (
            O => \N__40445\,
            I => \N__40442\
        );

    \I__9688\ : Span12Mux_h
    port map (
            O => \N__40442\,
            I => \N__40439\
        );

    \I__9687\ : Odrv12
    port map (
            O => \N__40439\,
            I => \ALU.N_293_0\
        );

    \I__9686\ : CascadeMux
    port map (
            O => \N__40436\,
            I => \ALU.d_RNI3V2CP1Z0Z_3_cascade_\
        );

    \I__9685\ : CascadeMux
    port map (
            O => \N__40433\,
            I => \N__40420\
        );

    \I__9684\ : InMux
    port map (
            O => \N__40432\,
            I => \N__40414\
        );

    \I__9683\ : InMux
    port map (
            O => \N__40431\,
            I => \N__40414\
        );

    \I__9682\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40411\
        );

    \I__9681\ : InMux
    port map (
            O => \N__40429\,
            I => \N__40406\
        );

    \I__9680\ : InMux
    port map (
            O => \N__40428\,
            I => \N__40403\
        );

    \I__9679\ : InMux
    port map (
            O => \N__40427\,
            I => \N__40398\
        );

    \I__9678\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40395\
        );

    \I__9677\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40392\
        );

    \I__9676\ : InMux
    port map (
            O => \N__40424\,
            I => \N__40385\
        );

    \I__9675\ : InMux
    port map (
            O => \N__40423\,
            I => \N__40380\
        );

    \I__9674\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40380\
        );

    \I__9673\ : InMux
    port map (
            O => \N__40419\,
            I => \N__40377\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__40414\,
            I => \N__40372\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__40411\,
            I => \N__40372\
        );

    \I__9670\ : InMux
    port map (
            O => \N__40410\,
            I => \N__40369\
        );

    \I__9669\ : CascadeMux
    port map (
            O => \N__40409\,
            I => \N__40363\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__40406\,
            I => \N__40357\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__40403\,
            I => \N__40357\
        );

    \I__9666\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40354\
        );

    \I__9665\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40351\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__40398\,
            I => \N__40348\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__40395\,
            I => \N__40343\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__40392\,
            I => \N__40343\
        );

    \I__9661\ : InMux
    port map (
            O => \N__40391\,
            I => \N__40340\
        );

    \I__9660\ : InMux
    port map (
            O => \N__40390\,
            I => \N__40337\
        );

    \I__9659\ : InMux
    port map (
            O => \N__40389\,
            I => \N__40332\
        );

    \I__9658\ : InMux
    port map (
            O => \N__40388\,
            I => \N__40332\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__40385\,
            I => \N__40329\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__40380\,
            I => \N__40326\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__40377\,
            I => \N__40319\
        );

    \I__9654\ : Span4Mux_v
    port map (
            O => \N__40372\,
            I => \N__40319\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__40369\,
            I => \N__40319\
        );

    \I__9652\ : InMux
    port map (
            O => \N__40368\,
            I => \N__40316\
        );

    \I__9651\ : InMux
    port map (
            O => \N__40367\,
            I => \N__40311\
        );

    \I__9650\ : InMux
    port map (
            O => \N__40366\,
            I => \N__40311\
        );

    \I__9649\ : InMux
    port map (
            O => \N__40363\,
            I => \N__40306\
        );

    \I__9648\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40306\
        );

    \I__9647\ : Span12Mux_h
    port map (
            O => \N__40357\,
            I => \N__40301\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__40354\,
            I => \N__40301\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__40351\,
            I => \N__40298\
        );

    \I__9644\ : Span4Mux_v
    port map (
            O => \N__40348\,
            I => \N__40293\
        );

    \I__9643\ : Span4Mux_v
    port map (
            O => \N__40343\,
            I => \N__40293\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__40340\,
            I => \N__40288\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40283\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40283\
        );

    \I__9639\ : Span4Mux_v
    port map (
            O => \N__40329\,
            I => \N__40278\
        );

    \I__9638\ : Span4Mux_h
    port map (
            O => \N__40326\,
            I => \N__40278\
        );

    \I__9637\ : Span4Mux_v
    port map (
            O => \N__40319\,
            I => \N__40271\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__40316\,
            I => \N__40271\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__40311\,
            I => \N__40266\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__40306\,
            I => \N__40266\
        );

    \I__9633\ : Span12Mux_v
    port map (
            O => \N__40301\,
            I => \N__40263\
        );

    \I__9632\ : Span12Mux_v
    port map (
            O => \N__40298\,
            I => \N__40258\
        );

    \I__9631\ : Sp12to4
    port map (
            O => \N__40293\,
            I => \N__40258\
        );

    \I__9630\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40253\
        );

    \I__9629\ : InMux
    port map (
            O => \N__40291\,
            I => \N__40253\
        );

    \I__9628\ : Span12Mux_h
    port map (
            O => \N__40288\,
            I => \N__40246\
        );

    \I__9627\ : Span12Mux_s5_h
    port map (
            O => \N__40283\,
            I => \N__40246\
        );

    \I__9626\ : Sp12to4
    port map (
            O => \N__40278\,
            I => \N__40246\
        );

    \I__9625\ : InMux
    port map (
            O => \N__40277\,
            I => \N__40241\
        );

    \I__9624\ : InMux
    port map (
            O => \N__40276\,
            I => \N__40241\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__40271\,
            I => \N__40236\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__40266\,
            I => \N__40236\
        );

    \I__9621\ : Odrv12
    port map (
            O => \N__40263\,
            I => \ALU.aluOut_5\
        );

    \I__9620\ : Odrv12
    port map (
            O => \N__40258\,
            I => \ALU.aluOut_5\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__40253\,
            I => \ALU.aluOut_5\
        );

    \I__9618\ : Odrv12
    port map (
            O => \N__40246\,
            I => \ALU.aluOut_5\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__40241\,
            I => \ALU.aluOut_5\
        );

    \I__9616\ : Odrv4
    port map (
            O => \N__40236\,
            I => \ALU.aluOut_5\
        );

    \I__9615\ : CascadeMux
    port map (
            O => \N__40223\,
            I => \N__40220\
        );

    \I__9614\ : InMux
    port map (
            O => \N__40220\,
            I => \N__40217\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__40217\,
            I => \N__40214\
        );

    \I__9612\ : Span4Mux_h
    port map (
            O => \N__40214\,
            I => \N__40211\
        );

    \I__9611\ : Span4Mux_v
    port map (
            O => \N__40211\,
            I => \N__40208\
        );

    \I__9610\ : Span4Mux_v
    port map (
            O => \N__40208\,
            I => \N__40205\
        );

    \I__9609\ : Span4Mux_h
    port map (
            O => \N__40205\,
            I => \N__40202\
        );

    \I__9608\ : Span4Mux_h
    port map (
            O => \N__40202\,
            I => \N__40199\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__40199\,
            I => \ALU.N_225_0_i\
        );

    \I__9606\ : InMux
    port map (
            O => \N__40196\,
            I => \ALU.un9_addsub_cry_4\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__40193\,
            I => \N__40190\
        );

    \I__9604\ : InMux
    port map (
            O => \N__40190\,
            I => \N__40187\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__40187\,
            I => \N__40184\
        );

    \I__9602\ : Span4Mux_h
    port map (
            O => \N__40184\,
            I => \N__40181\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__40181\,
            I => \N__40178\
        );

    \I__9600\ : Odrv4
    port map (
            O => \N__40178\,
            I => \ALU.N_219_0_i\
        );

    \I__9599\ : InMux
    port map (
            O => \N__40175\,
            I => \ALU.un9_addsub_cry_5\
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__40172\,
            I => \N__40169\
        );

    \I__9597\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40166\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__40166\,
            I => \N__40163\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__40163\,
            I => \N__40160\
        );

    \I__9594\ : Span4Mux_v
    port map (
            O => \N__40160\,
            I => \N__40157\
        );

    \I__9593\ : Span4Mux_v
    port map (
            O => \N__40157\,
            I => \N__40154\
        );

    \I__9592\ : Span4Mux_h
    port map (
            O => \N__40154\,
            I => \N__40151\
        );

    \I__9591\ : Span4Mux_h
    port map (
            O => \N__40151\,
            I => \N__40148\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__40148\,
            I => \ALU.N_213_0_i\
        );

    \I__9589\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40142\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__40142\,
            I => \N__40139\
        );

    \I__9587\ : Span4Mux_h
    port map (
            O => \N__40139\,
            I => \N__40136\
        );

    \I__9586\ : Span4Mux_h
    port map (
            O => \N__40136\,
            I => \N__40133\
        );

    \I__9585\ : Span4Mux_v
    port map (
            O => \N__40133\,
            I => \N__40130\
        );

    \I__9584\ : Span4Mux_v
    port map (
            O => \N__40130\,
            I => \N__40127\
        );

    \I__9583\ : Odrv4
    port map (
            O => \N__40127\,
            I => \ALU.un9_addsub_cry_6_c_RNI2EFHZ0Z8\
        );

    \I__9582\ : InMux
    port map (
            O => \N__40124\,
            I => \ALU.un9_addsub_cry_6\
        );

    \I__9581\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40116\
        );

    \I__9580\ : CascadeMux
    port map (
            O => \N__40120\,
            I => \N__40113\
        );

    \I__9579\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40108\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__40116\,
            I => \N__40104\
        );

    \I__9577\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40099\
        );

    \I__9576\ : CascadeMux
    port map (
            O => \N__40112\,
            I => \N__40095\
        );

    \I__9575\ : InMux
    port map (
            O => \N__40111\,
            I => \N__40090\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__40108\,
            I => \N__40087\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__40107\,
            I => \N__40076\
        );

    \I__9572\ : Span4Mux_v
    port map (
            O => \N__40104\,
            I => \N__40072\
        );

    \I__9571\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40066\
        );

    \I__9570\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40063\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__40099\,
            I => \N__40060\
        );

    \I__9568\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40057\
        );

    \I__9567\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40053\
        );

    \I__9566\ : InMux
    port map (
            O => \N__40094\,
            I => \N__40050\
        );

    \I__9565\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40047\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__40090\,
            I => \N__40040\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__40087\,
            I => \N__40037\
        );

    \I__9562\ : InMux
    port map (
            O => \N__40086\,
            I => \N__40032\
        );

    \I__9561\ : InMux
    port map (
            O => \N__40085\,
            I => \N__40032\
        );

    \I__9560\ : InMux
    port map (
            O => \N__40084\,
            I => \N__40029\
        );

    \I__9559\ : InMux
    port map (
            O => \N__40083\,
            I => \N__40022\
        );

    \I__9558\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40022\
        );

    \I__9557\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40022\
        );

    \I__9556\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40015\
        );

    \I__9555\ : InMux
    port map (
            O => \N__40079\,
            I => \N__40015\
        );

    \I__9554\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40015\
        );

    \I__9553\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40012\
        );

    \I__9552\ : Span4Mux_h
    port map (
            O => \N__40072\,
            I => \N__40009\
        );

    \I__9551\ : InMux
    port map (
            O => \N__40071\,
            I => \N__40006\
        );

    \I__9550\ : InMux
    port map (
            O => \N__40070\,
            I => \N__40001\
        );

    \I__9549\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40001\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__40066\,
            I => \N__39996\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__40063\,
            I => \N__39996\
        );

    \I__9546\ : Span4Mux_v
    port map (
            O => \N__40060\,
            I => \N__39993\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__40057\,
            I => \N__39990\
        );

    \I__9544\ : InMux
    port map (
            O => \N__40056\,
            I => \N__39987\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__40053\,
            I => \N__39984\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__40050\,
            I => \N__39979\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__40047\,
            I => \N__39979\
        );

    \I__9540\ : InMux
    port map (
            O => \N__40046\,
            I => \N__39976\
        );

    \I__9539\ : InMux
    port map (
            O => \N__40045\,
            I => \N__39971\
        );

    \I__9538\ : InMux
    port map (
            O => \N__40044\,
            I => \N__39971\
        );

    \I__9537\ : InMux
    port map (
            O => \N__40043\,
            I => \N__39968\
        );

    \I__9536\ : Span4Mux_v
    port map (
            O => \N__40040\,
            I => \N__39963\
        );

    \I__9535\ : Span4Mux_h
    port map (
            O => \N__40037\,
            I => \N__39963\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__40032\,
            I => \N__39960\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__40029\,
            I => \N__39953\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__40022\,
            I => \N__39953\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__40015\,
            I => \N__39953\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__40012\,
            I => \N__39950\
        );

    \I__9529\ : Span4Mux_h
    port map (
            O => \N__40009\,
            I => \N__39943\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__40006\,
            I => \N__39943\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__40001\,
            I => \N__39943\
        );

    \I__9526\ : Span4Mux_v
    port map (
            O => \N__39996\,
            I => \N__39940\
        );

    \I__9525\ : Span4Mux_h
    port map (
            O => \N__39993\,
            I => \N__39933\
        );

    \I__9524\ : Span4Mux_v
    port map (
            O => \N__39990\,
            I => \N__39933\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__39987\,
            I => \N__39933\
        );

    \I__9522\ : Span4Mux_s1_h
    port map (
            O => \N__39984\,
            I => \N__39928\
        );

    \I__9521\ : Span4Mux_v
    port map (
            O => \N__39979\,
            I => \N__39928\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__39976\,
            I => \N__39923\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__39971\,
            I => \N__39923\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__39968\,
            I => \N__39920\
        );

    \I__9517\ : Span4Mux_v
    port map (
            O => \N__39963\,
            I => \N__39913\
        );

    \I__9516\ : Span4Mux_v
    port map (
            O => \N__39960\,
            I => \N__39913\
        );

    \I__9515\ : Span4Mux_v
    port map (
            O => \N__39953\,
            I => \N__39913\
        );

    \I__9514\ : Span4Mux_v
    port map (
            O => \N__39950\,
            I => \N__39904\
        );

    \I__9513\ : Span4Mux_v
    port map (
            O => \N__39943\,
            I => \N__39904\
        );

    \I__9512\ : Span4Mux_h
    port map (
            O => \N__39940\,
            I => \N__39904\
        );

    \I__9511\ : Span4Mux_v
    port map (
            O => \N__39933\,
            I => \N__39904\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__39928\,
            I => \N__39899\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__39923\,
            I => \N__39899\
        );

    \I__9508\ : Odrv4
    port map (
            O => \N__39920\,
            I => \ALU.aluOut_8\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__39913\,
            I => \ALU.aluOut_8\
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__39904\,
            I => \ALU.aluOut_8\
        );

    \I__9505\ : Odrv4
    port map (
            O => \N__39899\,
            I => \ALU.aluOut_8\
        );

    \I__9504\ : CascadeMux
    port map (
            O => \N__39890\,
            I => \N__39887\
        );

    \I__9503\ : InMux
    port map (
            O => \N__39887\,
            I => \N__39884\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__39884\,
            I => \N__39881\
        );

    \I__9501\ : Span12Mux_h
    port map (
            O => \N__39881\,
            I => \N__39878\
        );

    \I__9500\ : Odrv12
    port map (
            O => \N__39878\,
            I => \ALU.N_201_0_i\
        );

    \I__9499\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39872\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__39872\,
            I => \N__39869\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__39869\,
            I => \N__39866\
        );

    \I__9496\ : Odrv4
    port map (
            O => \N__39866\,
            I => \ALU.un9_addsub_cry_7_c_RNIU7FZ0Z18\
        );

    \I__9495\ : InMux
    port map (
            O => \N__39863\,
            I => \bfn_13_8_0_\
        );

    \I__9494\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39856\
        );

    \I__9493\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39844\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__39856\,
            I => \N__39841\
        );

    \I__9491\ : InMux
    port map (
            O => \N__39855\,
            I => \N__39838\
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__39854\,
            I => \N__39833\
        );

    \I__9489\ : InMux
    port map (
            O => \N__39853\,
            I => \N__39829\
        );

    \I__9488\ : CascadeMux
    port map (
            O => \N__39852\,
            I => \N__39826\
        );

    \I__9487\ : InMux
    port map (
            O => \N__39851\,
            I => \N__39822\
        );

    \I__9486\ : InMux
    port map (
            O => \N__39850\,
            I => \N__39818\
        );

    \I__9485\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39815\
        );

    \I__9484\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39809\
        );

    \I__9483\ : InMux
    port map (
            O => \N__39847\,
            I => \N__39809\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__39844\,
            I => \N__39804\
        );

    \I__9481\ : Span4Mux_h
    port map (
            O => \N__39841\,
            I => \N__39799\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39799\
        );

    \I__9479\ : CascadeMux
    port map (
            O => \N__39837\,
            I => \N__39796\
        );

    \I__9478\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39792\
        );

    \I__9477\ : InMux
    port map (
            O => \N__39833\,
            I => \N__39789\
        );

    \I__9476\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39786\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__39829\,
            I => \N__39783\
        );

    \I__9474\ : InMux
    port map (
            O => \N__39826\,
            I => \N__39780\
        );

    \I__9473\ : InMux
    port map (
            O => \N__39825\,
            I => \N__39777\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__39822\,
            I => \N__39774\
        );

    \I__9471\ : InMux
    port map (
            O => \N__39821\,
            I => \N__39771\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__39818\,
            I => \N__39768\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39765\
        );

    \I__9468\ : InMux
    port map (
            O => \N__39814\,
            I => \N__39762\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__39809\,
            I => \N__39759\
        );

    \I__9466\ : InMux
    port map (
            O => \N__39808\,
            I => \N__39756\
        );

    \I__9465\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39753\
        );

    \I__9464\ : Span4Mux_h
    port map (
            O => \N__39804\,
            I => \N__39748\
        );

    \I__9463\ : Span4Mux_h
    port map (
            O => \N__39799\,
            I => \N__39745\
        );

    \I__9462\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39740\
        );

    \I__9461\ : InMux
    port map (
            O => \N__39795\,
            I => \N__39740\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__39792\,
            I => \N__39737\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__39789\,
            I => \N__39734\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__39786\,
            I => \N__39731\
        );

    \I__9457\ : Span4Mux_v
    port map (
            O => \N__39783\,
            I => \N__39728\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__39780\,
            I => \N__39725\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__39777\,
            I => \N__39722\
        );

    \I__9454\ : Span4Mux_v
    port map (
            O => \N__39774\,
            I => \N__39717\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__39771\,
            I => \N__39717\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__39768\,
            I => \N__39712\
        );

    \I__9451\ : Span4Mux_v
    port map (
            O => \N__39765\,
            I => \N__39712\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__39762\,
            I => \N__39709\
        );

    \I__9449\ : Span4Mux_v
    port map (
            O => \N__39759\,
            I => \N__39704\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__39756\,
            I => \N__39704\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__39753\,
            I => \N__39701\
        );

    \I__9446\ : InMux
    port map (
            O => \N__39752\,
            I => \N__39698\
        );

    \I__9445\ : InMux
    port map (
            O => \N__39751\,
            I => \N__39695\
        );

    \I__9444\ : Span4Mux_h
    port map (
            O => \N__39748\,
            I => \N__39692\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__39745\,
            I => \N__39689\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__39740\,
            I => \N__39686\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__39737\,
            I => \N__39681\
        );

    \I__9440\ : Span4Mux_h
    port map (
            O => \N__39734\,
            I => \N__39681\
        );

    \I__9439\ : Span4Mux_v
    port map (
            O => \N__39731\,
            I => \N__39676\
        );

    \I__9438\ : Span4Mux_h
    port map (
            O => \N__39728\,
            I => \N__39676\
        );

    \I__9437\ : Span4Mux_v
    port map (
            O => \N__39725\,
            I => \N__39665\
        );

    \I__9436\ : Span4Mux_v
    port map (
            O => \N__39722\,
            I => \N__39665\
        );

    \I__9435\ : Span4Mux_v
    port map (
            O => \N__39717\,
            I => \N__39665\
        );

    \I__9434\ : Span4Mux_h
    port map (
            O => \N__39712\,
            I => \N__39665\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__39709\,
            I => \N__39665\
        );

    \I__9432\ : Span4Mux_v
    port map (
            O => \N__39704\,
            I => \N__39656\
        );

    \I__9431\ : Span4Mux_s3_h
    port map (
            O => \N__39701\,
            I => \N__39656\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39656\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__39695\,
            I => \N__39656\
        );

    \I__9428\ : Odrv4
    port map (
            O => \N__39692\,
            I => \ALU.aluOut_9\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__39689\,
            I => \ALU.aluOut_9\
        );

    \I__9426\ : Odrv12
    port map (
            O => \N__39686\,
            I => \ALU.aluOut_9\
        );

    \I__9425\ : Odrv4
    port map (
            O => \N__39681\,
            I => \ALU.aluOut_9\
        );

    \I__9424\ : Odrv4
    port map (
            O => \N__39676\,
            I => \ALU.aluOut_9\
        );

    \I__9423\ : Odrv4
    port map (
            O => \N__39665\,
            I => \ALU.aluOut_9\
        );

    \I__9422\ : Odrv4
    port map (
            O => \N__39656\,
            I => \ALU.aluOut_9\
        );

    \I__9421\ : CascadeMux
    port map (
            O => \N__39641\,
            I => \N__39638\
        );

    \I__9420\ : InMux
    port map (
            O => \N__39638\,
            I => \N__39635\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__39635\,
            I => \N__39632\
        );

    \I__9418\ : Span4Mux_v
    port map (
            O => \N__39632\,
            I => \N__39629\
        );

    \I__9417\ : Sp12to4
    port map (
            O => \N__39629\,
            I => \N__39626\
        );

    \I__9416\ : Odrv12
    port map (
            O => \N__39626\,
            I => \ALU.N_207_0_i\
        );

    \I__9415\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39620\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__39620\,
            I => \N__39617\
        );

    \I__9413\ : Span4Mux_v
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__39614\,
            I => \ALU.un9_addsub_cry_8_c_RNIPV1SZ0Z8\
        );

    \I__9411\ : InMux
    port map (
            O => \N__39611\,
            I => \ALU.un9_addsub_cry_8\
        );

    \I__9410\ : CascadeMux
    port map (
            O => \N__39608\,
            I => \N__39602\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__39607\,
            I => \N__39596\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__39606\,
            I => \N__39590\
        );

    \I__9407\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39587\
        );

    \I__9406\ : InMux
    port map (
            O => \N__39602\,
            I => \N__39579\
        );

    \I__9405\ : InMux
    port map (
            O => \N__39601\,
            I => \N__39579\
        );

    \I__9404\ : InMux
    port map (
            O => \N__39600\,
            I => \N__39579\
        );

    \I__9403\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39572\
        );

    \I__9402\ : InMux
    port map (
            O => \N__39596\,
            I => \N__39572\
        );

    \I__9401\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39572\
        );

    \I__9400\ : InMux
    port map (
            O => \N__39594\,
            I => \N__39566\
        );

    \I__9399\ : InMux
    port map (
            O => \N__39593\,
            I => \N__39566\
        );

    \I__9398\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39563\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__39587\,
            I => \N__39560\
        );

    \I__9396\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39557\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__39579\,
            I => \N__39554\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__39572\,
            I => \N__39551\
        );

    \I__9393\ : InMux
    port map (
            O => \N__39571\,
            I => \N__39548\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__39566\,
            I => \N__39545\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__39563\,
            I => \N__39540\
        );

    \I__9390\ : Span4Mux_h
    port map (
            O => \N__39560\,
            I => \N__39540\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__39557\,
            I => \N__39537\
        );

    \I__9388\ : Span4Mux_v
    port map (
            O => \N__39554\,
            I => \N__39532\
        );

    \I__9387\ : Span4Mux_s1_h
    port map (
            O => \N__39551\,
            I => \N__39532\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__39548\,
            I => \N__39528\
        );

    \I__9385\ : Span4Mux_h
    port map (
            O => \N__39545\,
            I => \N__39525\
        );

    \I__9384\ : Span4Mux_h
    port map (
            O => \N__39540\,
            I => \N__39518\
        );

    \I__9383\ : Span4Mux_v
    port map (
            O => \N__39537\,
            I => \N__39518\
        );

    \I__9382\ : Span4Mux_h
    port map (
            O => \N__39532\,
            I => \N__39518\
        );

    \I__9381\ : InMux
    port map (
            O => \N__39531\,
            I => \N__39515\
        );

    \I__9380\ : Odrv12
    port map (
            O => \N__39528\,
            I => \ALU.N_192_0\
        );

    \I__9379\ : Odrv4
    port map (
            O => \N__39525\,
            I => \ALU.N_192_0\
        );

    \I__9378\ : Odrv4
    port map (
            O => \N__39518\,
            I => \ALU.N_192_0\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__39515\,
            I => \ALU.N_192_0\
        );

    \I__9376\ : CascadeMux
    port map (
            O => \N__39506\,
            I => \N__39503\
        );

    \I__9375\ : InMux
    port map (
            O => \N__39503\,
            I => \N__39500\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__39500\,
            I => \N__39497\
        );

    \I__9373\ : Sp12to4
    port map (
            O => \N__39497\,
            I => \N__39494\
        );

    \I__9372\ : Span12Mux_h
    port map (
            O => \N__39494\,
            I => \N__39491\
        );

    \I__9371\ : Odrv12
    port map (
            O => \N__39491\,
            I => \ALU.a_RNIV2S0FZ0Z_10\
        );

    \I__9370\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39485\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__39485\,
            I => \N__39482\
        );

    \I__9368\ : Odrv12
    port map (
            O => \N__39482\,
            I => \ALU.un9_addsub_cry_9_c_RNI22U6KZ0\
        );

    \I__9367\ : InMux
    port map (
            O => \N__39479\,
            I => \ALU.un9_addsub_cry_9\
        );

    \I__9366\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39473\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__39473\,
            I => \N__39468\
        );

    \I__9364\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39464\
        );

    \I__9363\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39460\
        );

    \I__9362\ : Span4Mux_v
    port map (
            O => \N__39468\,
            I => \N__39457\
        );

    \I__9361\ : InMux
    port map (
            O => \N__39467\,
            I => \N__39454\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__39464\,
            I => \N__39449\
        );

    \I__9359\ : InMux
    port map (
            O => \N__39463\,
            I => \N__39444\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__39460\,
            I => \N__39441\
        );

    \I__9357\ : Sp12to4
    port map (
            O => \N__39457\,
            I => \N__39435\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__39454\,
            I => \N__39435\
        );

    \I__9355\ : InMux
    port map (
            O => \N__39453\,
            I => \N__39430\
        );

    \I__9354\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39430\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__39449\,
            I => \N__39427\
        );

    \I__9352\ : InMux
    port map (
            O => \N__39448\,
            I => \N__39422\
        );

    \I__9351\ : InMux
    port map (
            O => \N__39447\,
            I => \N__39422\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__39444\,
            I => \N__39419\
        );

    \I__9349\ : Span4Mux_v
    port map (
            O => \N__39441\,
            I => \N__39416\
        );

    \I__9348\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39413\
        );

    \I__9347\ : Odrv12
    port map (
            O => \N__39435\,
            I => \ALU.N_186_0\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__39430\,
            I => \ALU.N_186_0\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__39427\,
            I => \ALU.N_186_0\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__39422\,
            I => \ALU.N_186_0\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__39419\,
            I => \ALU.N_186_0\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__39416\,
            I => \ALU.N_186_0\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__39413\,
            I => \ALU.N_186_0\
        );

    \I__9340\ : CascadeMux
    port map (
            O => \N__39398\,
            I => \N__39391\
        );

    \I__9339\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39379\
        );

    \I__9338\ : CascadeMux
    port map (
            O => \N__39396\,
            I => \N__39376\
        );

    \I__9337\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39372\
        );

    \I__9336\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39369\
        );

    \I__9335\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39365\
        );

    \I__9334\ : InMux
    port map (
            O => \N__39390\,
            I => \N__39362\
        );

    \I__9333\ : InMux
    port map (
            O => \N__39389\,
            I => \N__39359\
        );

    \I__9332\ : InMux
    port map (
            O => \N__39388\,
            I => \N__39356\
        );

    \I__9331\ : InMux
    port map (
            O => \N__39387\,
            I => \N__39351\
        );

    \I__9330\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39351\
        );

    \I__9329\ : InMux
    port map (
            O => \N__39385\,
            I => \N__39348\
        );

    \I__9328\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39345\
        );

    \I__9327\ : CascadeMux
    port map (
            O => \N__39383\,
            I => \N__39342\
        );

    \I__9326\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39338\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__39379\,
            I => \N__39335\
        );

    \I__9324\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39331\
        );

    \I__9323\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39328\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39323\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__39369\,
            I => \N__39323\
        );

    \I__9320\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39319\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39316\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__39362\,
            I => \N__39313\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__39359\,
            I => \N__39308\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__39356\,
            I => \N__39308\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39301\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__39348\,
            I => \N__39301\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__39345\,
            I => \N__39301\
        );

    \I__9312\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39296\
        );

    \I__9311\ : InMux
    port map (
            O => \N__39341\,
            I => \N__39296\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__39338\,
            I => \N__39293\
        );

    \I__9309\ : Span4Mux_v
    port map (
            O => \N__39335\,
            I => \N__39290\
        );

    \I__9308\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39287\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__39331\,
            I => \N__39279\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__39328\,
            I => \N__39279\
        );

    \I__9305\ : Span4Mux_v
    port map (
            O => \N__39323\,
            I => \N__39279\
        );

    \I__9304\ : InMux
    port map (
            O => \N__39322\,
            I => \N__39276\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__39319\,
            I => \N__39273\
        );

    \I__9302\ : Span4Mux_v
    port map (
            O => \N__39316\,
            I => \N__39270\
        );

    \I__9301\ : Span4Mux_v
    port map (
            O => \N__39313\,
            I => \N__39267\
        );

    \I__9300\ : Span4Mux_h
    port map (
            O => \N__39308\,
            I => \N__39260\
        );

    \I__9299\ : Span4Mux_v
    port map (
            O => \N__39301\,
            I => \N__39260\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__39296\,
            I => \N__39260\
        );

    \I__9297\ : Span4Mux_v
    port map (
            O => \N__39293\,
            I => \N__39253\
        );

    \I__9296\ : Span4Mux_h
    port map (
            O => \N__39290\,
            I => \N__39253\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__39287\,
            I => \N__39253\
        );

    \I__9294\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39250\
        );

    \I__9293\ : Span4Mux_v
    port map (
            O => \N__39279\,
            I => \N__39247\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__39276\,
            I => \N__39244\
        );

    \I__9291\ : Span4Mux_v
    port map (
            O => \N__39273\,
            I => \N__39241\
        );

    \I__9290\ : Span4Mux_h
    port map (
            O => \N__39270\,
            I => \N__39232\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__39267\,
            I => \N__39232\
        );

    \I__9288\ : Span4Mux_v
    port map (
            O => \N__39260\,
            I => \N__39232\
        );

    \I__9287\ : Span4Mux_v
    port map (
            O => \N__39253\,
            I => \N__39232\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__39250\,
            I => \N__39229\
        );

    \I__9285\ : Span4Mux_s3_h
    port map (
            O => \N__39247\,
            I => \N__39224\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__39244\,
            I => \N__39224\
        );

    \I__9283\ : Sp12to4
    port map (
            O => \N__39241\,
            I => \N__39219\
        );

    \I__9282\ : Sp12to4
    port map (
            O => \N__39232\,
            I => \N__39219\
        );

    \I__9281\ : Odrv12
    port map (
            O => \N__39229\,
            I => \ALU.aluOut_11\
        );

    \I__9280\ : Odrv4
    port map (
            O => \N__39224\,
            I => \ALU.aluOut_11\
        );

    \I__9279\ : Odrv12
    port map (
            O => \N__39219\,
            I => \ALU.aluOut_11\
        );

    \I__9278\ : InMux
    port map (
            O => \N__39212\,
            I => \N__39209\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__39209\,
            I => \N__39206\
        );

    \I__9276\ : Odrv4
    port map (
            O => \N__39206\,
            I => \ALU.un9_addsub_cry_10_c_RNI9C0KZ0Z9\
        );

    \I__9275\ : InMux
    port map (
            O => \N__39203\,
            I => \ALU.un9_addsub_cry_10\
        );

    \I__9274\ : InMux
    port map (
            O => \N__39200\,
            I => \N__39196\
        );

    \I__9273\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39193\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__39196\,
            I => \N__39188\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__39193\,
            I => \N__39188\
        );

    \I__9270\ : Odrv12
    port map (
            O => \N__39188\,
            I => \ALU.N_361\
        );

    \I__9269\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39182\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__39182\,
            I => \N__39177\
        );

    \I__9267\ : InMux
    port map (
            O => \N__39181\,
            I => \N__39174\
        );

    \I__9266\ : InMux
    port map (
            O => \N__39180\,
            I => \N__39171\
        );

    \I__9265\ : Span4Mux_h
    port map (
            O => \N__39177\,
            I => \N__39168\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__39174\,
            I => \N__39165\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__39171\,
            I => \N__39162\
        );

    \I__9262\ : Span4Mux_h
    port map (
            O => \N__39168\,
            I => \N__39157\
        );

    \I__9261\ : Span4Mux_h
    port map (
            O => \N__39165\,
            I => \N__39157\
        );

    \I__9260\ : Odrv4
    port map (
            O => \N__39162\,
            I => \ALU.N_244\
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__39157\,
            I => \ALU.N_244\
        );

    \I__9258\ : InMux
    port map (
            O => \N__39152\,
            I => \N__39134\
        );

    \I__9257\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39134\
        );

    \I__9256\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39129\
        );

    \I__9255\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39129\
        );

    \I__9254\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39122\
        );

    \I__9253\ : InMux
    port map (
            O => \N__39147\,
            I => \N__39122\
        );

    \I__9252\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39122\
        );

    \I__9251\ : InMux
    port map (
            O => \N__39145\,
            I => \N__39117\
        );

    \I__9250\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39117\
        );

    \I__9249\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39112\
        );

    \I__9248\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39112\
        );

    \I__9247\ : InMux
    port map (
            O => \N__39141\,
            I => \N__39109\
        );

    \I__9246\ : CascadeMux
    port map (
            O => \N__39140\,
            I => \N__39106\
        );

    \I__9245\ : CascadeMux
    port map (
            O => \N__39139\,
            I => \N__39102\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__39134\,
            I => \N__39099\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__39129\,
            I => \N__39088\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__39122\,
            I => \N__39088\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__39117\,
            I => \N__39088\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__39112\,
            I => \N__39088\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__39109\,
            I => \N__39088\
        );

    \I__9238\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39085\
        );

    \I__9237\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39071\
        );

    \I__9236\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39071\
        );

    \I__9235\ : Span4Mux_v
    port map (
            O => \N__39099\,
            I => \N__39062\
        );

    \I__9234\ : Span4Mux_v
    port map (
            O => \N__39088\,
            I => \N__39062\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__39085\,
            I => \N__39062\
        );

    \I__9232\ : CascadeMux
    port map (
            O => \N__39084\,
            I => \N__39058\
        );

    \I__9231\ : CascadeMux
    port map (
            O => \N__39083\,
            I => \N__39055\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__39082\,
            I => \N__39050\
        );

    \I__9229\ : CascadeMux
    port map (
            O => \N__39081\,
            I => \N__39047\
        );

    \I__9228\ : CascadeMux
    port map (
            O => \N__39080\,
            I => \N__39041\
        );

    \I__9227\ : CascadeMux
    port map (
            O => \N__39079\,
            I => \N__39038\
        );

    \I__9226\ : CascadeMux
    port map (
            O => \N__39078\,
            I => \N__39033\
        );

    \I__9225\ : CascadeMux
    port map (
            O => \N__39077\,
            I => \N__39030\
        );

    \I__9224\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39026\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__39071\,
            I => \N__39023\
        );

    \I__9222\ : InMux
    port map (
            O => \N__39070\,
            I => \N__39019\
        );

    \I__9221\ : CascadeMux
    port map (
            O => \N__39069\,
            I => \N__39007\
        );

    \I__9220\ : Span4Mux_h
    port map (
            O => \N__39062\,
            I => \N__39002\
        );

    \I__9219\ : InMux
    port map (
            O => \N__39061\,
            I => \N__38995\
        );

    \I__9218\ : InMux
    port map (
            O => \N__39058\,
            I => \N__38995\
        );

    \I__9217\ : InMux
    port map (
            O => \N__39055\,
            I => \N__38995\
        );

    \I__9216\ : InMux
    port map (
            O => \N__39054\,
            I => \N__38986\
        );

    \I__9215\ : InMux
    port map (
            O => \N__39053\,
            I => \N__38986\
        );

    \I__9214\ : InMux
    port map (
            O => \N__39050\,
            I => \N__38986\
        );

    \I__9213\ : InMux
    port map (
            O => \N__39047\,
            I => \N__38986\
        );

    \I__9212\ : InMux
    port map (
            O => \N__39046\,
            I => \N__38975\
        );

    \I__9211\ : InMux
    port map (
            O => \N__39045\,
            I => \N__38975\
        );

    \I__9210\ : InMux
    port map (
            O => \N__39044\,
            I => \N__38975\
        );

    \I__9209\ : InMux
    port map (
            O => \N__39041\,
            I => \N__38975\
        );

    \I__9208\ : InMux
    port map (
            O => \N__39038\,
            I => \N__38975\
        );

    \I__9207\ : InMux
    port map (
            O => \N__39037\,
            I => \N__38962\
        );

    \I__9206\ : InMux
    port map (
            O => \N__39036\,
            I => \N__38955\
        );

    \I__9205\ : InMux
    port map (
            O => \N__39033\,
            I => \N__38955\
        );

    \I__9204\ : InMux
    port map (
            O => \N__39030\,
            I => \N__38955\
        );

    \I__9203\ : InMux
    port map (
            O => \N__39029\,
            I => \N__38952\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__39026\,
            I => \N__38949\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__39023\,
            I => \N__38946\
        );

    \I__9200\ : InMux
    port map (
            O => \N__39022\,
            I => \N__38943\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__39019\,
            I => \N__38940\
        );

    \I__9198\ : InMux
    port map (
            O => \N__39018\,
            I => \N__38933\
        );

    \I__9197\ : InMux
    port map (
            O => \N__39017\,
            I => \N__38933\
        );

    \I__9196\ : InMux
    port map (
            O => \N__39016\,
            I => \N__38933\
        );

    \I__9195\ : InMux
    port map (
            O => \N__39015\,
            I => \N__38930\
        );

    \I__9194\ : InMux
    port map (
            O => \N__39014\,
            I => \N__38927\
        );

    \I__9193\ : InMux
    port map (
            O => \N__39013\,
            I => \N__38924\
        );

    \I__9192\ : InMux
    port map (
            O => \N__39012\,
            I => \N__38919\
        );

    \I__9191\ : InMux
    port map (
            O => \N__39011\,
            I => \N__38912\
        );

    \I__9190\ : InMux
    port map (
            O => \N__39010\,
            I => \N__38912\
        );

    \I__9189\ : InMux
    port map (
            O => \N__39007\,
            I => \N__38912\
        );

    \I__9188\ : InMux
    port map (
            O => \N__39006\,
            I => \N__38907\
        );

    \I__9187\ : InMux
    port map (
            O => \N__39005\,
            I => \N__38907\
        );

    \I__9186\ : Span4Mux_v
    port map (
            O => \N__39002\,
            I => \N__38902\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__38995\,
            I => \N__38902\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__38986\,
            I => \N__38897\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__38975\,
            I => \N__38897\
        );

    \I__9182\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38892\
        );

    \I__9181\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38892\
        );

    \I__9180\ : CascadeMux
    port map (
            O => \N__38972\,
            I => \N__38889\
        );

    \I__9179\ : CascadeMux
    port map (
            O => \N__38971\,
            I => \N__38884\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__38970\,
            I => \N__38881\
        );

    \I__9177\ : CascadeMux
    port map (
            O => \N__38969\,
            I => \N__38878\
        );

    \I__9176\ : CascadeMux
    port map (
            O => \N__38968\,
            I => \N__38875\
        );

    \I__9175\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38868\
        );

    \I__9174\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38868\
        );

    \I__9173\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38868\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__38962\,
            I => \N__38865\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__38955\,
            I => \N__38860\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__38952\,
            I => \N__38860\
        );

    \I__9169\ : Span4Mux_h
    port map (
            O => \N__38949\,
            I => \N__38855\
        );

    \I__9168\ : Span4Mux_v
    port map (
            O => \N__38946\,
            I => \N__38855\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__38943\,
            I => \N__38850\
        );

    \I__9166\ : Span4Mux_v
    port map (
            O => \N__38940\,
            I => \N__38850\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__38933\,
            I => \N__38847\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__38930\,
            I => \N__38840\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__38927\,
            I => \N__38840\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__38924\,
            I => \N__38840\
        );

    \I__9161\ : InMux
    port map (
            O => \N__38923\,
            I => \N__38835\
        );

    \I__9160\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38835\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__38919\,
            I => \N__38822\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__38912\,
            I => \N__38822\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__38907\,
            I => \N__38822\
        );

    \I__9156\ : Span4Mux_s2_v
    port map (
            O => \N__38902\,
            I => \N__38822\
        );

    \I__9155\ : Span4Mux_h
    port map (
            O => \N__38897\,
            I => \N__38822\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__38892\,
            I => \N__38822\
        );

    \I__9153\ : InMux
    port map (
            O => \N__38889\,
            I => \N__38819\
        );

    \I__9152\ : InMux
    port map (
            O => \N__38888\,
            I => \N__38814\
        );

    \I__9151\ : InMux
    port map (
            O => \N__38887\,
            I => \N__38814\
        );

    \I__9150\ : InMux
    port map (
            O => \N__38884\,
            I => \N__38807\
        );

    \I__9149\ : InMux
    port map (
            O => \N__38881\,
            I => \N__38807\
        );

    \I__9148\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38807\
        );

    \I__9147\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38804\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__38868\,
            I => \N__38801\
        );

    \I__9145\ : Span4Mux_v
    port map (
            O => \N__38865\,
            I => \N__38794\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__38860\,
            I => \N__38794\
        );

    \I__9143\ : Span4Mux_v
    port map (
            O => \N__38855\,
            I => \N__38794\
        );

    \I__9142\ : Span4Mux_h
    port map (
            O => \N__38850\,
            I => \N__38785\
        );

    \I__9141\ : Span4Mux_v
    port map (
            O => \N__38847\,
            I => \N__38785\
        );

    \I__9140\ : Span4Mux_v
    port map (
            O => \N__38840\,
            I => \N__38785\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__38835\,
            I => \N__38785\
        );

    \I__9138\ : Span4Mux_h
    port map (
            O => \N__38822\,
            I => \N__38782\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__38819\,
            I => \aluParams_1\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__38814\,
            I => \aluParams_1\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__38807\,
            I => \aluParams_1\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__38804\,
            I => \aluParams_1\
        );

    \I__9133\ : Odrv4
    port map (
            O => \N__38801\,
            I => \aluParams_1\
        );

    \I__9132\ : Odrv4
    port map (
            O => \N__38794\,
            I => \aluParams_1\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__38785\,
            I => \aluParams_1\
        );

    \I__9130\ : Odrv4
    port map (
            O => \N__38782\,
            I => \aluParams_1\
        );

    \I__9129\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38762\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__38762\,
            I => \N__38759\
        );

    \I__9127\ : Span4Mux_v
    port map (
            O => \N__38759\,
            I => \N__38756\
        );

    \I__9126\ : Span4Mux_h
    port map (
            O => \N__38756\,
            I => \N__38752\
        );

    \I__9125\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38749\
        );

    \I__9124\ : Odrv4
    port map (
            O => \N__38752\,
            I => \ALU.N_588\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__38749\,
            I => \ALU.N_588\
        );

    \I__9122\ : InMux
    port map (
            O => \N__38744\,
            I => \N__38740\
        );

    \I__9121\ : InMux
    port map (
            O => \N__38743\,
            I => \N__38736\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__38740\,
            I => \N__38719\
        );

    \I__9119\ : CascadeMux
    port map (
            O => \N__38739\,
            I => \N__38716\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__38736\,
            I => \N__38710\
        );

    \I__9117\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38707\
        );

    \I__9116\ : CascadeMux
    port map (
            O => \N__38734\,
            I => \N__38704\
        );

    \I__9115\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38701\
        );

    \I__9114\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38698\
        );

    \I__9113\ : InMux
    port map (
            O => \N__38731\,
            I => \N__38693\
        );

    \I__9112\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38690\
        );

    \I__9111\ : CascadeMux
    port map (
            O => \N__38729\,
            I => \N__38686\
        );

    \I__9110\ : InMux
    port map (
            O => \N__38728\,
            I => \N__38682\
        );

    \I__9109\ : CascadeMux
    port map (
            O => \N__38727\,
            I => \N__38679\
        );

    \I__9108\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38673\
        );

    \I__9107\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38668\
        );

    \I__9106\ : InMux
    port map (
            O => \N__38724\,
            I => \N__38668\
        );

    \I__9105\ : InMux
    port map (
            O => \N__38723\,
            I => \N__38663\
        );

    \I__9104\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38663\
        );

    \I__9103\ : Span4Mux_v
    port map (
            O => \N__38719\,
            I => \N__38660\
        );

    \I__9102\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38657\
        );

    \I__9101\ : CascadeMux
    port map (
            O => \N__38715\,
            I => \N__38654\
        );

    \I__9100\ : CascadeMux
    port map (
            O => \N__38714\,
            I => \N__38649\
        );

    \I__9099\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38643\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__38710\,
            I => \N__38640\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__38707\,
            I => \N__38637\
        );

    \I__9096\ : InMux
    port map (
            O => \N__38704\,
            I => \N__38634\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__38701\,
            I => \N__38631\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__38698\,
            I => \N__38628\
        );

    \I__9093\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38623\
        );

    \I__9092\ : InMux
    port map (
            O => \N__38696\,
            I => \N__38623\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__38693\,
            I => \N__38620\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__38690\,
            I => \N__38617\
        );

    \I__9089\ : InMux
    port map (
            O => \N__38689\,
            I => \N__38610\
        );

    \I__9088\ : InMux
    port map (
            O => \N__38686\,
            I => \N__38610\
        );

    \I__9087\ : InMux
    port map (
            O => \N__38685\,
            I => \N__38610\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__38682\,
            I => \N__38607\
        );

    \I__9085\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38604\
        );

    \I__9084\ : CascadeMux
    port map (
            O => \N__38678\,
            I => \N__38600\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__38677\,
            I => \N__38597\
        );

    \I__9082\ : CascadeMux
    port map (
            O => \N__38676\,
            I => \N__38594\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__38673\,
            I => \N__38584\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__38668\,
            I => \N__38584\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__38663\,
            I => \N__38584\
        );

    \I__9078\ : Sp12to4
    port map (
            O => \N__38660\,
            I => \N__38579\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__38657\,
            I => \N__38579\
        );

    \I__9076\ : InMux
    port map (
            O => \N__38654\,
            I => \N__38576\
        );

    \I__9075\ : InMux
    port map (
            O => \N__38653\,
            I => \N__38571\
        );

    \I__9074\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38571\
        );

    \I__9073\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38566\
        );

    \I__9072\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38566\
        );

    \I__9071\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38561\
        );

    \I__9070\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38561\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__38643\,
            I => \N__38556\
        );

    \I__9068\ : Span4Mux_v
    port map (
            O => \N__38640\,
            I => \N__38553\
        );

    \I__9067\ : Span4Mux_v
    port map (
            O => \N__38637\,
            I => \N__38548\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__38634\,
            I => \N__38548\
        );

    \I__9065\ : Span4Mux_s3_h
    port map (
            O => \N__38631\,
            I => \N__38541\
        );

    \I__9064\ : Span4Mux_v
    port map (
            O => \N__38628\,
            I => \N__38541\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__38623\,
            I => \N__38541\
        );

    \I__9062\ : Span4Mux_h
    port map (
            O => \N__38620\,
            I => \N__38529\
        );

    \I__9061\ : Span4Mux_h
    port map (
            O => \N__38617\,
            I => \N__38529\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__38610\,
            I => \N__38529\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__38607\,
            I => \N__38529\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__38604\,
            I => \N__38529\
        );

    \I__9057\ : CascadeMux
    port map (
            O => \N__38603\,
            I => \N__38525\
        );

    \I__9056\ : InMux
    port map (
            O => \N__38600\,
            I => \N__38522\
        );

    \I__9055\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38517\
        );

    \I__9054\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38517\
        );

    \I__9053\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38514\
        );

    \I__9052\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38509\
        );

    \I__9051\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38509\
        );

    \I__9050\ : Sp12to4
    port map (
            O => \N__38584\,
            I => \N__38504\
        );

    \I__9049\ : Span12Mux_h
    port map (
            O => \N__38579\,
            I => \N__38504\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__38576\,
            I => \N__38495\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38495\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__38566\,
            I => \N__38495\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__38561\,
            I => \N__38495\
        );

    \I__9044\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38490\
        );

    \I__9043\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38490\
        );

    \I__9042\ : Span4Mux_h
    port map (
            O => \N__38556\,
            I => \N__38485\
        );

    \I__9041\ : Span4Mux_v
    port map (
            O => \N__38553\,
            I => \N__38485\
        );

    \I__9040\ : Span4Mux_h
    port map (
            O => \N__38548\,
            I => \N__38480\
        );

    \I__9039\ : Span4Mux_h
    port map (
            O => \N__38541\,
            I => \N__38480\
        );

    \I__9038\ : InMux
    port map (
            O => \N__38540\,
            I => \N__38477\
        );

    \I__9037\ : Span4Mux_v
    port map (
            O => \N__38529\,
            I => \N__38474\
        );

    \I__9036\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38469\
        );

    \I__9035\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38469\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__38522\,
            I => \aluParams_2\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__38517\,
            I => \aluParams_2\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__38514\,
            I => \aluParams_2\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__38509\,
            I => \aluParams_2\
        );

    \I__9030\ : Odrv12
    port map (
            O => \N__38504\,
            I => \aluParams_2\
        );

    \I__9029\ : Odrv12
    port map (
            O => \N__38495\,
            I => \aluParams_2\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__38490\,
            I => \aluParams_2\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__38485\,
            I => \aluParams_2\
        );

    \I__9026\ : Odrv4
    port map (
            O => \N__38480\,
            I => \aluParams_2\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__38477\,
            I => \aluParams_2\
        );

    \I__9024\ : Odrv4
    port map (
            O => \N__38474\,
            I => \aluParams_2\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__38469\,
            I => \aluParams_2\
        );

    \I__9022\ : InMux
    port map (
            O => \N__38444\,
            I => \N__38441\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__38441\,
            I => \N__38438\
        );

    \I__9020\ : Span4Mux_v
    port map (
            O => \N__38438\,
            I => \N__38433\
        );

    \I__9019\ : InMux
    port map (
            O => \N__38437\,
            I => \N__38428\
        );

    \I__9018\ : InMux
    port map (
            O => \N__38436\,
            I => \N__38425\
        );

    \I__9017\ : Sp12to4
    port map (
            O => \N__38433\,
            I => \N__38422\
        );

    \I__9016\ : InMux
    port map (
            O => \N__38432\,
            I => \N__38417\
        );

    \I__9015\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38417\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__38428\,
            I => \N__38414\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__38425\,
            I => \ALU.N_590\
        );

    \I__9012\ : Odrv12
    port map (
            O => \N__38422\,
            I => \ALU.N_590\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__38417\,
            I => \ALU.N_590\
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__38414\,
            I => \ALU.N_590\
        );

    \I__9009\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38402\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__38402\,
            I => \N__38398\
        );

    \I__9007\ : CascadeMux
    port map (
            O => \N__38401\,
            I => \N__38395\
        );

    \I__9006\ : Span4Mux_v
    port map (
            O => \N__38398\,
            I => \N__38392\
        );

    \I__9005\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38388\
        );

    \I__9004\ : Span4Mux_h
    port map (
            O => \N__38392\,
            I => \N__38385\
        );

    \I__9003\ : InMux
    port map (
            O => \N__38391\,
            I => \N__38382\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__38388\,
            I => \ALU.eZ0Z_9\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__38385\,
            I => \ALU.eZ0Z_9\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__38382\,
            I => \ALU.eZ0Z_9\
        );

    \I__8999\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__38372\,
            I => \N__38368\
        );

    \I__8997\ : InMux
    port map (
            O => \N__38371\,
            I => \N__38365\
        );

    \I__8996\ : Span4Mux_v
    port map (
            O => \N__38368\,
            I => \N__38361\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__38365\,
            I => \N__38358\
        );

    \I__8994\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38355\
        );

    \I__8993\ : Span4Mux_h
    port map (
            O => \N__38361\,
            I => \N__38350\
        );

    \I__8992\ : Span4Mux_v
    port map (
            O => \N__38358\,
            I => \N__38350\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__38355\,
            I => \ALU.aZ0Z_9\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__38350\,
            I => \ALU.aZ0Z_9\
        );

    \I__8989\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38342\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__38342\,
            I => \ALU.e_RNIR49HZ0Z_9\
        );

    \I__8987\ : CascadeMux
    port map (
            O => \N__38339\,
            I => \N__38333\
        );

    \I__8986\ : InMux
    port map (
            O => \N__38338\,
            I => \N__38326\
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__38337\,
            I => \N__38319\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__38336\,
            I => \N__38312\
        );

    \I__8983\ : InMux
    port map (
            O => \N__38333\,
            I => \N__38303\
        );

    \I__8982\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38300\
        );

    \I__8981\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38292\
        );

    \I__8980\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38292\
        );

    \I__8979\ : InMux
    port map (
            O => \N__38329\,
            I => \N__38292\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__38326\,
            I => \N__38288\
        );

    \I__8977\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38285\
        );

    \I__8976\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38282\
        );

    \I__8975\ : InMux
    port map (
            O => \N__38323\,
            I => \N__38275\
        );

    \I__8974\ : InMux
    port map (
            O => \N__38322\,
            I => \N__38275\
        );

    \I__8973\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38275\
        );

    \I__8972\ : InMux
    port map (
            O => \N__38318\,
            I => \N__38269\
        );

    \I__8971\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38264\
        );

    \I__8970\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38264\
        );

    \I__8969\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38257\
        );

    \I__8968\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38257\
        );

    \I__8967\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38257\
        );

    \I__8966\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38250\
        );

    \I__8965\ : InMux
    port map (
            O => \N__38309\,
            I => \N__38250\
        );

    \I__8964\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38250\
        );

    \I__8963\ : InMux
    port map (
            O => \N__38307\,
            I => \N__38242\
        );

    \I__8962\ : InMux
    port map (
            O => \N__38306\,
            I => \N__38242\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__38303\,
            I => \N__38239\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__38300\,
            I => \N__38236\
        );

    \I__8959\ : InMux
    port map (
            O => \N__38299\,
            I => \N__38233\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38230\
        );

    \I__8957\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38227\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__38288\,
            I => \N__38222\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38219\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__38282\,
            I => \N__38214\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__38275\,
            I => \N__38214\
        );

    \I__8952\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38210\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__38273\,
            I => \N__38207\
        );

    \I__8950\ : InMux
    port map (
            O => \N__38272\,
            I => \N__38204\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__38269\,
            I => \N__38199\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__38264\,
            I => \N__38199\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38196\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__38250\,
            I => \N__38193\
        );

    \I__8945\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38183\
        );

    \I__8944\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38183\
        );

    \I__8943\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38183\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38180\
        );

    \I__8941\ : Span4Mux_v
    port map (
            O => \N__38239\,
            I => \N__38173\
        );

    \I__8940\ : Span4Mux_v
    port map (
            O => \N__38236\,
            I => \N__38170\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38163\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__38230\,
            I => \N__38163\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38163\
        );

    \I__8936\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38158\
        );

    \I__8935\ : InMux
    port map (
            O => \N__38225\,
            I => \N__38158\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__38222\,
            I => \N__38153\
        );

    \I__8933\ : Span4Mux_h
    port map (
            O => \N__38219\,
            I => \N__38153\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__38214\,
            I => \N__38150\
        );

    \I__8931\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38147\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__38210\,
            I => \N__38144\
        );

    \I__8929\ : InMux
    port map (
            O => \N__38207\,
            I => \N__38141\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__38204\,
            I => \N__38138\
        );

    \I__8927\ : Span4Mux_v
    port map (
            O => \N__38199\,
            I => \N__38131\
        );

    \I__8926\ : Span4Mux_v
    port map (
            O => \N__38196\,
            I => \N__38131\
        );

    \I__8925\ : Span4Mux_s1_h
    port map (
            O => \N__38193\,
            I => \N__38131\
        );

    \I__8924\ : InMux
    port map (
            O => \N__38192\,
            I => \N__38126\
        );

    \I__8923\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38126\
        );

    \I__8922\ : InMux
    port map (
            O => \N__38190\,
            I => \N__38123\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__38183\,
            I => \N__38120\
        );

    \I__8920\ : Span12Mux_s4_v
    port map (
            O => \N__38180\,
            I => \N__38117\
        );

    \I__8919\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38114\
        );

    \I__8918\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38111\
        );

    \I__8917\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38108\
        );

    \I__8916\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38105\
        );

    \I__8915\ : Span4Mux_s2_h
    port map (
            O => \N__38173\,
            I => \N__38100\
        );

    \I__8914\ : Span4Mux_v
    port map (
            O => \N__38170\,
            I => \N__38100\
        );

    \I__8913\ : Span4Mux_v
    port map (
            O => \N__38163\,
            I => \N__38095\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__38158\,
            I => \N__38095\
        );

    \I__8911\ : Span4Mux_h
    port map (
            O => \N__38153\,
            I => \N__38092\
        );

    \I__8910\ : Span4Mux_v
    port map (
            O => \N__38150\,
            I => \N__38085\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__38147\,
            I => \N__38085\
        );

    \I__8908\ : Span4Mux_v
    port map (
            O => \N__38144\,
            I => \N__38085\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__38141\,
            I => \N__38076\
        );

    \I__8906\ : Span4Mux_h
    port map (
            O => \N__38138\,
            I => \N__38076\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__38131\,
            I => \N__38076\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__38126\,
            I => \N__38076\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__38123\,
            I => \ALU.N_252_0\
        );

    \I__8902\ : Odrv12
    port map (
            O => \N__38120\,
            I => \ALU.N_252_0\
        );

    \I__8901\ : Odrv12
    port map (
            O => \N__38117\,
            I => \ALU.N_252_0\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__38114\,
            I => \ALU.N_252_0\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__38111\,
            I => \ALU.N_252_0\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__38108\,
            I => \ALU.N_252_0\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__38105\,
            I => \ALU.N_252_0\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__38100\,
            I => \ALU.N_252_0\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__38095\,
            I => \ALU.N_252_0\
        );

    \I__8894\ : Odrv4
    port map (
            O => \N__38092\,
            I => \ALU.N_252_0\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__38085\,
            I => \ALU.N_252_0\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__38076\,
            I => \ALU.N_252_0\
        );

    \I__8891\ : CascadeMux
    port map (
            O => \N__38051\,
            I => \N__38048\
        );

    \I__8890\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38042\
        );

    \I__8889\ : CascadeMux
    port map (
            O => \N__38047\,
            I => \N__38038\
        );

    \I__8888\ : CascadeMux
    port map (
            O => \N__38046\,
            I => \N__38030\
        );

    \I__8887\ : CascadeMux
    port map (
            O => \N__38045\,
            I => \N__38019\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__38042\,
            I => \N__38016\
        );

    \I__8885\ : InMux
    port map (
            O => \N__38041\,
            I => \N__38013\
        );

    \I__8884\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38006\
        );

    \I__8883\ : InMux
    port map (
            O => \N__38037\,
            I => \N__38006\
        );

    \I__8882\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38006\
        );

    \I__8881\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38003\
        );

    \I__8880\ : InMux
    port map (
            O => \N__38034\,
            I => \N__37998\
        );

    \I__8879\ : InMux
    port map (
            O => \N__38033\,
            I => \N__37987\
        );

    \I__8878\ : InMux
    port map (
            O => \N__38030\,
            I => \N__37987\
        );

    \I__8877\ : InMux
    port map (
            O => \N__38029\,
            I => \N__37987\
        );

    \I__8876\ : InMux
    port map (
            O => \N__38028\,
            I => \N__37982\
        );

    \I__8875\ : InMux
    port map (
            O => \N__38027\,
            I => \N__37976\
        );

    \I__8874\ : InMux
    port map (
            O => \N__38026\,
            I => \N__37976\
        );

    \I__8873\ : InMux
    port map (
            O => \N__38025\,
            I => \N__37969\
        );

    \I__8872\ : InMux
    port map (
            O => \N__38024\,
            I => \N__37969\
        );

    \I__8871\ : InMux
    port map (
            O => \N__38023\,
            I => \N__37969\
        );

    \I__8870\ : InMux
    port map (
            O => \N__38022\,
            I => \N__37963\
        );

    \I__8869\ : InMux
    port map (
            O => \N__38019\,
            I => \N__37963\
        );

    \I__8868\ : Span4Mux_h
    port map (
            O => \N__38016\,
            I => \N__37956\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__37956\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__38006\,
            I => \N__37953\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__38003\,
            I => \N__37950\
        );

    \I__8864\ : InMux
    port map (
            O => \N__38002\,
            I => \N__37947\
        );

    \I__8863\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37944\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__37998\,
            I => \N__37941\
        );

    \I__8861\ : InMux
    port map (
            O => \N__37997\,
            I => \N__37938\
        );

    \I__8860\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37926\
        );

    \I__8859\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37926\
        );

    \I__8858\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37926\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__37987\,
            I => \N__37923\
        );

    \I__8856\ : InMux
    port map (
            O => \N__37986\,
            I => \N__37918\
        );

    \I__8855\ : InMux
    port map (
            O => \N__37985\,
            I => \N__37918\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__37982\,
            I => \N__37915\
        );

    \I__8853\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37912\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__37976\,
            I => \N__37907\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37907\
        );

    \I__8850\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37904\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37901\
        );

    \I__8848\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37898\
        );

    \I__8847\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37895\
        );

    \I__8846\ : Span4Mux_v
    port map (
            O => \N__37956\,
            I => \N__37891\
        );

    \I__8845\ : Span4Mux_v
    port map (
            O => \N__37953\,
            I => \N__37888\
        );

    \I__8844\ : Span4Mux_v
    port map (
            O => \N__37950\,
            I => \N__37883\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__37947\,
            I => \N__37883\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__37944\,
            I => \N__37876\
        );

    \I__8841\ : Span4Mux_h
    port map (
            O => \N__37941\,
            I => \N__37876\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37876\
        );

    \I__8839\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37867\
        );

    \I__8838\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37867\
        );

    \I__8837\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37867\
        );

    \I__8836\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37867\
        );

    \I__8835\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37864\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__37926\,
            I => \N__37861\
        );

    \I__8833\ : Span4Mux_v
    port map (
            O => \N__37923\,
            I => \N__37856\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__37918\,
            I => \N__37856\
        );

    \I__8831\ : Span4Mux_v
    port map (
            O => \N__37915\,
            I => \N__37847\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__37912\,
            I => \N__37847\
        );

    \I__8829\ : Span4Mux_h
    port map (
            O => \N__37907\,
            I => \N__37847\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__37904\,
            I => \N__37847\
        );

    \I__8827\ : Span12Mux_s3_v
    port map (
            O => \N__37901\,
            I => \N__37840\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__37898\,
            I => \N__37840\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__37895\,
            I => \N__37840\
        );

    \I__8824\ : InMux
    port map (
            O => \N__37894\,
            I => \N__37837\
        );

    \I__8823\ : Span4Mux_h
    port map (
            O => \N__37891\,
            I => \N__37834\
        );

    \I__8822\ : Span4Mux_h
    port map (
            O => \N__37888\,
            I => \N__37827\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__37883\,
            I => \N__37827\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__37876\,
            I => \N__37827\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__37867\,
            I => \N__37824\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__37864\,
            I => \N__37819\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__37861\,
            I => \N__37819\
        );

    \I__8816\ : Span4Mux_v
    port map (
            O => \N__37856\,
            I => \N__37816\
        );

    \I__8815\ : Span4Mux_v
    port map (
            O => \N__37847\,
            I => \N__37813\
        );

    \I__8814\ : Odrv12
    port map (
            O => \N__37840\,
            I => \ALU.aluOut_0\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__37837\,
            I => \ALU.aluOut_0\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__37834\,
            I => \ALU.aluOut_0\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__37827\,
            I => \ALU.aluOut_0\
        );

    \I__8810\ : Odrv12
    port map (
            O => \N__37824\,
            I => \ALU.aluOut_0\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__37819\,
            I => \ALU.aluOut_0\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__37816\,
            I => \ALU.aluOut_0\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__37813\,
            I => \ALU.aluOut_0\
        );

    \I__8806\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37793\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__37793\,
            I => \N__37790\
        );

    \I__8804\ : Odrv4
    port map (
            O => \N__37790\,
            I => \ALU.a0_b_2\
        );

    \I__8803\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37783\
        );

    \I__8802\ : CascadeMux
    port map (
            O => \N__37786\,
            I => \N__37780\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__37783\,
            I => \N__37777\
        );

    \I__8800\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37774\
        );

    \I__8799\ : Span4Mux_v
    port map (
            O => \N__37777\,
            I => \N__37770\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__37774\,
            I => \N__37764\
        );

    \I__8797\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37754\
        );

    \I__8796\ : Span4Mux_h
    port map (
            O => \N__37770\,
            I => \N__37751\
        );

    \I__8795\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37746\
        );

    \I__8794\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37746\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__37767\,
            I => \N__37743\
        );

    \I__8792\ : Span4Mux_h
    port map (
            O => \N__37764\,
            I => \N__37738\
        );

    \I__8791\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37733\
        );

    \I__8790\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37733\
        );

    \I__8789\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37725\
        );

    \I__8788\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37725\
        );

    \I__8787\ : InMux
    port map (
            O => \N__37759\,
            I => \N__37722\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__37758\,
            I => \N__37719\
        );

    \I__8785\ : InMux
    port map (
            O => \N__37757\,
            I => \N__37712\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__37754\,
            I => \N__37709\
        );

    \I__8783\ : Span4Mux_h
    port map (
            O => \N__37751\,
            I => \N__37704\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__37746\,
            I => \N__37704\
        );

    \I__8781\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37699\
        );

    \I__8780\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37696\
        );

    \I__8779\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37693\
        );

    \I__8778\ : Span4Mux_v
    port map (
            O => \N__37738\,
            I => \N__37688\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__37733\,
            I => \N__37688\
        );

    \I__8776\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37683\
        );

    \I__8775\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37683\
        );

    \I__8774\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37680\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N__37675\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__37722\,
            I => \N__37675\
        );

    \I__8771\ : InMux
    port map (
            O => \N__37719\,
            I => \N__37672\
        );

    \I__8770\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37669\
        );

    \I__8769\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37664\
        );

    \I__8768\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37664\
        );

    \I__8767\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37661\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__37712\,
            I => \N__37648\
        );

    \I__8765\ : Span4Mux_h
    port map (
            O => \N__37709\,
            I => \N__37641\
        );

    \I__8764\ : Span4Mux_v
    port map (
            O => \N__37704\,
            I => \N__37641\
        );

    \I__8763\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37636\
        );

    \I__8762\ : InMux
    port map (
            O => \N__37702\,
            I => \N__37636\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37633\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__37696\,
            I => \N__37628\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__37693\,
            I => \N__37628\
        );

    \I__8758\ : Span4Mux_h
    port map (
            O => \N__37688\,
            I => \N__37623\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__37683\,
            I => \N__37620\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__37680\,
            I => \N__37617\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__37675\,
            I => \N__37614\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__37672\,
            I => \N__37611\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__37669\,
            I => \N__37608\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37603\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__37661\,
            I => \N__37603\
        );

    \I__8750\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37596\
        );

    \I__8749\ : InMux
    port map (
            O => \N__37659\,
            I => \N__37596\
        );

    \I__8748\ : InMux
    port map (
            O => \N__37658\,
            I => \N__37596\
        );

    \I__8747\ : InMux
    port map (
            O => \N__37657\,
            I => \N__37593\
        );

    \I__8746\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37586\
        );

    \I__8745\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37586\
        );

    \I__8744\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37586\
        );

    \I__8743\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37583\
        );

    \I__8742\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37578\
        );

    \I__8741\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37578\
        );

    \I__8740\ : Span4Mux_h
    port map (
            O => \N__37648\,
            I => \N__37575\
        );

    \I__8739\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37570\
        );

    \I__8738\ : InMux
    port map (
            O => \N__37646\,
            I => \N__37570\
        );

    \I__8737\ : Span4Mux_v
    port map (
            O => \N__37641\,
            I => \N__37567\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__37636\,
            I => \N__37560\
        );

    \I__8735\ : Span4Mux_v
    port map (
            O => \N__37633\,
            I => \N__37560\
        );

    \I__8734\ : Span4Mux_v
    port map (
            O => \N__37628\,
            I => \N__37560\
        );

    \I__8733\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37555\
        );

    \I__8732\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37555\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__37623\,
            I => \N__37538\
        );

    \I__8730\ : Span4Mux_s3_h
    port map (
            O => \N__37620\,
            I => \N__37538\
        );

    \I__8729\ : Span4Mux_v
    port map (
            O => \N__37617\,
            I => \N__37538\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__37614\,
            I => \N__37538\
        );

    \I__8727\ : Span4Mux_s3_h
    port map (
            O => \N__37611\,
            I => \N__37538\
        );

    \I__8726\ : Span4Mux_v
    port map (
            O => \N__37608\,
            I => \N__37538\
        );

    \I__8725\ : Span4Mux_v
    port map (
            O => \N__37603\,
            I => \N__37538\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37538\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__37593\,
            I => \N__37533\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__37586\,
            I => \N__37533\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__37583\,
            I => \ALU.N_249_0_i\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__37578\,
            I => \ALU.N_249_0_i\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__37575\,
            I => \ALU.N_249_0_i\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__37570\,
            I => \ALU.N_249_0_i\
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__37567\,
            I => \ALU.N_249_0_i\
        );

    \I__8716\ : Odrv4
    port map (
            O => \N__37560\,
            I => \ALU.N_249_0_i\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__37555\,
            I => \ALU.N_249_0_i\
        );

    \I__8714\ : Odrv4
    port map (
            O => \N__37538\,
            I => \ALU.N_249_0_i\
        );

    \I__8713\ : Odrv12
    port map (
            O => \N__37533\,
            I => \ALU.N_249_0_i\
        );

    \I__8712\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37510\
        );

    \I__8711\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37507\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__37510\,
            I => \N__37504\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__37507\,
            I => \N__37497\
        );

    \I__8708\ : Span4Mux_v
    port map (
            O => \N__37504\,
            I => \N__37494\
        );

    \I__8707\ : InMux
    port map (
            O => \N__37503\,
            I => \N__37491\
        );

    \I__8706\ : CascadeMux
    port map (
            O => \N__37502\,
            I => \N__37481\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__37501\,
            I => \N__37476\
        );

    \I__8704\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37473\
        );

    \I__8703\ : Span4Mux_v
    port map (
            O => \N__37497\,
            I => \N__37468\
        );

    \I__8702\ : Span4Mux_s2_h
    port map (
            O => \N__37494\,
            I => \N__37463\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__37491\,
            I => \N__37463\
        );

    \I__8700\ : InMux
    port map (
            O => \N__37490\,
            I => \N__37456\
        );

    \I__8699\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37456\
        );

    \I__8698\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37456\
        );

    \I__8697\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37451\
        );

    \I__8696\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37451\
        );

    \I__8695\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37448\
        );

    \I__8694\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37444\
        );

    \I__8693\ : InMux
    port map (
            O => \N__37481\,
            I => \N__37439\
        );

    \I__8692\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37439\
        );

    \I__8691\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37436\
        );

    \I__8690\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37433\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37430\
        );

    \I__8688\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37420\
        );

    \I__8687\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37420\
        );

    \I__8686\ : Span4Mux_s2_h
    port map (
            O => \N__37468\,
            I => \N__37406\
        );

    \I__8685\ : Span4Mux_v
    port map (
            O => \N__37463\,
            I => \N__37406\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37406\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__37451\,
            I => \N__37406\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__37448\,
            I => \N__37406\
        );

    \I__8681\ : InMux
    port map (
            O => \N__37447\,
            I => \N__37403\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__37444\,
            I => \N__37400\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__37439\,
            I => \N__37397\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37392\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__37433\,
            I => \N__37392\
        );

    \I__8676\ : Span4Mux_v
    port map (
            O => \N__37430\,
            I => \N__37388\
        );

    \I__8675\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37383\
        );

    \I__8674\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37383\
        );

    \I__8673\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37380\
        );

    \I__8672\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37377\
        );

    \I__8671\ : CascadeMux
    port map (
            O => \N__37425\,
            I => \N__37373\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__37420\,
            I => \N__37368\
        );

    \I__8669\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37365\
        );

    \I__8668\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37362\
        );

    \I__8667\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37359\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__37406\,
            I => \N__37356\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__37403\,
            I => \N__37353\
        );

    \I__8664\ : Span4Mux_s2_h
    port map (
            O => \N__37400\,
            I => \N__37350\
        );

    \I__8663\ : Span4Mux_v
    port map (
            O => \N__37397\,
            I => \N__37342\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__37392\,
            I => \N__37342\
        );

    \I__8661\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37339\
        );

    \I__8660\ : Span4Mux_v
    port map (
            O => \N__37388\,
            I => \N__37334\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__37383\,
            I => \N__37334\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__37380\,
            I => \N__37329\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37329\
        );

    \I__8656\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37326\
        );

    \I__8655\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37319\
        );

    \I__8654\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37319\
        );

    \I__8653\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37319\
        );

    \I__8652\ : Span4Mux_h
    port map (
            O => \N__37368\,
            I => \N__37313\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__37365\,
            I => \N__37313\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__37362\,
            I => \N__37302\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__37359\,
            I => \N__37302\
        );

    \I__8648\ : Span4Mux_s2_h
    port map (
            O => \N__37356\,
            I => \N__37302\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__37353\,
            I => \N__37302\
        );

    \I__8646\ : Span4Mux_v
    port map (
            O => \N__37350\,
            I => \N__37302\
        );

    \I__8645\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37295\
        );

    \I__8644\ : InMux
    port map (
            O => \N__37348\,
            I => \N__37295\
        );

    \I__8643\ : InMux
    port map (
            O => \N__37347\,
            I => \N__37295\
        );

    \I__8642\ : Span4Mux_h
    port map (
            O => \N__37342\,
            I => \N__37290\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__37339\,
            I => \N__37290\
        );

    \I__8640\ : Span4Mux_h
    port map (
            O => \N__37334\,
            I => \N__37287\
        );

    \I__8639\ : Span4Mux_v
    port map (
            O => \N__37329\,
            I => \N__37280\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__37326\,
            I => \N__37280\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37280\
        );

    \I__8636\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37277\
        );

    \I__8635\ : Span4Mux_v
    port map (
            O => \N__37313\,
            I => \N__37272\
        );

    \I__8634\ : Span4Mux_h
    port map (
            O => \N__37302\,
            I => \N__37272\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__37295\,
            I => \ALU.aluOut_1\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__37290\,
            I => \ALU.aluOut_1\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__37287\,
            I => \ALU.aluOut_1\
        );

    \I__8630\ : Odrv4
    port map (
            O => \N__37280\,
            I => \ALU.aluOut_1\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__37277\,
            I => \ALU.aluOut_1\
        );

    \I__8628\ : Odrv4
    port map (
            O => \N__37272\,
            I => \ALU.aluOut_1\
        );

    \I__8627\ : InMux
    port map (
            O => \N__37259\,
            I => \ALU.un9_addsub_cry_0\
        );

    \I__8626\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37251\
        );

    \I__8625\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37246\
        );

    \I__8624\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37246\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37241\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__37246\,
            I => \N__37238\
        );

    \I__8621\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37228\
        );

    \I__8620\ : InMux
    port map (
            O => \N__37244\,
            I => \N__37225\
        );

    \I__8619\ : Span4Mux_v
    port map (
            O => \N__37241\,
            I => \N__37222\
        );

    \I__8618\ : Span4Mux_v
    port map (
            O => \N__37238\,
            I => \N__37219\
        );

    \I__8617\ : CascadeMux
    port map (
            O => \N__37237\,
            I => \N__37215\
        );

    \I__8616\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37211\
        );

    \I__8615\ : InMux
    port map (
            O => \N__37235\,
            I => \N__37206\
        );

    \I__8614\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37206\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__37233\,
            I => \N__37196\
        );

    \I__8612\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37191\
        );

    \I__8611\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37188\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37183\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__37225\,
            I => \N__37183\
        );

    \I__8608\ : Span4Mux_v
    port map (
            O => \N__37222\,
            I => \N__37180\
        );

    \I__8607\ : Span4Mux_v
    port map (
            O => \N__37219\,
            I => \N__37177\
        );

    \I__8606\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37174\
        );

    \I__8605\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37169\
        );

    \I__8604\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37169\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__37211\,
            I => \N__37164\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__37206\,
            I => \N__37164\
        );

    \I__8601\ : InMux
    port map (
            O => \N__37205\,
            I => \N__37159\
        );

    \I__8600\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37159\
        );

    \I__8599\ : CascadeMux
    port map (
            O => \N__37203\,
            I => \N__37153\
        );

    \I__8598\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37146\
        );

    \I__8597\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37146\
        );

    \I__8596\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37146\
        );

    \I__8595\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37142\
        );

    \I__8594\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37139\
        );

    \I__8593\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37136\
        );

    \I__8592\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37133\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__37191\,
            I => \N__37130\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__37188\,
            I => \N__37125\
        );

    \I__8589\ : Span4Mux_h
    port map (
            O => \N__37183\,
            I => \N__37125\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__37180\,
            I => \N__37122\
        );

    \I__8587\ : Span4Mux_h
    port map (
            O => \N__37177\,
            I => \N__37119\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__37174\,
            I => \N__37105\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__37169\,
            I => \N__37105\
        );

    \I__8584\ : Span4Mux_v
    port map (
            O => \N__37164\,
            I => \N__37105\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__37159\,
            I => \N__37105\
        );

    \I__8582\ : CascadeMux
    port map (
            O => \N__37158\,
            I => \N__37102\
        );

    \I__8581\ : CascadeMux
    port map (
            O => \N__37157\,
            I => \N__37099\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__37156\,
            I => \N__37095\
        );

    \I__8579\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37091\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__37146\,
            I => \N__37088\
        );

    \I__8577\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37085\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37080\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__37139\,
            I => \N__37080\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__37136\,
            I => \N__37077\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__37133\,
            I => \N__37074\
        );

    \I__8572\ : Span4Mux_h
    port map (
            O => \N__37130\,
            I => \N__37069\
        );

    \I__8571\ : Span4Mux_v
    port map (
            O => \N__37125\,
            I => \N__37069\
        );

    \I__8570\ : Span4Mux_v
    port map (
            O => \N__37122\,
            I => \N__37064\
        );

    \I__8569\ : Span4Mux_h
    port map (
            O => \N__37119\,
            I => \N__37064\
        );

    \I__8568\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37059\
        );

    \I__8567\ : InMux
    port map (
            O => \N__37117\,
            I => \N__37059\
        );

    \I__8566\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37052\
        );

    \I__8565\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37052\
        );

    \I__8564\ : InMux
    port map (
            O => \N__37114\,
            I => \N__37052\
        );

    \I__8563\ : Span4Mux_h
    port map (
            O => \N__37105\,
            I => \N__37049\
        );

    \I__8562\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37044\
        );

    \I__8561\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37044\
        );

    \I__8560\ : InMux
    port map (
            O => \N__37098\,
            I => \N__37037\
        );

    \I__8559\ : InMux
    port map (
            O => \N__37095\,
            I => \N__37037\
        );

    \I__8558\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37037\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__37091\,
            I => \N__37030\
        );

    \I__8556\ : Span12Mux_s7_v
    port map (
            O => \N__37088\,
            I => \N__37030\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__37085\,
            I => \N__37030\
        );

    \I__8554\ : Span4Mux_s1_h
    port map (
            O => \N__37080\,
            I => \N__37021\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__37077\,
            I => \N__37021\
        );

    \I__8552\ : Span4Mux_v
    port map (
            O => \N__37074\,
            I => \N__37021\
        );

    \I__8551\ : Span4Mux_v
    port map (
            O => \N__37069\,
            I => \N__37021\
        );

    \I__8550\ : Odrv4
    port map (
            O => \N__37064\,
            I => \ALU.N_240_0\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__37059\,
            I => \ALU.N_240_0\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__37052\,
            I => \ALU.N_240_0\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__37049\,
            I => \ALU.N_240_0\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__37044\,
            I => \ALU.N_240_0\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__37037\,
            I => \ALU.N_240_0\
        );

    \I__8544\ : Odrv12
    port map (
            O => \N__37030\,
            I => \ALU.N_240_0\
        );

    \I__8543\ : Odrv4
    port map (
            O => \N__37021\,
            I => \ALU.N_240_0\
        );

    \I__8542\ : CascadeMux
    port map (
            O => \N__37004\,
            I => \N__36990\
        );

    \I__8541\ : CascadeMux
    port map (
            O => \N__37003\,
            I => \N__36986\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__37002\,
            I => \N__36976\
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__37001\,
            I => \N__36973\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__37000\,
            I => \N__36970\
        );

    \I__8537\ : CascadeMux
    port map (
            O => \N__36999\,
            I => \N__36967\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__36998\,
            I => \N__36959\
        );

    \I__8535\ : CascadeMux
    port map (
            O => \N__36997\,
            I => \N__36954\
        );

    \I__8534\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36949\
        );

    \I__8533\ : InMux
    port map (
            O => \N__36995\,
            I => \N__36946\
        );

    \I__8532\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36941\
        );

    \I__8531\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36933\
        );

    \I__8530\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36930\
        );

    \I__8529\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36925\
        );

    \I__8528\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36925\
        );

    \I__8527\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36922\
        );

    \I__8526\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36915\
        );

    \I__8525\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36915\
        );

    \I__8524\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36915\
        );

    \I__8523\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36912\
        );

    \I__8522\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36905\
        );

    \I__8521\ : InMux
    port map (
            O => \N__36979\,
            I => \N__36905\
        );

    \I__8520\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36905\
        );

    \I__8519\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36902\
        );

    \I__8518\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36897\
        );

    \I__8517\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36897\
        );

    \I__8516\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36890\
        );

    \I__8515\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36890\
        );

    \I__8514\ : InMux
    port map (
            O => \N__36964\,
            I => \N__36890\
        );

    \I__8513\ : InMux
    port map (
            O => \N__36963\,
            I => \N__36887\
        );

    \I__8512\ : InMux
    port map (
            O => \N__36962\,
            I => \N__36884\
        );

    \I__8511\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36879\
        );

    \I__8510\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36879\
        );

    \I__8509\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36875\
        );

    \I__8508\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36868\
        );

    \I__8507\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36868\
        );

    \I__8506\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36868\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__36949\,
            I => \N__36865\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__36946\,
            I => \N__36862\
        );

    \I__8503\ : CascadeMux
    port map (
            O => \N__36945\,
            I => \N__36858\
        );

    \I__8502\ : CascadeMux
    port map (
            O => \N__36944\,
            I => \N__36855\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36852\
        );

    \I__8500\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36845\
        );

    \I__8499\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36845\
        );

    \I__8498\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36845\
        );

    \I__8497\ : InMux
    port map (
            O => \N__36937\,
            I => \N__36839\
        );

    \I__8496\ : InMux
    port map (
            O => \N__36936\,
            I => \N__36839\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__36933\,
            I => \N__36836\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__36930\,
            I => \N__36833\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__36925\,
            I => \N__36828\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__36922\,
            I => \N__36828\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__36915\,
            I => \N__36825\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__36912\,
            I => \N__36820\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__36905\,
            I => \N__36820\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__36902\,
            I => \N__36817\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__36897\,
            I => \N__36814\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__36890\,
            I => \N__36804\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__36887\,
            I => \N__36804\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36804\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__36879\,
            I => \N__36804\
        );

    \I__8482\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36801\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__36875\,
            I => \N__36796\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36796\
        );

    \I__8479\ : Span4Mux_v
    port map (
            O => \N__36865\,
            I => \N__36791\
        );

    \I__8478\ : Span4Mux_v
    port map (
            O => \N__36862\,
            I => \N__36791\
        );

    \I__8477\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36784\
        );

    \I__8476\ : InMux
    port map (
            O => \N__36858\,
            I => \N__36784\
        );

    \I__8475\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36784\
        );

    \I__8474\ : Span4Mux_s2_h
    port map (
            O => \N__36852\,
            I => \N__36779\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36779\
        );

    \I__8472\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36776\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__36839\,
            I => \N__36773\
        );

    \I__8470\ : Span4Mux_h
    port map (
            O => \N__36836\,
            I => \N__36770\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__36833\,
            I => \N__36765\
        );

    \I__8468\ : Span4Mux_v
    port map (
            O => \N__36828\,
            I => \N__36765\
        );

    \I__8467\ : Span4Mux_h
    port map (
            O => \N__36825\,
            I => \N__36760\
        );

    \I__8466\ : Span4Mux_v
    port map (
            O => \N__36820\,
            I => \N__36760\
        );

    \I__8465\ : Span4Mux_h
    port map (
            O => \N__36817\,
            I => \N__36757\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__36814\,
            I => \N__36754\
        );

    \I__8463\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36751\
        );

    \I__8462\ : Span4Mux_v
    port map (
            O => \N__36804\,
            I => \N__36748\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__36801\,
            I => \N__36741\
        );

    \I__8460\ : Span4Mux_v
    port map (
            O => \N__36796\,
            I => \N__36741\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__36791\,
            I => \N__36741\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36734\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__36779\,
            I => \N__36734\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__36776\,
            I => \N__36734\
        );

    \I__8455\ : Span12Mux_s3_v
    port map (
            O => \N__36773\,
            I => \N__36731\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__36770\,
            I => \N__36728\
        );

    \I__8453\ : Span4Mux_h
    port map (
            O => \N__36765\,
            I => \N__36725\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__36760\,
            I => \N__36722\
        );

    \I__8451\ : Span4Mux_v
    port map (
            O => \N__36757\,
            I => \N__36709\
        );

    \I__8450\ : Span4Mux_h
    port map (
            O => \N__36754\,
            I => \N__36709\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__36751\,
            I => \N__36709\
        );

    \I__8448\ : Span4Mux_h
    port map (
            O => \N__36748\,
            I => \N__36709\
        );

    \I__8447\ : Span4Mux_v
    port map (
            O => \N__36741\,
            I => \N__36709\
        );

    \I__8446\ : Span4Mux_v
    port map (
            O => \N__36734\,
            I => \N__36709\
        );

    \I__8445\ : Odrv12
    port map (
            O => \N__36731\,
            I => \ALU.aluOut_2\
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__36728\,
            I => \ALU.aluOut_2\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__36725\,
            I => \ALU.aluOut_2\
        );

    \I__8442\ : Odrv4
    port map (
            O => \N__36722\,
            I => \ALU.aluOut_2\
        );

    \I__8441\ : Odrv4
    port map (
            O => \N__36709\,
            I => \ALU.aluOut_2\
        );

    \I__8440\ : InMux
    port map (
            O => \N__36698\,
            I => \ALU.un9_addsub_cry_1\
        );

    \I__8439\ : CascadeMux
    port map (
            O => \N__36695\,
            I => \N__36692\
        );

    \I__8438\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36689\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36686\
        );

    \I__8436\ : Span12Mux_h
    port map (
            O => \N__36686\,
            I => \N__36683\
        );

    \I__8435\ : Odrv12
    port map (
            O => \N__36683\,
            I => \ALU.N_237_0_i\
        );

    \I__8434\ : InMux
    port map (
            O => \N__36680\,
            I => \ALU.un9_addsub_cry_2\
        );

    \I__8433\ : CascadeMux
    port map (
            O => \N__36677\,
            I => \N__36674\
        );

    \I__8432\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36671\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36668\
        );

    \I__8430\ : Odrv12
    port map (
            O => \N__36668\,
            I => \ALU.N_231_0_i\
        );

    \I__8429\ : InMux
    port map (
            O => \N__36665\,
            I => \ALU.un9_addsub_cry_3\
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__36662\,
            I => \N__36659\
        );

    \I__8427\ : InMux
    port map (
            O => \N__36659\,
            I => \N__36656\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36653\
        );

    \I__8425\ : Span4Mux_h
    port map (
            O => \N__36653\,
            I => \N__36650\
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__36650\,
            I => \ALU.madd_axb_0_l_ofx\
        );

    \I__8423\ : CascadeMux
    port map (
            O => \N__36647\,
            I => \ALU.mult_1_cascade_\
        );

    \I__8422\ : InMux
    port map (
            O => \N__36644\,
            I => \N__36641\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__36641\,
            I => \N__36638\
        );

    \I__8420\ : Span4Mux_v
    port map (
            O => \N__36638\,
            I => \N__36635\
        );

    \I__8419\ : Span4Mux_h
    port map (
            O => \N__36635\,
            I => \N__36632\
        );

    \I__8418\ : Span4Mux_v
    port map (
            O => \N__36632\,
            I => \N__36629\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__36629\,
            I => \ALU.a_15_m5_1\
        );

    \I__8416\ : CascadeMux
    port map (
            O => \N__36626\,
            I => \ALU.d_RNIEICQ63Z0Z_1_cascade_\
        );

    \I__8415\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36617\
        );

    \I__8414\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36617\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__36617\,
            I => \ALU.bZ0Z_1\
        );

    \I__8412\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36610\
        );

    \I__8411\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36607\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__36610\,
            I => \N__36602\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__36607\,
            I => \N__36599\
        );

    \I__8408\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36596\
        );

    \I__8407\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36593\
        );

    \I__8406\ : Span4Mux_h
    port map (
            O => \N__36602\,
            I => \N__36587\
        );

    \I__8405\ : Span4Mux_h
    port map (
            O => \N__36599\,
            I => \N__36584\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__36596\,
            I => \N__36581\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36578\
        );

    \I__8402\ : InMux
    port map (
            O => \N__36592\,
            I => \N__36575\
        );

    \I__8401\ : InMux
    port map (
            O => \N__36591\,
            I => \N__36572\
        );

    \I__8400\ : InMux
    port map (
            O => \N__36590\,
            I => \N__36569\
        );

    \I__8399\ : Odrv4
    port map (
            O => \N__36587\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__36584\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8397\ : Odrv4
    port map (
            O => \N__36581\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8396\ : Odrv12
    port map (
            O => \N__36578\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__36575\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__36572\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__36569\,
            I => \ALU.d_RNIEICQ63Z0Z_1\
        );

    \I__8392\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36548\
        );

    \I__8391\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36548\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__36545\,
            I => \ALU.dZ0Z_1\
        );

    \I__8388\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36539\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__36539\,
            I => \N__36536\
        );

    \I__8386\ : Span4Mux_h
    port map (
            O => \N__36536\,
            I => \N__36532\
        );

    \I__8385\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36529\
        );

    \I__8384\ : Span4Mux_h
    port map (
            O => \N__36532\,
            I => \N__36526\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__36529\,
            I => \N__36523\
        );

    \I__8382\ : Odrv4
    port map (
            O => \N__36526\,
            I => \ALU.hZ0Z_4\
        );

    \I__8381\ : Odrv12
    port map (
            O => \N__36523\,
            I => \ALU.hZ0Z_4\
        );

    \I__8380\ : InMux
    port map (
            O => \N__36518\,
            I => \N__36514\
        );

    \I__8379\ : InMux
    port map (
            O => \N__36517\,
            I => \N__36511\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__36514\,
            I => \FTDI.un3_TX_0_i\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__36511\,
            I => \FTDI.un3_TX_0_i\
        );

    \I__8376\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36503\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__36503\,
            I => \FTDI.un3_TX_axb_3\
        );

    \I__8374\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36497\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__36497\,
            I => \N__36494\
        );

    \I__8372\ : Span4Mux_s2_v
    port map (
            O => \N__36494\,
            I => \N__36491\
        );

    \I__8371\ : Odrv4
    port map (
            O => \N__36491\,
            I => \FTDI.TXshiftZ0Z_0\
        );

    \I__8370\ : InMux
    port map (
            O => \N__36488\,
            I => \FTDI.un3_TX_cry_3\
        );

    \I__8369\ : IoInMux
    port map (
            O => \N__36485\,
            I => \N__36482\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__36482\,
            I => \N__36479\
        );

    \I__8367\ : Span4Mux_s1_v
    port map (
            O => \N__36479\,
            I => \N__36476\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__36476\,
            I => \N__36473\
        );

    \I__8365\ : Span4Mux_h
    port map (
            O => \N__36473\,
            I => \N__36470\
        );

    \I__8364\ : Odrv4
    port map (
            O => \N__36470\,
            I => \FTDI_TX_0_i\
        );

    \I__8363\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36461\
        );

    \I__8362\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36461\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__36461\,
            I => \ALU.fZ0Z_1\
        );

    \I__8360\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__36455\,
            I => \N__36452\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__36452\,
            I => \N__36448\
        );

    \I__8357\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36445\
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__36448\,
            I => \ALU.fZ0Z_2\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__36445\,
            I => \ALU.fZ0Z_2\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__36440\,
            I => \N__36437\
        );

    \I__8353\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36434\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36430\
        );

    \I__8351\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36427\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__36430\,
            I => \N__36424\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__36427\,
            I => \ALU.fZ0Z_5\
        );

    \I__8348\ : Odrv4
    port map (
            O => \N__36424\,
            I => \ALU.fZ0Z_5\
        );

    \I__8347\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36416\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__36416\,
            I => \N__36412\
        );

    \I__8345\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36409\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__36412\,
            I => \N__36406\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__36409\,
            I => \N__36403\
        );

    \I__8342\ : Span4Mux_h
    port map (
            O => \N__36406\,
            I => \N__36400\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__36403\,
            I => \ALU.fZ0Z_6\
        );

    \I__8340\ : Odrv4
    port map (
            O => \N__36400\,
            I => \ALU.fZ0Z_6\
        );

    \I__8339\ : CascadeMux
    port map (
            O => \N__36395\,
            I => \N__36392\
        );

    \I__8338\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__8337\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36386\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__36386\,
            I => \N__36383\
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__36383\,
            I => \ALU.fZ0Z_7\
        );

    \I__8334\ : CEMux
    port map (
            O => \N__36380\,
            I => \N__36377\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__36377\,
            I => \N__36373\
        );

    \I__8332\ : CEMux
    port map (
            O => \N__36376\,
            I => \N__36370\
        );

    \I__8331\ : Span4Mux_v
    port map (
            O => \N__36373\,
            I => \N__36367\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__36370\,
            I => \N__36364\
        );

    \I__8329\ : Span4Mux_v
    port map (
            O => \N__36367\,
            I => \N__36360\
        );

    \I__8328\ : Span4Mux_v
    port map (
            O => \N__36364\,
            I => \N__36357\
        );

    \I__8327\ : CEMux
    port map (
            O => \N__36363\,
            I => \N__36354\
        );

    \I__8326\ : Span4Mux_h
    port map (
            O => \N__36360\,
            I => \N__36351\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__36357\,
            I => \N__36348\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__36354\,
            I => \N__36345\
        );

    \I__8323\ : Span4Mux_h
    port map (
            O => \N__36351\,
            I => \N__36342\
        );

    \I__8322\ : Sp12to4
    port map (
            O => \N__36348\,
            I => \N__36339\
        );

    \I__8321\ : Span4Mux_h
    port map (
            O => \N__36345\,
            I => \N__36336\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__36342\,
            I => \ALU.f_cnvZ0Z_0\
        );

    \I__8319\ : Odrv12
    port map (
            O => \N__36339\,
            I => \ALU.f_cnvZ0Z_0\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__36336\,
            I => \ALU.f_cnvZ0Z_0\
        );

    \I__8317\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36326\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__36326\,
            I => \N__36322\
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__36325\,
            I => \N__36319\
        );

    \I__8314\ : Span4Mux_h
    port map (
            O => \N__36322\,
            I => \N__36316\
        );

    \I__8313\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36313\
        );

    \I__8312\ : Span4Mux_v
    port map (
            O => \N__36316\,
            I => \N__36308\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__36313\,
            I => \N__36308\
        );

    \I__8310\ : Span4Mux_h
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__36305\,
            I => \ALU.N_1700_i\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__36302\,
            I => \ALU.d_RNIO75MAZ0Z_0_cascade_\
        );

    \I__8307\ : CascadeMux
    port map (
            O => \N__36299\,
            I => \N__36296\
        );

    \I__8306\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36293\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__36293\,
            I => \N__36290\
        );

    \I__8304\ : Span4Mux_h
    port map (
            O => \N__36290\,
            I => \N__36287\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__36287\,
            I => \N__36283\
        );

    \I__8302\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36280\
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__36283\,
            I => \ALU.bZ0Z_0\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__36280\,
            I => \ALU.bZ0Z_0\
        );

    \I__8299\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36272\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__36272\,
            I => \N__36269\
        );

    \I__8297\ : Span4Mux_v
    port map (
            O => \N__36269\,
            I => \N__36265\
        );

    \I__8296\ : InMux
    port map (
            O => \N__36268\,
            I => \N__36261\
        );

    \I__8295\ : Span4Mux_h
    port map (
            O => \N__36265\,
            I => \N__36254\
        );

    \I__8294\ : InMux
    port map (
            O => \N__36264\,
            I => \N__36251\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__36261\,
            I => \N__36248\
        );

    \I__8292\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36245\
        );

    \I__8291\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36242\
        );

    \I__8290\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36239\
        );

    \I__8289\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36236\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__36254\,
            I => \N__36231\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__36251\,
            I => \N__36231\
        );

    \I__8286\ : Span4Mux_h
    port map (
            O => \N__36248\,
            I => \N__36228\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__36245\,
            I => \N__36223\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36223\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__36239\,
            I => \N__36218\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__36236\,
            I => \N__36218\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__36231\,
            I => \ALU.a_15_ns_1_9\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__36228\,
            I => \ALU.a_15_ns_1_9\
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__36223\,
            I => \ALU.a_15_ns_1_9\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__36218\,
            I => \ALU.a_15_ns_1_9\
        );

    \I__8277\ : CascadeMux
    port map (
            O => \N__36209\,
            I => \N__36206\
        );

    \I__8276\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36199\
        );

    \I__8275\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36196\
        );

    \I__8274\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36191\
        );

    \I__8273\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36188\
        );

    \I__8272\ : CascadeMux
    port map (
            O => \N__36202\,
            I => \N__36185\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__36182\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__36196\,
            I => \N__36179\
        );

    \I__8269\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36175\
        );

    \I__8268\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36172\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__36191\,
            I => \N__36167\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36167\
        );

    \I__8265\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36164\
        );

    \I__8264\ : Span4Mux_v
    port map (
            O => \N__36182\,
            I => \N__36161\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__36179\,
            I => \N__36158\
        );

    \I__8262\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36155\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__36175\,
            I => \N__36152\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__36172\,
            I => \N__36147\
        );

    \I__8259\ : Span4Mux_h
    port map (
            O => \N__36167\,
            I => \N__36147\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__36164\,
            I => \N__36140\
        );

    \I__8257\ : Span4Mux_h
    port map (
            O => \N__36161\,
            I => \N__36140\
        );

    \I__8256\ : Span4Mux_v
    port map (
            O => \N__36158\,
            I => \N__36140\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__36155\,
            I => \ALU.mult_9\
        );

    \I__8254\ : Odrv4
    port map (
            O => \N__36152\,
            I => \ALU.mult_9\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__36147\,
            I => \ALU.mult_9\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__36140\,
            I => \ALU.mult_9\
        );

    \I__8251\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36128\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__36128\,
            I => \N__36125\
        );

    \I__8249\ : Span4Mux_h
    port map (
            O => \N__36125\,
            I => \N__36120\
        );

    \I__8248\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36115\
        );

    \I__8247\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36115\
        );

    \I__8246\ : Span4Mux_h
    port map (
            O => \N__36120\,
            I => \N__36112\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36109\
        );

    \I__8244\ : Odrv4
    port map (
            O => \N__36112\,
            I => \ALU.gZ0Z_9\
        );

    \I__8243\ : Odrv12
    port map (
            O => \N__36109\,
            I => \ALU.gZ0Z_9\
        );

    \I__8242\ : CEMux
    port map (
            O => \N__36104\,
            I => \N__36101\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__36101\,
            I => \N__36097\
        );

    \I__8240\ : CEMux
    port map (
            O => \N__36100\,
            I => \N__36094\
        );

    \I__8239\ : Span4Mux_v
    port map (
            O => \N__36097\,
            I => \N__36090\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__36094\,
            I => \N__36087\
        );

    \I__8237\ : CEMux
    port map (
            O => \N__36093\,
            I => \N__36084\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__36090\,
            I => \N__36081\
        );

    \I__8235\ : Span4Mux_v
    port map (
            O => \N__36087\,
            I => \N__36076\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__36084\,
            I => \N__36076\
        );

    \I__8233\ : Span4Mux_h
    port map (
            O => \N__36081\,
            I => \N__36073\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__36076\,
            I => \N__36070\
        );

    \I__8231\ : Span4Mux_v
    port map (
            O => \N__36073\,
            I => \N__36066\
        );

    \I__8230\ : Span4Mux_h
    port map (
            O => \N__36070\,
            I => \N__36063\
        );

    \I__8229\ : CEMux
    port map (
            O => \N__36069\,
            I => \N__36060\
        );

    \I__8228\ : Span4Mux_v
    port map (
            O => \N__36066\,
            I => \N__36057\
        );

    \I__8227\ : Sp12to4
    port map (
            O => \N__36063\,
            I => \N__36054\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__36060\,
            I => \N__36051\
        );

    \I__8225\ : Sp12to4
    port map (
            O => \N__36057\,
            I => \N__36046\
        );

    \I__8224\ : Span12Mux_v
    port map (
            O => \N__36054\,
            I => \N__36046\
        );

    \I__8223\ : Span4Mux_v
    port map (
            O => \N__36051\,
            I => \N__36043\
        );

    \I__8222\ : Odrv12
    port map (
            O => \N__36046\,
            I => \ALU.g_cnvZ0Z_0\
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__36043\,
            I => \ALU.g_cnvZ0Z_0\
        );

    \I__8220\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36035\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__36032\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__36032\,
            I => \N__36028\
        );

    \I__8217\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36025\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__36028\,
            I => \ALU.eZ0Z_13\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__36025\,
            I => \ALU.eZ0Z_13\
        );

    \I__8214\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36016\
        );

    \I__8213\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36013\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__36016\,
            I => \N__36010\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__36013\,
            I => \ALU.aZ0Z_13\
        );

    \I__8210\ : Odrv4
    port map (
            O => \N__36010\,
            I => \ALU.aZ0Z_13\
        );

    \I__8209\ : CascadeMux
    port map (
            O => \N__36005\,
            I => \N__36000\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__36004\,
            I => \N__35997\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__36003\,
            I => \N__35993\
        );

    \I__8206\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35990\
        );

    \I__8205\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35986\
        );

    \I__8204\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35982\
        );

    \I__8203\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35979\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35976\
        );

    \I__8201\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35973\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__35986\,
            I => \N__35970\
        );

    \I__8199\ : CascadeMux
    port map (
            O => \N__35985\,
            I => \N__35967\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35962\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__35979\,
            I => \N__35959\
        );

    \I__8196\ : Span4Mux_v
    port map (
            O => \N__35976\,
            I => \N__35954\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__35973\,
            I => \N__35954\
        );

    \I__8194\ : Span4Mux_v
    port map (
            O => \N__35970\,
            I => \N__35951\
        );

    \I__8193\ : InMux
    port map (
            O => \N__35967\,
            I => \N__35948\
        );

    \I__8192\ : CascadeMux
    port map (
            O => \N__35966\,
            I => \N__35945\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__35965\,
            I => \N__35942\
        );

    \I__8190\ : Span4Mux_v
    port map (
            O => \N__35962\,
            I => \N__35937\
        );

    \I__8189\ : Span4Mux_v
    port map (
            O => \N__35959\,
            I => \N__35937\
        );

    \I__8188\ : Span4Mux_h
    port map (
            O => \N__35954\,
            I => \N__35934\
        );

    \I__8187\ : Span4Mux_h
    port map (
            O => \N__35951\,
            I => \N__35931\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__35948\,
            I => \N__35928\
        );

    \I__8185\ : InMux
    port map (
            O => \N__35945\,
            I => \N__35923\
        );

    \I__8184\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35923\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__35937\,
            I => \aluOperand1_2_rep2\
        );

    \I__8182\ : Odrv4
    port map (
            O => \N__35934\,
            I => \aluOperand1_2_rep2\
        );

    \I__8181\ : Odrv4
    port map (
            O => \N__35931\,
            I => \aluOperand1_2_rep2\
        );

    \I__8180\ : Odrv12
    port map (
            O => \N__35928\,
            I => \aluOperand1_2_rep2\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__35923\,
            I => \aluOperand1_2_rep2\
        );

    \I__8178\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35907\
        );

    \I__8177\ : CascadeMux
    port map (
            O => \N__35911\,
            I => \N__35903\
        );

    \I__8176\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35900\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__35907\,
            I => \N__35894\
        );

    \I__8174\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35889\
        );

    \I__8173\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35889\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__35900\,
            I => \N__35886\
        );

    \I__8171\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35883\
        );

    \I__8170\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35880\
        );

    \I__8169\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35877\
        );

    \I__8168\ : Span4Mux_h
    port map (
            O => \N__35894\,
            I => \N__35872\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__35889\,
            I => \N__35863\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__35886\,
            I => \N__35863\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__35883\,
            I => \N__35863\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35860\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__35877\,
            I => \N__35857\
        );

    \I__8162\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35854\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__35875\,
            I => \N__35849\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__35872\,
            I => \N__35846\
        );

    \I__8159\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35841\
        );

    \I__8158\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35841\
        );

    \I__8157\ : Span4Mux_h
    port map (
            O => \N__35863\,
            I => \N__35838\
        );

    \I__8156\ : Span4Mux_h
    port map (
            O => \N__35860\,
            I => \N__35833\
        );

    \I__8155\ : Span4Mux_h
    port map (
            O => \N__35857\,
            I => \N__35833\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__35854\,
            I => \N__35830\
        );

    \I__8153\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35823\
        );

    \I__8152\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35823\
        );

    \I__8151\ : InMux
    port map (
            O => \N__35849\,
            I => \N__35823\
        );

    \I__8150\ : Odrv4
    port map (
            O => \N__35846\,
            I => \aluOperand1_1_rep1\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__35841\,
            I => \aluOperand1_1_rep1\
        );

    \I__8148\ : Odrv4
    port map (
            O => \N__35838\,
            I => \aluOperand1_1_rep1\
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__35833\,
            I => \aluOperand1_1_rep1\
        );

    \I__8146\ : Odrv12
    port map (
            O => \N__35830\,
            I => \aluOperand1_1_rep1\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__35823\,
            I => \aluOperand1_1_rep1\
        );

    \I__8144\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35806\
        );

    \I__8143\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35803\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__35806\,
            I => \ALU.cZ0Z_13\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__35803\,
            I => \ALU.cZ0Z_13\
        );

    \I__8140\ : CascadeMux
    port map (
            O => \N__35798\,
            I => \ALU.dout_3_ns_1_13_cascade_\
        );

    \I__8139\ : InMux
    port map (
            O => \N__35795\,
            I => \N__35791\
        );

    \I__8138\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35788\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__35791\,
            I => \ALU.gZ0Z_13\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__35788\,
            I => \ALU.gZ0Z_13\
        );

    \I__8135\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35776\
        );

    \I__8134\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35776\
        );

    \I__8133\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35773\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__35776\,
            I => \N__35770\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__35773\,
            I => \N__35767\
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__35770\,
            I => \ALU.bZ0Z_13\
        );

    \I__8129\ : Odrv4
    port map (
            O => \N__35767\,
            I => \ALU.bZ0Z_13\
        );

    \I__8128\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35758\
        );

    \I__8127\ : InMux
    port map (
            O => \N__35761\,
            I => \N__35755\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35749\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35745\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__35754\,
            I => \N__35742\
        );

    \I__8123\ : CascadeMux
    port map (
            O => \N__35753\,
            I => \N__35739\
        );

    \I__8122\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35734\
        );

    \I__8121\ : Span4Mux_h
    port map (
            O => \N__35749\,
            I => \N__35731\
        );

    \I__8120\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35728\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__35745\,
            I => \N__35725\
        );

    \I__8118\ : InMux
    port map (
            O => \N__35742\,
            I => \N__35720\
        );

    \I__8117\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35720\
        );

    \I__8116\ : CascadeMux
    port map (
            O => \N__35738\,
            I => \N__35717\
        );

    \I__8115\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35714\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__35734\,
            I => \N__35710\
        );

    \I__8113\ : Span4Mux_v
    port map (
            O => \N__35731\,
            I => \N__35703\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__35728\,
            I => \N__35700\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__35725\,
            I => \N__35695\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35692\
        );

    \I__8109\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35689\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__35714\,
            I => \N__35686\
        );

    \I__8107\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35683\
        );

    \I__8106\ : Span4Mux_h
    port map (
            O => \N__35710\,
            I => \N__35680\
        );

    \I__8105\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35677\
        );

    \I__8104\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35672\
        );

    \I__8103\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35672\
        );

    \I__8102\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35668\
        );

    \I__8101\ : Span4Mux_v
    port map (
            O => \N__35703\,
            I => \N__35663\
        );

    \I__8100\ : Span4Mux_v
    port map (
            O => \N__35700\,
            I => \N__35663\
        );

    \I__8099\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35658\
        );

    \I__8098\ : InMux
    port map (
            O => \N__35698\,
            I => \N__35658\
        );

    \I__8097\ : Span4Mux_v
    port map (
            O => \N__35695\,
            I => \N__35653\
        );

    \I__8096\ : Span4Mux_h
    port map (
            O => \N__35692\,
            I => \N__35653\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35648\
        );

    \I__8094\ : Span4Mux_v
    port map (
            O => \N__35686\,
            I => \N__35648\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35645\
        );

    \I__8092\ : Span4Mux_h
    port map (
            O => \N__35680\,
            I => \N__35638\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__35677\,
            I => \N__35638\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__35672\,
            I => \N__35638\
        );

    \I__8089\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35635\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__35668\,
            I => \N__35632\
        );

    \I__8087\ : Odrv4
    port map (
            O => \N__35663\,
            I => \aluOperand1_1_rep2\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__35658\,
            I => \aluOperand1_1_rep2\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__35653\,
            I => \aluOperand1_1_rep2\
        );

    \I__8084\ : Odrv4
    port map (
            O => \N__35648\,
            I => \aluOperand1_1_rep2\
        );

    \I__8083\ : Odrv12
    port map (
            O => \N__35645\,
            I => \aluOperand1_1_rep2\
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__35638\,
            I => \aluOperand1_1_rep2\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__35635\,
            I => \aluOperand1_1_rep2\
        );

    \I__8080\ : Odrv4
    port map (
            O => \N__35632\,
            I => \aluOperand1_1_rep2\
        );

    \I__8079\ : CascadeMux
    port map (
            O => \N__35615\,
            I => \N__35611\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__35614\,
            I => \N__35608\
        );

    \I__8077\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35604\
        );

    \I__8076\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35599\
        );

    \I__8075\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35599\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35596\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35591\
        );

    \I__8072\ : Span4Mux_v
    port map (
            O => \N__35596\,
            I => \N__35591\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__35591\,
            I => \ALU.fZ0Z_13\
        );

    \I__8070\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35583\
        );

    \I__8069\ : CascadeMux
    port map (
            O => \N__35587\,
            I => \N__35578\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__35586\,
            I => \N__35573\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__35583\,
            I => \N__35570\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__35582\,
            I => \N__35567\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__35581\,
            I => \N__35564\
        );

    \I__8064\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35561\
        );

    \I__8063\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35558\
        );

    \I__8062\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35555\
        );

    \I__8061\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35551\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__35570\,
            I => \N__35548\
        );

    \I__8059\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35545\
        );

    \I__8058\ : InMux
    port map (
            O => \N__35564\,
            I => \N__35542\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35539\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__35558\,
            I => \N__35536\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__35555\,
            I => \N__35533\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__35554\,
            I => \N__35528\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35525\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__35548\,
            I => \N__35522\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__35545\,
            I => \N__35519\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__35542\,
            I => \N__35516\
        );

    \I__8049\ : Span4Mux_h
    port map (
            O => \N__35539\,
            I => \N__35513\
        );

    \I__8048\ : Span4Mux_v
    port map (
            O => \N__35536\,
            I => \N__35510\
        );

    \I__8047\ : Span4Mux_h
    port map (
            O => \N__35533\,
            I => \N__35507\
        );

    \I__8046\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35504\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__35531\,
            I => \N__35501\
        );

    \I__8044\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35498\
        );

    \I__8043\ : Span4Mux_h
    port map (
            O => \N__35525\,
            I => \N__35495\
        );

    \I__8042\ : Span4Mux_v
    port map (
            O => \N__35522\,
            I => \N__35488\
        );

    \I__8041\ : Span4Mux_v
    port map (
            O => \N__35519\,
            I => \N__35488\
        );

    \I__8040\ : Span4Mux_v
    port map (
            O => \N__35516\,
            I => \N__35488\
        );

    \I__8039\ : Span4Mux_v
    port map (
            O => \N__35513\,
            I => \N__35483\
        );

    \I__8038\ : Span4Mux_h
    port map (
            O => \N__35510\,
            I => \N__35483\
        );

    \I__8037\ : Span4Mux_v
    port map (
            O => \N__35507\,
            I => \N__35478\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__35504\,
            I => \N__35478\
        );

    \I__8035\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35475\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__35498\,
            I => \aluOperand1_2\
        );

    \I__8033\ : Odrv4
    port map (
            O => \N__35495\,
            I => \aluOperand1_2\
        );

    \I__8032\ : Odrv4
    port map (
            O => \N__35488\,
            I => \aluOperand1_2\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__35483\,
            I => \aluOperand1_2\
        );

    \I__8030\ : Odrv4
    port map (
            O => \N__35478\,
            I => \aluOperand1_2\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__35475\,
            I => \aluOperand1_2\
        );

    \I__8028\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35458\
        );

    \I__8027\ : InMux
    port map (
            O => \N__35461\,
            I => \N__35455\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35452\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__35455\,
            I => \N__35447\
        );

    \I__8024\ : Span4Mux_v
    port map (
            O => \N__35452\,
            I => \N__35447\
        );

    \I__8023\ : Span4Mux_h
    port map (
            O => \N__35447\,
            I => \N__35443\
        );

    \I__8022\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35440\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__35443\,
            I => \ALU.hZ0Z_13\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__35440\,
            I => \ALU.hZ0Z_13\
        );

    \I__8019\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35431\
        );

    \I__8018\ : InMux
    port map (
            O => \N__35434\,
            I => \N__35428\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__35431\,
            I => \N__35425\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__35428\,
            I => \N__35421\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__35425\,
            I => \N__35418\
        );

    \I__8014\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35415\
        );

    \I__8013\ : Span4Mux_h
    port map (
            O => \N__35421\,
            I => \N__35410\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__35418\,
            I => \N__35410\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__35415\,
            I => \ALU.dZ0Z_13\
        );

    \I__8010\ : Odrv4
    port map (
            O => \N__35410\,
            I => \ALU.dZ0Z_13\
        );

    \I__8009\ : CascadeMux
    port map (
            O => \N__35405\,
            I => \ALU.dout_6_ns_1_13_cascade_\
        );

    \I__8008\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35396\
        );

    \I__8007\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35396\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__35396\,
            I => \N__35391\
        );

    \I__8005\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35386\
        );

    \I__8004\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35386\
        );

    \I__8003\ : Span4Mux_v
    port map (
            O => \N__35391\,
            I => \N__35379\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__35386\,
            I => \N__35379\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__35385\,
            I => \N__35371\
        );

    \I__8000\ : CascadeMux
    port map (
            O => \N__35384\,
            I => \N__35368\
        );

    \I__7999\ : Span4Mux_v
    port map (
            O => \N__35379\,
            I => \N__35362\
        );

    \I__7998\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35357\
        );

    \I__7997\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35357\
        );

    \I__7996\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35353\
        );

    \I__7995\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35347\
        );

    \I__7994\ : InMux
    port map (
            O => \N__35374\,
            I => \N__35347\
        );

    \I__7993\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35344\
        );

    \I__7992\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35341\
        );

    \I__7991\ : InMux
    port map (
            O => \N__35367\,
            I => \N__35338\
        );

    \I__7990\ : InMux
    port map (
            O => \N__35366\,
            I => \N__35335\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__35365\,
            I => \N__35332\
        );

    \I__7988\ : Span4Mux_h
    port map (
            O => \N__35362\,
            I => \N__35329\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__35357\,
            I => \N__35326\
        );

    \I__7986\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35323\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35320\
        );

    \I__7984\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35317\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__35347\,
            I => \N__35314\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__35344\,
            I => \N__35311\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__35341\,
            I => \N__35308\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__35338\,
            I => \N__35303\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__35335\,
            I => \N__35303\
        );

    \I__7978\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35300\
        );

    \I__7977\ : Span4Mux_h
    port map (
            O => \N__35329\,
            I => \N__35294\
        );

    \I__7976\ : Span4Mux_h
    port map (
            O => \N__35326\,
            I => \N__35289\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__35323\,
            I => \N__35289\
        );

    \I__7974\ : Span4Mux_v
    port map (
            O => \N__35320\,
            I => \N__35280\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__35317\,
            I => \N__35280\
        );

    \I__7972\ : Span4Mux_v
    port map (
            O => \N__35314\,
            I => \N__35280\
        );

    \I__7971\ : Span4Mux_v
    port map (
            O => \N__35311\,
            I => \N__35280\
        );

    \I__7970\ : Span4Mux_v
    port map (
            O => \N__35308\,
            I => \N__35275\
        );

    \I__7969\ : Span4Mux_v
    port map (
            O => \N__35303\,
            I => \N__35275\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__35300\,
            I => \N__35272\
        );

    \I__7967\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35265\
        );

    \I__7966\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35265\
        );

    \I__7965\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35265\
        );

    \I__7964\ : Odrv4
    port map (
            O => \N__35294\,
            I => \aluOperand1_1\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__35289\,
            I => \aluOperand1_1\
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__35280\,
            I => \aluOperand1_1\
        );

    \I__7961\ : Odrv4
    port map (
            O => \N__35275\,
            I => \aluOperand1_1\
        );

    \I__7960\ : Odrv12
    port map (
            O => \N__35272\,
            I => \aluOperand1_1\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__35265\,
            I => \aluOperand1_1\
        );

    \I__7958\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__35249\,
            I => \ALU.N_712\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__35246\,
            I => \ALU.N_760_cascade_\
        );

    \I__7955\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35236\
        );

    \I__7954\ : InMux
    port map (
            O => \N__35242\,
            I => \N__35236\
        );

    \I__7953\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35233\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__35236\,
            I => \N__35226\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__35233\,
            I => \N__35217\
        );

    \I__7950\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35214\
        );

    \I__7949\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35211\
        );

    \I__7948\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35208\
        );

    \I__7947\ : InMux
    port map (
            O => \N__35229\,
            I => \N__35203\
        );

    \I__7946\ : Span4Mux_v
    port map (
            O => \N__35226\,
            I => \N__35199\
        );

    \I__7945\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35196\
        );

    \I__7944\ : InMux
    port map (
            O => \N__35224\,
            I => \N__35193\
        );

    \I__7943\ : InMux
    port map (
            O => \N__35223\,
            I => \N__35190\
        );

    \I__7942\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35187\
        );

    \I__7941\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35184\
        );

    \I__7940\ : InMux
    port map (
            O => \N__35220\,
            I => \N__35180\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__35217\,
            I => \N__35175\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__35214\,
            I => \N__35175\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35170\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__35208\,
            I => \N__35170\
        );

    \I__7935\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35167\
        );

    \I__7934\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35164\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35161\
        );

    \I__7932\ : InMux
    port map (
            O => \N__35202\,
            I => \N__35158\
        );

    \I__7931\ : Span4Mux_v
    port map (
            O => \N__35199\,
            I => \N__35151\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__35196\,
            I => \N__35151\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__35193\,
            I => \N__35151\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__35190\,
            I => \N__35148\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__35187\,
            I => \N__35145\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__35184\,
            I => \N__35142\
        );

    \I__7925\ : InMux
    port map (
            O => \N__35183\,
            I => \N__35139\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35136\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__35175\,
            I => \N__35125\
        );

    \I__7922\ : Span4Mux_v
    port map (
            O => \N__35170\,
            I => \N__35125\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__35167\,
            I => \N__35125\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__35164\,
            I => \N__35125\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__35161\,
            I => \N__35122\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__35158\,
            I => \N__35119\
        );

    \I__7917\ : Span4Mux_h
    port map (
            O => \N__35151\,
            I => \N__35116\
        );

    \I__7916\ : Span12Mux_v
    port map (
            O => \N__35148\,
            I => \N__35113\
        );

    \I__7915\ : Span12Mux_v
    port map (
            O => \N__35145\,
            I => \N__35110\
        );

    \I__7914\ : Span4Mux_h
    port map (
            O => \N__35142\,
            I => \N__35107\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35102\
        );

    \I__7912\ : Span4Mux_v
    port map (
            O => \N__35136\,
            I => \N__35102\
        );

    \I__7911\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35097\
        );

    \I__7910\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35097\
        );

    \I__7909\ : Span4Mux_h
    port map (
            O => \N__35125\,
            I => \N__35094\
        );

    \I__7908\ : Span4Mux_h
    port map (
            O => \N__35122\,
            I => \N__35087\
        );

    \I__7907\ : Span4Mux_v
    port map (
            O => \N__35119\,
            I => \N__35087\
        );

    \I__7906\ : Span4Mux_v
    port map (
            O => \N__35116\,
            I => \N__35087\
        );

    \I__7905\ : Odrv12
    port map (
            O => \N__35113\,
            I => \aluOperand1_0\
        );

    \I__7904\ : Odrv12
    port map (
            O => \N__35110\,
            I => \aluOperand1_0\
        );

    \I__7903\ : Odrv4
    port map (
            O => \N__35107\,
            I => \aluOperand1_0\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__35102\,
            I => \aluOperand1_0\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__35097\,
            I => \aluOperand1_0\
        );

    \I__7900\ : Odrv4
    port map (
            O => \N__35094\,
            I => \aluOperand1_0\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__35087\,
            I => \aluOperand1_0\
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__35072\,
            I => \ALU.aluOut_13_cascade_\
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__35069\,
            I => \N__35066\
        );

    \I__7896\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35062\
        );

    \I__7895\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35059\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__35054\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__35059\,
            I => \N__35054\
        );

    \I__7892\ : Odrv12
    port map (
            O => \N__35054\,
            I => \ALU.a13_b_0\
        );

    \I__7891\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35048\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__35045\
        );

    \I__7889\ : Span4Mux_h
    port map (
            O => \N__35045\,
            I => \N__35041\
        );

    \I__7888\ : InMux
    port map (
            O => \N__35044\,
            I => \N__35038\
        );

    \I__7887\ : Odrv4
    port map (
            O => \N__35041\,
            I => \ALU.fZ0Z_0\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__35038\,
            I => \ALU.fZ0Z_0\
        );

    \I__7885\ : InMux
    port map (
            O => \N__35033\,
            I => \N__35023\
        );

    \I__7884\ : InMux
    port map (
            O => \N__35032\,
            I => \N__35020\
        );

    \I__7883\ : InMux
    port map (
            O => \N__35031\,
            I => \N__35017\
        );

    \I__7882\ : InMux
    port map (
            O => \N__35030\,
            I => \N__35014\
        );

    \I__7881\ : InMux
    port map (
            O => \N__35029\,
            I => \N__35009\
        );

    \I__7880\ : InMux
    port map (
            O => \N__35028\,
            I => \N__35006\
        );

    \I__7879\ : InMux
    port map (
            O => \N__35027\,
            I => \N__35003\
        );

    \I__7878\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35000\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__34995\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__35020\,
            I => \N__34995\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N__34988\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34988\
        );

    \I__7873\ : InMux
    port map (
            O => \N__35013\,
            I => \N__34983\
        );

    \I__7872\ : InMux
    port map (
            O => \N__35012\,
            I => \N__34983\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__34980\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__35006\,
            I => \N__34977\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__35003\,
            I => \N__34972\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__35000\,
            I => \N__34972\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__34995\,
            I => \N__34969\
        );

    \I__7866\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34966\
        );

    \I__7865\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34963\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__34988\,
            I => \N__34960\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__34983\,
            I => \N__34957\
        );

    \I__7862\ : Span4Mux_h
    port map (
            O => \N__34980\,
            I => \N__34954\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__34977\,
            I => \N__34947\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__34972\,
            I => \N__34947\
        );

    \I__7859\ : Span4Mux_v
    port map (
            O => \N__34969\,
            I => \N__34947\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__34966\,
            I => \aluOperand2_1_rep1\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__34963\,
            I => \aluOperand2_1_rep1\
        );

    \I__7856\ : Odrv4
    port map (
            O => \N__34960\,
            I => \aluOperand2_1_rep1\
        );

    \I__7855\ : Odrv12
    port map (
            O => \N__34957\,
            I => \aluOperand2_1_rep1\
        );

    \I__7854\ : Odrv4
    port map (
            O => \N__34954\,
            I => \aluOperand2_1_rep1\
        );

    \I__7853\ : Odrv4
    port map (
            O => \N__34947\,
            I => \aluOperand2_1_rep1\
        );

    \I__7852\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34930\
        );

    \I__7851\ : InMux
    port map (
            O => \N__34933\,
            I => \N__34927\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34924\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34921\
        );

    \I__7848\ : Span4Mux_h
    port map (
            O => \N__34924\,
            I => \N__34918\
        );

    \I__7847\ : Span4Mux_h
    port map (
            O => \N__34921\,
            I => \N__34914\
        );

    \I__7846\ : Span4Mux_h
    port map (
            O => \N__34918\,
            I => \N__34911\
        );

    \I__7845\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34908\
        );

    \I__7844\ : Odrv4
    port map (
            O => \N__34914\,
            I => \ALU.cZ0Z_10\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__34911\,
            I => \ALU.cZ0Z_10\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__34908\,
            I => \ALU.cZ0Z_10\
        );

    \I__7841\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34898\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__34898\,
            I => \N__34895\
        );

    \I__7839\ : Span4Mux_v
    port map (
            O => \N__34895\,
            I => \N__34892\
        );

    \I__7838\ : Span4Mux_v
    port map (
            O => \N__34892\,
            I => \N__34888\
        );

    \I__7837\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34885\
        );

    \I__7836\ : Span4Mux_h
    port map (
            O => \N__34888\,
            I => \N__34877\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__34885\,
            I => \N__34877\
        );

    \I__7834\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34872\
        );

    \I__7833\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34872\
        );

    \I__7832\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34869\
        );

    \I__7831\ : Span4Mux_v
    port map (
            O => \N__34877\,
            I => \N__34864\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__34872\,
            I => \N__34859\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__34869\,
            I => \N__34856\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__34868\,
            I => \N__34851\
        );

    \I__7827\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34848\
        );

    \I__7826\ : Span4Mux_h
    port map (
            O => \N__34864\,
            I => \N__34845\
        );

    \I__7825\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34840\
        );

    \I__7824\ : InMux
    port map (
            O => \N__34862\,
            I => \N__34840\
        );

    \I__7823\ : Span4Mux_h
    port map (
            O => \N__34859\,
            I => \N__34837\
        );

    \I__7822\ : Span4Mux_h
    port map (
            O => \N__34856\,
            I => \N__34834\
        );

    \I__7821\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34827\
        );

    \I__7820\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34827\
        );

    \I__7819\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34827\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__34848\,
            I => \aluOperand2_fast_2\
        );

    \I__7817\ : Odrv4
    port map (
            O => \N__34845\,
            I => \aluOperand2_fast_2\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__34840\,
            I => \aluOperand2_fast_2\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__34837\,
            I => \aluOperand2_fast_2\
        );

    \I__7814\ : Odrv4
    port map (
            O => \N__34834\,
            I => \aluOperand2_fast_2\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__34827\,
            I => \aluOperand2_fast_2\
        );

    \I__7812\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34811\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__34811\,
            I => \N__34808\
        );

    \I__7810\ : Span4Mux_h
    port map (
            O => \N__34808\,
            I => \N__34805\
        );

    \I__7809\ : Span4Mux_h
    port map (
            O => \N__34805\,
            I => \N__34802\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__34802\,
            I => \ALU.g0_7_m4_1\
        );

    \I__7807\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34791\
        );

    \I__7806\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34788\
        );

    \I__7805\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34784\
        );

    \I__7804\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34777\
        );

    \I__7803\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34777\
        );

    \I__7802\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34777\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__34791\,
            I => \N__34774\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__34788\,
            I => \N__34771\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__34787\,
            I => \N__34766\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__34784\,
            I => \N__34759\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__34777\,
            I => \N__34759\
        );

    \I__7796\ : Span4Mux_v
    port map (
            O => \N__34774\,
            I => \N__34756\
        );

    \I__7795\ : Span4Mux_v
    port map (
            O => \N__34771\,
            I => \N__34753\
        );

    \I__7794\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34748\
        );

    \I__7793\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34748\
        );

    \I__7792\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34741\
        );

    \I__7791\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34741\
        );

    \I__7790\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34741\
        );

    \I__7789\ : Span4Mux_v
    port map (
            O => \N__34759\,
            I => \N__34738\
        );

    \I__7788\ : Sp12to4
    port map (
            O => \N__34756\,
            I => \N__34735\
        );

    \I__7787\ : Sp12to4
    port map (
            O => \N__34753\,
            I => \N__34732\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__34748\,
            I => \N_287_0\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__34741\,
            I => \N_287_0\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__34738\,
            I => \N_287_0\
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__34735\,
            I => \N_287_0\
        );

    \I__7782\ : Odrv12
    port map (
            O => \N__34732\,
            I => \N_287_0\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__34721\,
            I => \N__34717\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__34720\,
            I => \N__34711\
        );

    \I__7779\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34705\
        );

    \I__7778\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34698\
        );

    \I__7777\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34698\
        );

    \I__7776\ : InMux
    port map (
            O => \N__34714\,
            I => \N__34698\
        );

    \I__7775\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34695\
        );

    \I__7774\ : CEMux
    port map (
            O => \N__34710\,
            I => \N__34692\
        );

    \I__7773\ : CascadeMux
    port map (
            O => \N__34709\,
            I => \N__34688\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__34708\,
            I => \N__34682\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34678\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__34698\,
            I => \N__34675\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34672\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34669\
        );

    \I__7767\ : CEMux
    port map (
            O => \N__34691\,
            I => \N__34665\
        );

    \I__7766\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34662\
        );

    \I__7765\ : InMux
    port map (
            O => \N__34687\,
            I => \N__34657\
        );

    \I__7764\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34657\
        );

    \I__7763\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34652\
        );

    \I__7762\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34652\
        );

    \I__7761\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34649\
        );

    \I__7760\ : Span4Mux_h
    port map (
            O => \N__34678\,
            I => \N__34646\
        );

    \I__7759\ : Span4Mux_v
    port map (
            O => \N__34675\,
            I => \N__34643\
        );

    \I__7758\ : Span4Mux_h
    port map (
            O => \N__34672\,
            I => \N__34640\
        );

    \I__7757\ : Span4Mux_s3_h
    port map (
            O => \N__34669\,
            I => \N__34637\
        );

    \I__7756\ : InMux
    port map (
            O => \N__34668\,
            I => \N__34634\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__34665\,
            I => \N__34631\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__34662\,
            I => \N__34624\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__34657\,
            I => \N__34624\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__34652\,
            I => \N__34624\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34621\
        );

    \I__7750\ : Span4Mux_h
    port map (
            O => \N__34646\,
            I => \N__34618\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__34643\,
            I => \N__34613\
        );

    \I__7748\ : Span4Mux_h
    port map (
            O => \N__34640\,
            I => \N__34610\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__34637\,
            I => \N__34605\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__34634\,
            I => \N__34605\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__34631\,
            I => \N__34601\
        );

    \I__7744\ : Span12Mux_h
    port map (
            O => \N__34624\,
            I => \N__34594\
        );

    \I__7743\ : Sp12to4
    port map (
            O => \N__34621\,
            I => \N__34594\
        );

    \I__7742\ : Sp12to4
    port map (
            O => \N__34618\,
            I => \N__34594\
        );

    \I__7741\ : InMux
    port map (
            O => \N__34617\,
            I => \N__34589\
        );

    \I__7740\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34589\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__34613\,
            I => \N__34582\
        );

    \I__7738\ : Span4Mux_v
    port map (
            O => \N__34610\,
            I => \N__34582\
        );

    \I__7737\ : Span4Mux_s3_h
    port map (
            O => \N__34605\,
            I => \N__34582\
        );

    \I__7736\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34579\
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__34601\,
            I => \G_566\
        );

    \I__7734\ : Odrv12
    port map (
            O => \N__34594\,
            I => \G_566\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__34589\,
            I => \G_566\
        );

    \I__7732\ : Odrv4
    port map (
            O => \N__34582\,
            I => \G_566\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__34579\,
            I => \G_566\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__34568\,
            I => \N__34563\
        );

    \I__7729\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34558\
        );

    \I__7728\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34558\
        );

    \I__7727\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34555\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34552\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__34555\,
            I => \N__34549\
        );

    \I__7724\ : Span4Mux_v
    port map (
            O => \N__34552\,
            I => \N__34546\
        );

    \I__7723\ : Span4Mux_v
    port map (
            O => \N__34549\,
            I => \N__34542\
        );

    \I__7722\ : Sp12to4
    port map (
            O => \N__34546\,
            I => \N__34539\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__34545\,
            I => \N__34536\
        );

    \I__7720\ : Span4Mux_v
    port map (
            O => \N__34542\,
            I => \N__34533\
        );

    \I__7719\ : Span12Mux_h
    port map (
            O => \N__34539\,
            I => \N__34530\
        );

    \I__7718\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34527\
        );

    \I__7717\ : Sp12to4
    port map (
            O => \N__34533\,
            I => \N__34524\
        );

    \I__7716\ : Span12Mux_v
    port map (
            O => \N__34530\,
            I => \N__34521\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__34527\,
            I => \testWordZ0Z_11\
        );

    \I__7714\ : Odrv12
    port map (
            O => \N__34524\,
            I => \testWordZ0Z_11\
        );

    \I__7713\ : Odrv12
    port map (
            O => \N__34521\,
            I => \testWordZ0Z_11\
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__34514\,
            I => \N__34509\
        );

    \I__7711\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34505\
        );

    \I__7710\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34502\
        );

    \I__7709\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34497\
        );

    \I__7708\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34497\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34489\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__34502\,
            I => \N__34489\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__34497\,
            I => \N__34485\
        );

    \I__7704\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34482\
        );

    \I__7703\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34479\
        );

    \I__7702\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34476\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__34489\,
            I => \N__34470\
        );

    \I__7700\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34465\
        );

    \I__7699\ : Span4Mux_v
    port map (
            O => \N__34485\,
            I => \N__34462\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34459\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__34479\,
            I => \N__34454\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__34476\,
            I => \N__34454\
        );

    \I__7695\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34447\
        );

    \I__7694\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34447\
        );

    \I__7693\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34447\
        );

    \I__7692\ : Span4Mux_h
    port map (
            O => \N__34470\,
            I => \N__34444\
        );

    \I__7691\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34439\
        );

    \I__7690\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34439\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__34465\,
            I => \N__34434\
        );

    \I__7688\ : Span4Mux_h
    port map (
            O => \N__34462\,
            I => \N__34434\
        );

    \I__7687\ : Span4Mux_h
    port map (
            O => \N__34459\,
            I => \N__34431\
        );

    \I__7686\ : Span4Mux_h
    port map (
            O => \N__34454\,
            I => \N__34424\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__34447\,
            I => \N__34424\
        );

    \I__7684\ : Span4Mux_h
    port map (
            O => \N__34444\,
            I => \N__34424\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__34439\,
            I => \aluOperand2_1\
        );

    \I__7682\ : Odrv4
    port map (
            O => \N__34434\,
            I => \aluOperand2_1\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__34431\,
            I => \aluOperand2_1\
        );

    \I__7680\ : Odrv4
    port map (
            O => \N__34424\,
            I => \aluOperand2_1\
        );

    \I__7679\ : CascadeMux
    port map (
            O => \N__34415\,
            I => \N__34412\
        );

    \I__7678\ : InMux
    port map (
            O => \N__34412\,
            I => \N__34408\
        );

    \I__7677\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34405\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__34408\,
            I => \N__34399\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__34405\,
            I => \N__34396\
        );

    \I__7674\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34391\
        );

    \I__7673\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34388\
        );

    \I__7672\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34385\
        );

    \I__7671\ : Span4Mux_v
    port map (
            O => \N__34399\,
            I => \N__34381\
        );

    \I__7670\ : Span4Mux_h
    port map (
            O => \N__34396\,
            I => \N__34378\
        );

    \I__7669\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34375\
        );

    \I__7668\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34372\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34369\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__34388\,
            I => \N__34364\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__34385\,
            I => \N__34364\
        );

    \I__7664\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34361\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__34381\,
            I => \ALU.mult_10\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__34378\,
            I => \ALU.mult_10\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__34375\,
            I => \ALU.mult_10\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__34372\,
            I => \ALU.mult_10\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__34369\,
            I => \ALU.mult_10\
        );

    \I__7658\ : Odrv12
    port map (
            O => \N__34364\,
            I => \ALU.mult_10\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__34361\,
            I => \ALU.mult_10\
        );

    \I__7656\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34339\
        );

    \I__7655\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34336\
        );

    \I__7654\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34333\
        );

    \I__7653\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34330\
        );

    \I__7652\ : InMux
    port map (
            O => \N__34342\,
            I => \N__34327\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__34339\,
            I => \N__34317\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__34336\,
            I => \N__34317\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__34333\,
            I => \N__34317\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34317\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__34327\,
            I => \N__34314\
        );

    \I__7646\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34311\
        );

    \I__7645\ : Span4Mux_v
    port map (
            O => \N__34317\,
            I => \N__34307\
        );

    \I__7644\ : Span4Mux_v
    port map (
            O => \N__34314\,
            I => \N__34304\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__34311\,
            I => \N__34301\
        );

    \I__7642\ : InMux
    port map (
            O => \N__34310\,
            I => \N__34298\
        );

    \I__7641\ : Span4Mux_h
    port map (
            O => \N__34307\,
            I => \N__34295\
        );

    \I__7640\ : Sp12to4
    port map (
            O => \N__34304\,
            I => \N__34288\
        );

    \I__7639\ : Span12Mux_v
    port map (
            O => \N__34301\,
            I => \N__34288\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__34298\,
            I => \N__34288\
        );

    \I__7637\ : Odrv4
    port map (
            O => \N__34295\,
            I => \aluOperation_RNINNN4N3_0\
        );

    \I__7636\ : Odrv12
    port map (
            O => \N__34288\,
            I => \aluOperation_RNINNN4N3_0\
        );

    \I__7635\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34279\
        );

    \I__7634\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34276\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__34279\,
            I => \N__34273\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34270\
        );

    \I__7631\ : Span4Mux_v
    port map (
            O => \N__34273\,
            I => \N__34264\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__34270\,
            I => \N__34264\
        );

    \I__7629\ : CascadeMux
    port map (
            O => \N__34269\,
            I => \N__34261\
        );

    \I__7628\ : Span4Mux_h
    port map (
            O => \N__34264\,
            I => \N__34258\
        );

    \I__7627\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34255\
        );

    \I__7626\ : Odrv4
    port map (
            O => \N__34258\,
            I => \ALU.gZ0Z_10\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__34255\,
            I => \ALU.gZ0Z_10\
        );

    \I__7624\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34242\
        );

    \I__7623\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34239\
        );

    \I__7622\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34236\
        );

    \I__7621\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34233\
        );

    \I__7620\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34230\
        );

    \I__7619\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34227\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__34242\,
            I => \N__34224\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__34239\,
            I => \N__34215\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__34236\,
            I => \N__34215\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__34233\,
            I => \N__34215\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34215\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__34227\,
            I => \N__34211\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__34224\,
            I => \N__34208\
        );

    \I__7611\ : Span4Mux_v
    port map (
            O => \N__34215\,
            I => \N__34205\
        );

    \I__7610\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34202\
        );

    \I__7609\ : Span4Mux_h
    port map (
            O => \N__34211\,
            I => \N__34199\
        );

    \I__7608\ : Span4Mux_h
    port map (
            O => \N__34208\,
            I => \N__34196\
        );

    \I__7607\ : Sp12to4
    port map (
            O => \N__34205\,
            I => \N__34193\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__34202\,
            I => \N__34190\
        );

    \I__7605\ : Odrv4
    port map (
            O => \N__34199\,
            I => \aluOperation_RNI5QD2L3_0\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__34196\,
            I => \aluOperation_RNI5QD2L3_0\
        );

    \I__7603\ : Odrv12
    port map (
            O => \N__34193\,
            I => \aluOperation_RNI5QD2L3_0\
        );

    \I__7602\ : Odrv12
    port map (
            O => \N__34190\,
            I => \aluOperation_RNI5QD2L3_0\
        );

    \I__7601\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34176\
        );

    \I__7600\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34171\
        );

    \I__7599\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34168\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__34176\,
            I => \N__34164\
        );

    \I__7597\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34161\
        );

    \I__7596\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34157\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34154\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__34168\,
            I => \N__34151\
        );

    \I__7593\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34148\
        );

    \I__7592\ : Span4Mux_h
    port map (
            O => \N__34164\,
            I => \N__34144\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__34161\,
            I => \N__34141\
        );

    \I__7590\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34138\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__34157\,
            I => \N__34135\
        );

    \I__7588\ : Span4Mux_v
    port map (
            O => \N__34154\,
            I => \N__34128\
        );

    \I__7587\ : Span4Mux_h
    port map (
            O => \N__34151\,
            I => \N__34128\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__34148\,
            I => \N__34128\
        );

    \I__7585\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34125\
        );

    \I__7584\ : Odrv4
    port map (
            O => \N__34144\,
            I => \ALU.mult_11\
        );

    \I__7583\ : Odrv4
    port map (
            O => \N__34141\,
            I => \ALU.mult_11\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__34138\,
            I => \ALU.mult_11\
        );

    \I__7581\ : Odrv4
    port map (
            O => \N__34135\,
            I => \ALU.mult_11\
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__34128\,
            I => \ALU.mult_11\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__34125\,
            I => \ALU.mult_11\
        );

    \I__7578\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34109\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__34109\,
            I => \N__34106\
        );

    \I__7576\ : Span4Mux_v
    port map (
            O => \N__34106\,
            I => \N__34102\
        );

    \I__7575\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34099\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__34102\,
            I => \N__34094\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34094\
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__34094\,
            I => \ALU.gZ0Z_11\
        );

    \I__7571\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34083\
        );

    \I__7570\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34080\
        );

    \I__7569\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34077\
        );

    \I__7568\ : CascadeMux
    port map (
            O => \N__34088\,
            I => \N__34073\
        );

    \I__7567\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34070\
        );

    \I__7566\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34067\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__34064\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34059\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__34077\,
            I => \N__34059\
        );

    \I__7562\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34056\
        );

    \I__7561\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34053\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__34070\,
            I => \N__34048\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__34048\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__34064\,
            I => \N__34045\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__34059\,
            I => \N__34042\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__34056\,
            I => \aluOperation_RNIGPL5M3_0\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__34053\,
            I => \aluOperation_RNIGPL5M3_0\
        );

    \I__7554\ : Odrv4
    port map (
            O => \N__34048\,
            I => \aluOperation_RNIGPL5M3_0\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__34045\,
            I => \aluOperation_RNIGPL5M3_0\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__34042\,
            I => \aluOperation_RNIGPL5M3_0\
        );

    \I__7551\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34027\
        );

    \I__7550\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34022\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__34017\
        );

    \I__7548\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34014\
        );

    \I__7547\ : InMux
    port map (
            O => \N__34025\,
            I => \N__34011\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__34022\,
            I => \N__34007\
        );

    \I__7545\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34004\
        );

    \I__7544\ : InMux
    port map (
            O => \N__34020\,
            I => \N__34001\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__34017\,
            I => \N__33997\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__34014\,
            I => \N__33994\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__34011\,
            I => \N__33991\
        );

    \I__7540\ : InMux
    port map (
            O => \N__34010\,
            I => \N__33988\
        );

    \I__7539\ : Span4Mux_v
    port map (
            O => \N__34007\,
            I => \N__33983\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__34004\,
            I => \N__33983\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__34001\,
            I => \N__33980\
        );

    \I__7536\ : InMux
    port map (
            O => \N__34000\,
            I => \N__33977\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__33997\,
            I => \ALU.mult_12\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__33994\,
            I => \ALU.mult_12\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__33991\,
            I => \ALU.mult_12\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__33988\,
            I => \ALU.mult_12\
        );

    \I__7531\ : Odrv4
    port map (
            O => \N__33983\,
            I => \ALU.mult_12\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__33980\,
            I => \ALU.mult_12\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__33977\,
            I => \ALU.mult_12\
        );

    \I__7528\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33959\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__33959\,
            I => \N__33955\
        );

    \I__7526\ : InMux
    port map (
            O => \N__33958\,
            I => \N__33952\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__33955\,
            I => \N__33947\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__33952\,
            I => \N__33947\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__33947\,
            I => \N__33944\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__33944\,
            I => \ALU.gZ0Z_12\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__33941\,
            I => \N__33936\
        );

    \I__7520\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33931\
        );

    \I__7519\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33928\
        );

    \I__7518\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33925\
        );

    \I__7517\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33922\
        );

    \I__7516\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33917\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__33931\,
            I => \N__33914\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__33928\,
            I => \N__33911\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33906\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__33922\,
            I => \N__33906\
        );

    \I__7511\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33903\
        );

    \I__7510\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33900\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__33917\,
            I => \N__33895\
        );

    \I__7508\ : Span4Mux_h
    port map (
            O => \N__33914\,
            I => \N__33895\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__33911\,
            I => \N__33890\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__33906\,
            I => \N__33890\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__33903\,
            I => \aluOperation_RNI2J9SL3_0\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__33900\,
            I => \aluOperation_RNI2J9SL3_0\
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__33895\,
            I => \aluOperation_RNI2J9SL3_0\
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__33890\,
            I => \aluOperation_RNI2J9SL3_0\
        );

    \I__7501\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33877\
        );

    \I__7500\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33874\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33868\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33865\
        );

    \I__7497\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33860\
        );

    \I__7496\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33857\
        );

    \I__7495\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33854\
        );

    \I__7494\ : Span4Mux_h
    port map (
            O => \N__33868\,
            I => \N__33848\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__33865\,
            I => \N__33848\
        );

    \I__7492\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33845\
        );

    \I__7491\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33842\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33839\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__33857\,
            I => \N__33834\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__33854\,
            I => \N__33834\
        );

    \I__7487\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33831\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__33848\,
            I => \ALU.mult_13\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__33845\,
            I => \ALU.mult_13\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__33842\,
            I => \ALU.mult_13\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__33839\,
            I => \ALU.mult_13\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__33834\,
            I => \ALU.mult_13\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__33831\,
            I => \ALU.mult_13\
        );

    \I__7480\ : InMux
    port map (
            O => \N__33818\,
            I => \N__33809\
        );

    \I__7479\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33806\
        );

    \I__7478\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33803\
        );

    \I__7477\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33800\
        );

    \I__7476\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33797\
        );

    \I__7475\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33794\
        );

    \I__7474\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33791\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__33809\,
            I => \N__33788\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__33806\,
            I => \N__33785\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33782\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__33800\,
            I => \N__33769\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__33797\,
            I => \N__33769\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__33794\,
            I => \N__33769\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33769\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__33788\,
            I => \N__33769\
        );

    \I__7465\ : Span4Mux_v
    port map (
            O => \N__33785\,
            I => \N__33769\
        );

    \I__7464\ : Span4Mux_h
    port map (
            O => \N__33782\,
            I => \N__33766\
        );

    \I__7463\ : Span4Mux_v
    port map (
            O => \N__33769\,
            I => \N__33763\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__33766\,
            I => \aluOperation_RNIR872K3_0\
        );

    \I__7461\ : Odrv4
    port map (
            O => \N__33763\,
            I => \aluOperation_RNIR872K3_0\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33758\,
            I => \N__33753\
        );

    \I__7459\ : InMux
    port map (
            O => \N__33757\,
            I => \N__33750\
        );

    \I__7458\ : InMux
    port map (
            O => \N__33756\,
            I => \N__33744\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__33753\,
            I => \N__33741\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__33750\,
            I => \N__33737\
        );

    \I__7455\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33734\
        );

    \I__7454\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33731\
        );

    \I__7453\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33728\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33724\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__33741\,
            I => \N__33721\
        );

    \I__7450\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33718\
        );

    \I__7449\ : Span4Mux_h
    port map (
            O => \N__33737\,
            I => \N__33713\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__33734\,
            I => \N__33713\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__33731\,
            I => \N__33708\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__33728\,
            I => \N__33708\
        );

    \I__7445\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33705\
        );

    \I__7444\ : Odrv4
    port map (
            O => \N__33724\,
            I => \ALU.mult_14\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__33721\,
            I => \ALU.mult_14\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__33718\,
            I => \ALU.mult_14\
        );

    \I__7441\ : Odrv4
    port map (
            O => \N__33713\,
            I => \ALU.mult_14\
        );

    \I__7440\ : Odrv4
    port map (
            O => \N__33708\,
            I => \ALU.mult_14\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__33705\,
            I => \ALU.mult_14\
        );

    \I__7438\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33689\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33686\
        );

    \I__7436\ : Span4Mux_h
    port map (
            O => \N__33686\,
            I => \N__33682\
        );

    \I__7435\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33679\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__33682\,
            I => \N__33676\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__33679\,
            I => \N__33673\
        );

    \I__7432\ : Span4Mux_h
    port map (
            O => \N__33676\,
            I => \N__33670\
        );

    \I__7431\ : Span12Mux_s11_h
    port map (
            O => \N__33673\,
            I => \N__33667\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__33670\,
            I => \ALU.gZ0Z_14\
        );

    \I__7429\ : Odrv12
    port map (
            O => \N__33667\,
            I => \ALU.gZ0Z_14\
        );

    \I__7428\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33656\
        );

    \I__7427\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33650\
        );

    \I__7426\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33647\
        );

    \I__7425\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33644\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__33656\,
            I => \N__33641\
        );

    \I__7423\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33638\
        );

    \I__7422\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33635\
        );

    \I__7421\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33632\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33623\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__33647\,
            I => \N__33623\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__33644\,
            I => \N__33623\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__33641\,
            I => \N__33623\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33620\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__33635\,
            I => \N__33615\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__33632\,
            I => \N__33615\
        );

    \I__7413\ : Span4Mux_v
    port map (
            O => \N__33623\,
            I => \N__33612\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__33620\,
            I => \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93\
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__33615\,
            I => \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93\
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__33612\,
            I => \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93\
        );

    \I__7409\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33598\
        );

    \I__7408\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33595\
        );

    \I__7407\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33592\
        );

    \I__7406\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33586\
        );

    \I__7405\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33583\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__33598\,
            I => \N__33580\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__33595\,
            I => \N__33577\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__33592\,
            I => \N__33574\
        );

    \I__7401\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33571\
        );

    \I__7400\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33568\
        );

    \I__7399\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33565\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33562\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__33583\,
            I => \N__33557\
        );

    \I__7396\ : Span4Mux_h
    port map (
            O => \N__33580\,
            I => \N__33557\
        );

    \I__7395\ : Span4Mux_h
    port map (
            O => \N__33577\,
            I => \N__33552\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__33574\,
            I => \N__33552\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__33571\,
            I => \ALU.mult_15\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__33568\,
            I => \ALU.mult_15\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__33565\,
            I => \ALU.mult_15\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__33562\,
            I => \ALU.mult_15\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__33557\,
            I => \ALU.mult_15\
        );

    \I__7388\ : Odrv4
    port map (
            O => \N__33552\,
            I => \ALU.mult_15\
        );

    \I__7387\ : InMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__33536\,
            I => \N__33532\
        );

    \I__7385\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33529\
        );

    \I__7384\ : Span4Mux_v
    port map (
            O => \N__33532\,
            I => \N__33526\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__33529\,
            I => \ALU.gZ0Z_15\
        );

    \I__7382\ : Odrv4
    port map (
            O => \N__33526\,
            I => \ALU.gZ0Z_15\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__33521\,
            I => \ALU.a_15_m4_15_cascade_\
        );

    \I__7380\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33515\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__33515\,
            I => \N__33512\
        );

    \I__7378\ : Span4Mux_v
    port map (
            O => \N__33512\,
            I => \N__33509\
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__33509\,
            I => \ALU.a_15_m3_15\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__33506\,
            I => \ALU.c_RNIR4QHM2Z0Z_15_cascade_\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__33503\,
            I => \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93_cascade_\
        );

    \I__7374\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33497\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__33497\,
            I => \N__33494\
        );

    \I__7372\ : Span4Mux_h
    port map (
            O => \N__33494\,
            I => \N__33491\
        );

    \I__7371\ : Span4Mux_h
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__7370\ : Span4Mux_v
    port map (
            O => \N__33488\,
            I => \N__33484\
        );

    \I__7369\ : InMux
    port map (
            O => \N__33487\,
            I => \N__33481\
        );

    \I__7368\ : Odrv4
    port map (
            O => \N__33484\,
            I => \ALU.hZ0Z_15\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__33481\,
            I => \ALU.hZ0Z_15\
        );

    \I__7366\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33473\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__33473\,
            I => \N__33469\
        );

    \I__7364\ : InMux
    port map (
            O => \N__33472\,
            I => \N__33466\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__33469\,
            I => \N__33463\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33460\
        );

    \I__7361\ : Span4Mux_v
    port map (
            O => \N__33463\,
            I => \N__33457\
        );

    \I__7360\ : Span4Mux_v
    port map (
            O => \N__33460\,
            I => \N__33454\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__33457\,
            I => \ALU.dZ0Z_15\
        );

    \I__7358\ : Odrv4
    port map (
            O => \N__33454\,
            I => \ALU.dZ0Z_15\
        );

    \I__7357\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__33446\,
            I => \ALU.d_RNISBLUZ0Z_15\
        );

    \I__7355\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33439\
        );

    \I__7354\ : CEMux
    port map (
            O => \N__33442\,
            I => \N__33435\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__33439\,
            I => \N__33431\
        );

    \I__7352\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33428\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__33435\,
            I => \N__33425\
        );

    \I__7350\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33422\
        );

    \I__7349\ : Sp12to4
    port map (
            O => \N__33431\,
            I => \N__33419\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__33428\,
            I => \N__33416\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__33425\,
            I => \N__33411\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33411\
        );

    \I__7345\ : Span12Mux_v
    port map (
            O => \N__33419\,
            I => \N__33408\
        );

    \I__7344\ : Span12Mux_s4_v
    port map (
            O => \N__33416\,
            I => \N__33405\
        );

    \I__7343\ : Span4Mux_s0_v
    port map (
            O => \N__33411\,
            I => \N__33402\
        );

    \I__7342\ : Odrv12
    port map (
            O => \N__33408\,
            I => \CONTROL.aluOperation_cnvZ0Z_0\
        );

    \I__7341\ : Odrv12
    port map (
            O => \N__33405\,
            I => \CONTROL.aluOperation_cnvZ0Z_0\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__33402\,
            I => \CONTROL.aluOperation_cnvZ0Z_0\
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__7338\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33389\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__33389\,
            I => \N__33386\
        );

    \I__7336\ : Span4Mux_h
    port map (
            O => \N__33386\,
            I => \N__33381\
        );

    \I__7335\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33376\
        );

    \I__7334\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33376\
        );

    \I__7333\ : Span4Mux_h
    port map (
            O => \N__33381\,
            I => \N__33373\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__33376\,
            I => \N__33370\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__33373\,
            I => \N__33367\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__33370\,
            I => \N__33362\
        );

    \I__7329\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33362\
        );

    \I__7328\ : Odrv4
    port map (
            O => \N__33362\,
            I => \N_723\
        );

    \I__7327\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33351\
        );

    \I__7326\ : InMux
    port map (
            O => \N__33358\,
            I => \N__33342\
        );

    \I__7325\ : InMux
    port map (
            O => \N__33357\,
            I => \N__33342\
        );

    \I__7324\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33342\
        );

    \I__7323\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33342\
        );

    \I__7322\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33339\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__33351\,
            I => \N__33336\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__33342\,
            I => \N__33332\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__33339\,
            I => \N__33325\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__33336\,
            I => \N__33325\
        );

    \I__7317\ : CascadeMux
    port map (
            O => \N__33335\,
            I => \N__33322\
        );

    \I__7316\ : Span4Mux_h
    port map (
            O => \N__33332\,
            I => \N__33319\
        );

    \I__7315\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33313\
        );

    \I__7314\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33310\
        );

    \I__7313\ : Span4Mux_h
    port map (
            O => \N__33325\,
            I => \N__33307\
        );

    \I__7312\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33304\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__33319\,
            I => \N__33297\
        );

    \I__7310\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33287\
        );

    \I__7309\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33287\
        );

    \I__7308\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33287\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33282\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__33310\,
            I => \N__33282\
        );

    \I__7305\ : Span4Mux_h
    port map (
            O => \N__33307\,
            I => \N__33279\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__33304\,
            I => \N__33276\
        );

    \I__7303\ : CascadeMux
    port map (
            O => \N__33303\,
            I => \N__33272\
        );

    \I__7302\ : CascadeMux
    port map (
            O => \N__33302\,
            I => \N__33268\
        );

    \I__7301\ : CascadeMux
    port map (
            O => \N__33301\,
            I => \N__33265\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__33300\,
            I => \N__33256\
        );

    \I__7299\ : IoSpan4Mux
    port map (
            O => \N__33297\,
            I => \N__33253\
        );

    \I__7298\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33246\
        );

    \I__7297\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33246\
        );

    \I__7296\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33246\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__33287\,
            I => \N__33240\
        );

    \I__7294\ : Span4Mux_v
    port map (
            O => \N__33282\,
            I => \N__33240\
        );

    \I__7293\ : Span4Mux_h
    port map (
            O => \N__33279\,
            I => \N__33237\
        );

    \I__7292\ : Span4Mux_h
    port map (
            O => \N__33276\,
            I => \N__33234\
        );

    \I__7291\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33227\
        );

    \I__7290\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33227\
        );

    \I__7289\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33227\
        );

    \I__7288\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33220\
        );

    \I__7287\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33220\
        );

    \I__7286\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33220\
        );

    \I__7285\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33213\
        );

    \I__7284\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33213\
        );

    \I__7283\ : InMux
    port map (
            O => \N__33261\,
            I => \N__33213\
        );

    \I__7282\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33210\
        );

    \I__7281\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33205\
        );

    \I__7280\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33205\
        );

    \I__7279\ : Span4Mux_s0_v
    port map (
            O => \N__33253\,
            I => \N__33200\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33200\
        );

    \I__7277\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33197\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__33240\,
            I => \N__33192\
        );

    \I__7275\ : Span4Mux_v
    port map (
            O => \N__33237\,
            I => \N__33192\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__33234\,
            I => \testWordZ0Z_5\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__33227\,
            I => \testWordZ0Z_5\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__33220\,
            I => \testWordZ0Z_5\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__33213\,
            I => \testWordZ0Z_5\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__33210\,
            I => \testWordZ0Z_5\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__33205\,
            I => \testWordZ0Z_5\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__33200\,
            I => \testWordZ0Z_5\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__33197\,
            I => \testWordZ0Z_5\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__33192\,
            I => \testWordZ0Z_5\
        );

    \I__7265\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__33170\,
            I => \N__33167\
        );

    \I__7263\ : Span4Mux_h
    port map (
            O => \N__33167\,
            I => \N__33164\
        );

    \I__7262\ : Span4Mux_h
    port map (
            O => \N__33164\,
            I => \N__33160\
        );

    \I__7261\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33157\
        );

    \I__7260\ : Span4Mux_v
    port map (
            O => \N__33160\,
            I => \N__33154\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__33157\,
            I => \aluOperation_5\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__33154\,
            I => \aluOperation_5\
        );

    \I__7257\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33145\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__33148\,
            I => \N__33142\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33139\
        );

    \I__7254\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33136\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__33139\,
            I => \N__33133\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__33136\,
            I => \N__33130\
        );

    \I__7251\ : Span4Mux_v
    port map (
            O => \N__33133\,
            I => \N__33127\
        );

    \I__7250\ : Span4Mux_h
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__7249\ : Span4Mux_h
    port map (
            O => \N__33127\,
            I => \N__33121\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__33124\,
            I => \N__33118\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__33121\,
            I => \ALU.a2_b_0\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__33118\,
            I => \ALU.a2_b_0\
        );

    \I__7245\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33110\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__33110\,
            I => \N__33107\
        );

    \I__7243\ : Odrv12
    port map (
            O => \N__33107\,
            I => \ALU.madd_axb_1_l_ofx\
        );

    \I__7242\ : CascadeMux
    port map (
            O => \N__33104\,
            I => \N__33100\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__33103\,
            I => \N__33097\
        );

    \I__7240\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33093\
        );

    \I__7239\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33090\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__33096\,
            I => \N__33086\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__33093\,
            I => \N__33081\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__33090\,
            I => \N__33078\
        );

    \I__7235\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33075\
        );

    \I__7234\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33072\
        );

    \I__7233\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33069\
        );

    \I__7232\ : InMux
    port map (
            O => \N__33084\,
            I => \N__33066\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__33081\,
            I => \N__33055\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__33078\,
            I => \N__33055\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__33075\,
            I => \N__33055\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33052\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33049\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__33066\,
            I => \N__33045\
        );

    \I__7225\ : InMux
    port map (
            O => \N__33065\,
            I => \N__33042\
        );

    \I__7224\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33037\
        );

    \I__7223\ : InMux
    port map (
            O => \N__33063\,
            I => \N__33037\
        );

    \I__7222\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33034\
        );

    \I__7221\ : Span4Mux_h
    port map (
            O => \N__33055\,
            I => \N__33031\
        );

    \I__7220\ : Sp12to4
    port map (
            O => \N__33052\,
            I => \N__33026\
        );

    \I__7219\ : Sp12to4
    port map (
            O => \N__33049\,
            I => \N__33026\
        );

    \I__7218\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33023\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__33045\,
            I => \N__33020\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__33042\,
            I => \N__33013\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__33037\,
            I => \N__33013\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__33034\,
            I => \N__33013\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__33031\,
            I => \N__33010\
        );

    \I__7212\ : Span12Mux_v
    port map (
            O => \N__33026\,
            I => \N__33007\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__33023\,
            I => \aluOperand2_0_rep2\
        );

    \I__7210\ : Odrv4
    port map (
            O => \N__33020\,
            I => \aluOperand2_0_rep2\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__33013\,
            I => \aluOperand2_0_rep2\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__33010\,
            I => \aluOperand2_0_rep2\
        );

    \I__7207\ : Odrv12
    port map (
            O => \N__33007\,
            I => \aluOperand2_0_rep2\
        );

    \I__7206\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32987\
        );

    \I__7205\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32984\
        );

    \I__7204\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32980\
        );

    \I__7203\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32975\
        );

    \I__7202\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32975\
        );

    \I__7201\ : InMux
    port map (
            O => \N__32991\,
            I => \N__32972\
        );

    \I__7200\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32967\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__32987\,
            I => \N__32964\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__32984\,
            I => \N__32960\
        );

    \I__7197\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32956\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__32980\,
            I => \N__32953\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32950\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32972\,
            I => \N__32947\
        );

    \I__7193\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32943\
        );

    \I__7192\ : InMux
    port map (
            O => \N__32970\,
            I => \N__32940\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__32967\,
            I => \N__32935\
        );

    \I__7190\ : Span4Mux_s3_h
    port map (
            O => \N__32964\,
            I => \N__32935\
        );

    \I__7189\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32932\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__32960\,
            I => \N__32929\
        );

    \I__7187\ : CascadeMux
    port map (
            O => \N__32959\,
            I => \N__32926\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32921\
        );

    \I__7185\ : Span4Mux_h
    port map (
            O => \N__32953\,
            I => \N__32921\
        );

    \I__7184\ : Span4Mux_v
    port map (
            O => \N__32950\,
            I => \N__32918\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__32947\,
            I => \N__32915\
        );

    \I__7182\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32912\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__32943\,
            I => \N__32909\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__32940\,
            I => \N__32906\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__32935\,
            I => \N__32903\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32899\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__32929\,
            I => \N__32896\
        );

    \I__7176\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32893\
        );

    \I__7175\ : Span4Mux_h
    port map (
            O => \N__32921\,
            I => \N__32890\
        );

    \I__7174\ : Span4Mux_h
    port map (
            O => \N__32918\,
            I => \N__32885\
        );

    \I__7173\ : Span4Mux_h
    port map (
            O => \N__32915\,
            I => \N__32885\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32876\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__32909\,
            I => \N__32876\
        );

    \I__7170\ : Span4Mux_h
    port map (
            O => \N__32906\,
            I => \N__32876\
        );

    \I__7169\ : Span4Mux_h
    port map (
            O => \N__32903\,
            I => \N__32876\
        );

    \I__7168\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32873\
        );

    \I__7167\ : Span12Mux_v
    port map (
            O => \N__32899\,
            I => \N__32870\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__32896\,
            I => \N__32867\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__32893\,
            I => \aluOperand2_0\
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__32890\,
            I => \aluOperand2_0\
        );

    \I__7163\ : Odrv4
    port map (
            O => \N__32885\,
            I => \aluOperand2_0\
        );

    \I__7162\ : Odrv4
    port map (
            O => \N__32876\,
            I => \aluOperand2_0\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__32873\,
            I => \aluOperand2_0\
        );

    \I__7160\ : Odrv12
    port map (
            O => \N__32870\,
            I => \aluOperand2_0\
        );

    \I__7159\ : Odrv4
    port map (
            O => \N__32867\,
            I => \aluOperand2_0\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__32852\,
            I => \ALU.g_RNIVGLLZ0Z_9_cascade_\
        );

    \I__7157\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__32846\,
            I => \N__32843\
        );

    \I__7155\ : Odrv12
    port map (
            O => \N__32843\,
            I => \ALU.operand2_7_ns_1_9\
        );

    \I__7154\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32836\
        );

    \I__7153\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32833\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32830\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__32833\,
            I => \N__32827\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__32830\,
            I => \N__32824\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__32827\,
            I => \N__32821\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__32824\,
            I => \N__32818\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__32821\,
            I => \N__32814\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__32818\,
            I => \N__32811\
        );

    \I__7145\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32808\
        );

    \I__7144\ : Span4Mux_h
    port map (
            O => \N__32814\,
            I => \N__32805\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__32811\,
            I => \ALU.hZ0Z_9\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__32808\,
            I => \ALU.hZ0Z_9\
        );

    \I__7141\ : Odrv4
    port map (
            O => \N__32805\,
            I => \ALU.hZ0Z_9\
        );

    \I__7140\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32793\
        );

    \I__7139\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32790\
        );

    \I__7138\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32787\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__32793\,
            I => \N__32784\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32781\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32778\
        );

    \I__7134\ : Span4Mux_v
    port map (
            O => \N__32784\,
            I => \N__32775\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__32781\,
            I => \N__32772\
        );

    \I__7132\ : Span4Mux_v
    port map (
            O => \N__32778\,
            I => \N__32767\
        );

    \I__7131\ : Span4Mux_v
    port map (
            O => \N__32775\,
            I => \N__32767\
        );

    \I__7130\ : Span4Mux_h
    port map (
            O => \N__32772\,
            I => \N__32764\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__32767\,
            I => \ALU.dZ0Z_9\
        );

    \I__7128\ : Odrv4
    port map (
            O => \N__32764\,
            I => \ALU.dZ0Z_9\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__7126\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32753\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__7124\ : Span4Mux_h
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__7123\ : Span4Mux_h
    port map (
            O => \N__32747\,
            I => \N__32744\
        );

    \I__7122\ : Odrv4
    port map (
            O => \N__32744\,
            I => \ALU.g0_0_0_m2_1\
        );

    \I__7121\ : CascadeMux
    port map (
            O => \N__32741\,
            I => \ALU.N_11_cascade_\
        );

    \I__7120\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__7118\ : Span4Mux_s3_h
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__32726\,
            I => \N__32723\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__32723\,
            I => \ALU.N_13\
        );

    \I__7114\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32717\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__32717\,
            I => \N__32712\
        );

    \I__7112\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32707\
        );

    \I__7111\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32707\
        );

    \I__7110\ : Span4Mux_h
    port map (
            O => \N__32712\,
            I => \N__32704\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__32707\,
            I => \N__32701\
        );

    \I__7108\ : Span4Mux_h
    port map (
            O => \N__32704\,
            I => \N__32696\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__32701\,
            I => \N__32696\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__32696\,
            I => \ALU.cZ0Z_9\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__7104\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__32687\,
            I => \ALU.g0_0_0_m2_0_1\
        );

    \I__7102\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32678\
        );

    \I__7100\ : Odrv4
    port map (
            O => \N__32678\,
            I => \ALU.N_12\
        );

    \I__7099\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32671\
        );

    \I__7098\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32667\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__32671\,
            I => \N__32662\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__32670\,
            I => \N__32658\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32655\
        );

    \I__7094\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32652\
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__32665\,
            I => \N__32649\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__32662\,
            I => \N__32646\
        );

    \I__7091\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32641\
        );

    \I__7090\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32641\
        );

    \I__7089\ : Span12Mux_h
    port map (
            O => \N__32655\,
            I => \N__32638\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__32652\,
            I => \N__32635\
        );

    \I__7087\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32632\
        );

    \I__7086\ : Span4Mux_v
    port map (
            O => \N__32646\,
            I => \N__32627\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32627\
        );

    \I__7084\ : Odrv12
    port map (
            O => \N__32638\,
            I => \ALU.aluOut_15\
        );

    \I__7083\ : Odrv12
    port map (
            O => \N__32635\,
            I => \ALU.aluOut_15\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__32632\,
            I => \ALU.aluOut_15\
        );

    \I__7081\ : Odrv4
    port map (
            O => \N__32627\,
            I => \ALU.aluOut_15\
        );

    \I__7080\ : CascadeMux
    port map (
            O => \N__32618\,
            I => \ALU.a_15_m2_ns_1Z0Z_15_cascade_\
        );

    \I__7079\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32612\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__32612\,
            I => \N__32609\
        );

    \I__7077\ : Span4Mux_h
    port map (
            O => \N__32609\,
            I => \N__32605\
        );

    \I__7076\ : InMux
    port map (
            O => \N__32608\,
            I => \N__32601\
        );

    \I__7075\ : Span4Mux_h
    port map (
            O => \N__32605\,
            I => \N__32598\
        );

    \I__7074\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32595\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__32601\,
            I => \N__32592\
        );

    \I__7072\ : Odrv4
    port map (
            O => \N__32598\,
            I => \ALU.N_7_0\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__32595\,
            I => \ALU.N_7_0\
        );

    \I__7070\ : Odrv12
    port map (
            O => \N__32592\,
            I => \ALU.N_7_0\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__32585\,
            I => \ALU.a_15_m2_15_cascade_\
        );

    \I__7068\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32579\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__32579\,
            I => \N__32576\
        );

    \I__7066\ : Span4Mux_h
    port map (
            O => \N__32576\,
            I => \N__32573\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__32573\,
            I => \N__32570\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__32570\,
            I => \ALU.lshift_15\
        );

    \I__7063\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32564\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__32564\,
            I => \N__32561\
        );

    \I__7061\ : Odrv12
    port map (
            O => \N__32561\,
            I => \TXbufferZ0Z_7\
        );

    \I__7060\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32555\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__32555\,
            I => \FTDI.TXshiftZ0Z_7\
        );

    \I__7058\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32546\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__32546\,
            I => \N__32543\
        );

    \I__7055\ : Span4Mux_h
    port map (
            O => \N__32543\,
            I => \N__32540\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__32540\,
            I => \ALU.un2_addsub_cry_10_c_RNIUS1OJZ0\
        );

    \I__7053\ : CascadeMux
    port map (
            O => \N__32537\,
            I => \ALU.a_15_m2_ns_1Z0Z_11_cascade_\
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__32534\,
            I => \ALU.a_15_m2_11_cascade_\
        );

    \I__7051\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32528\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__32525\,
            I => \N__32522\
        );

    \I__7048\ : Span4Mux_h
    port map (
            O => \N__32522\,
            I => \N__32519\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__32519\,
            I => \ALU.lshift_11\
        );

    \I__7046\ : CascadeMux
    port map (
            O => \N__32516\,
            I => \ALU.a_15_m4_11_cascade_\
        );

    \I__7045\ : InMux
    port map (
            O => \N__32513\,
            I => \N__32510\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32507\
        );

    \I__7043\ : Span4Mux_h
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__7042\ : Odrv4
    port map (
            O => \N__32504\,
            I => \ALU.a_15_m3_11\
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__32501\,
            I => \c_RNID7K8N2_11_cascade_\
        );

    \I__7040\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32495\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__32495\,
            I => \un2_addsub_cry_10_c_RNIEBKOT\
        );

    \I__7038\ : CascadeMux
    port map (
            O => \N__32492\,
            I => \aluOperation_RNI5QD2L3_0_cascade_\
        );

    \I__7037\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32486\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__32486\,
            I => \N__32483\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__32483\,
            I => \N__32479\
        );

    \I__7034\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32476\
        );

    \I__7033\ : Span4Mux_h
    port map (
            O => \N__32479\,
            I => \N__32471\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__32476\,
            I => \N__32471\
        );

    \I__7031\ : Odrv4
    port map (
            O => \N__32471\,
            I => \ALU.aZ0Z_11\
        );

    \I__7030\ : CEMux
    port map (
            O => \N__32468\,
            I => \N__32464\
        );

    \I__7029\ : CEMux
    port map (
            O => \N__32467\,
            I => \N__32461\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__32464\,
            I => \N__32458\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32454\
        );

    \I__7026\ : Span4Mux_v
    port map (
            O => \N__32458\,
            I => \N__32451\
        );

    \I__7025\ : CEMux
    port map (
            O => \N__32457\,
            I => \N__32448\
        );

    \I__7024\ : Span4Mux_v
    port map (
            O => \N__32454\,
            I => \N__32445\
        );

    \I__7023\ : Span4Mux_v
    port map (
            O => \N__32451\,
            I => \N__32439\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32439\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__32445\,
            I => \N__32436\
        );

    \I__7020\ : CEMux
    port map (
            O => \N__32444\,
            I => \N__32432\
        );

    \I__7019\ : Span4Mux_h
    port map (
            O => \N__32439\,
            I => \N__32429\
        );

    \I__7018\ : Span4Mux_v
    port map (
            O => \N__32436\,
            I => \N__32426\
        );

    \I__7017\ : CEMux
    port map (
            O => \N__32435\,
            I => \N__32423\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__32432\,
            I => \N__32420\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__32429\,
            I => \N__32417\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__32426\,
            I => \N__32414\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32411\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__32420\,
            I => \N__32408\
        );

    \I__7011\ : Span4Mux_v
    port map (
            O => \N__32417\,
            I => \N__32405\
        );

    \I__7010\ : IoSpan4Mux
    port map (
            O => \N__32414\,
            I => \N__32402\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__32411\,
            I => \N__32399\
        );

    \I__7008\ : Sp12to4
    port map (
            O => \N__32408\,
            I => \N__32396\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__32405\,
            I => \N__32393\
        );

    \I__7006\ : Span4Mux_s1_v
    port map (
            O => \N__32402\,
            I => \N__32390\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__32399\,
            I => \N__32387\
        );

    \I__7004\ : Span12Mux_s10_h
    port map (
            O => \N__32396\,
            I => \N__32384\
        );

    \I__7003\ : Span4Mux_h
    port map (
            O => \N__32393\,
            I => \N__32379\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__32390\,
            I => \N__32379\
        );

    \I__7001\ : Span4Mux_h
    port map (
            O => \N__32387\,
            I => \N__32376\
        );

    \I__7000\ : Span12Mux_v
    port map (
            O => \N__32384\,
            I => \N__32373\
        );

    \I__6999\ : Span4Mux_h
    port map (
            O => \N__32379\,
            I => \N__32370\
        );

    \I__6998\ : Odrv4
    port map (
            O => \N__32376\,
            I => \ALU.e_cnvZ0Z_0\
        );

    \I__6997\ : Odrv12
    port map (
            O => \N__32373\,
            I => \ALU.e_cnvZ0Z_0\
        );

    \I__6996\ : Odrv4
    port map (
            O => \N__32370\,
            I => \ALU.e_cnvZ0Z_0\
        );

    \I__6995\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32359\
        );

    \I__6994\ : IoInMux
    port map (
            O => \N__32362\,
            I => \N__32356\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__32359\,
            I => \N__32353\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__32356\,
            I => \N__32350\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__32353\,
            I => \N__32347\
        );

    \I__6990\ : Span4Mux_s3_v
    port map (
            O => \N__32350\,
            I => \N__32344\
        );

    \I__6989\ : Sp12to4
    port map (
            O => \N__32347\,
            I => \N__32341\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__32344\,
            I => \N__32338\
        );

    \I__6987\ : Span12Mux_s10_v
    port map (
            O => \N__32341\,
            I => \N__32335\
        );

    \I__6986\ : Sp12to4
    port map (
            O => \N__32338\,
            I => \N__32332\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__32335\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6984\ : Odrv12
    port map (
            O => \N__32332\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__32327\,
            I => \N__32323\
        );

    \I__6982\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32316\
        );

    \I__6981\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32313\
        );

    \I__6980\ : InMux
    port map (
            O => \N__32322\,
            I => \N__32308\
        );

    \I__6979\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32308\
        );

    \I__6978\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32303\
        );

    \I__6977\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32303\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__32316\,
            I => \FTDI.un3_TX_0\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__32313\,
            I => \FTDI.un3_TX_0\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__32308\,
            I => \FTDI.un3_TX_0\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__32303\,
            I => \FTDI.un3_TX_0\
        );

    \I__6972\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32288\
        );

    \I__6971\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32285\
        );

    \I__6970\ : InMux
    port map (
            O => \N__32292\,
            I => \N__32282\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__32291\,
            I => \N__32279\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__32288\,
            I => \N__32276\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__32285\,
            I => \N__32273\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__32282\,
            I => \N__32270\
        );

    \I__6965\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32267\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__32276\,
            I => \N__32263\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__32273\,
            I => \N__32260\
        );

    \I__6962\ : Span4Mux_h
    port map (
            O => \N__32270\,
            I => \N__32257\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__32267\,
            I => \N__32254\
        );

    \I__6960\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32251\
        );

    \I__6959\ : Sp12to4
    port map (
            O => \N__32263\,
            I => \N__32248\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__32260\,
            I => \N__32245\
        );

    \I__6957\ : Span4Mux_v
    port map (
            O => \N__32257\,
            I => \N__32242\
        );

    \I__6956\ : Span4Mux_v
    port map (
            O => \N__32254\,
            I => \N__32239\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__32251\,
            I => \RXbuffer_4\
        );

    \I__6954\ : Odrv12
    port map (
            O => \N__32248\,
            I => \RXbuffer_4\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__32245\,
            I => \RXbuffer_4\
        );

    \I__6952\ : Odrv4
    port map (
            O => \N__32242\,
            I => \RXbuffer_4\
        );

    \I__6951\ : Odrv4
    port map (
            O => \N__32239\,
            I => \RXbuffer_4\
        );

    \I__6950\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__32225\,
            I => \N__32221\
        );

    \I__6948\ : InMux
    port map (
            O => \N__32224\,
            I => \N__32218\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__32221\,
            I => \N__32215\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__32218\,
            I => \N__32210\
        );

    \I__6945\ : Span4Mux_h
    port map (
            O => \N__32215\,
            I => \N__32207\
        );

    \I__6944\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32204\
        );

    \I__6943\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32201\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__32210\,
            I => \N__32198\
        );

    \I__6941\ : Span4Mux_h
    port map (
            O => \N__32207\,
            I => \N__32193\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__32204\,
            I => \N__32193\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32188\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__32198\,
            I => \N__32188\
        );

    \I__6937\ : Span4Mux_v
    port map (
            O => \N__32193\,
            I => \N__32185\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__32188\,
            I => \N__32181\
        );

    \I__6935\ : Span4Mux_h
    port map (
            O => \N__32185\,
            I => \N__32178\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__32184\,
            I => \N__32175\
        );

    \I__6933\ : Span4Mux_h
    port map (
            O => \N__32181\,
            I => \N__32172\
        );

    \I__6932\ : Span4Mux_h
    port map (
            O => \N__32178\,
            I => \N__32169\
        );

    \I__6931\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32166\
        );

    \I__6930\ : Span4Mux_h
    port map (
            O => \N__32172\,
            I => \N__32163\
        );

    \I__6929\ : Span4Mux_v
    port map (
            O => \N__32169\,
            I => \N__32160\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__32166\,
            I => \testWordZ0Z_12\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__32163\,
            I => \testWordZ0Z_12\
        );

    \I__6926\ : Odrv4
    port map (
            O => \N__32160\,
            I => \testWordZ0Z_12\
        );

    \I__6925\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__32147\,
            I => \TXbufferZ0Z_0\
        );

    \I__6922\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32141\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__32141\,
            I => \N__32138\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__32138\,
            I => \TXbufferZ0Z_3\
        );

    \I__6919\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__32132\,
            I => \FTDI.TXshiftZ0Z_5\
        );

    \I__6917\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32126\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__32126\,
            I => \N__32123\
        );

    \I__6915\ : Odrv12
    port map (
            O => \N__32123\,
            I => \TXbufferZ0Z_4\
        );

    \I__6914\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__32114\,
            I => \FTDI.TXshiftZ0Z_4\
        );

    \I__6911\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32108\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__32108\,
            I => \FTDI.TXshiftZ0Z_3\
        );

    \I__6909\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32099\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__32099\,
            I => \TXbufferZ0Z_2\
        );

    \I__6906\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__32093\,
            I => \N__32090\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__32090\,
            I => \TXbufferZ0Z_6\
        );

    \I__6903\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32084\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__32084\,
            I => \FTDI.TXshiftZ0Z_6\
        );

    \I__6901\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32074\
        );

    \I__6900\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32074\
        );

    \I__6899\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32070\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__32074\,
            I => \N__32062\
        );

    \I__6897\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32059\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__32070\,
            I => \N__32056\
        );

    \I__6895\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32053\
        );

    \I__6894\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32050\
        );

    \I__6893\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32044\
        );

    \I__6892\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32044\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__32065\,
            I => \N__32041\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__32062\,
            I => \N__32036\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__32059\,
            I => \N__32033\
        );

    \I__6888\ : Span4Mux_h
    port map (
            O => \N__32056\,
            I => \N__32028\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__32053\,
            I => \N__32028\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__32022\
        );

    \I__6885\ : InMux
    port map (
            O => \N__32049\,
            I => \N__32019\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__32044\,
            I => \N__32016\
        );

    \I__6883\ : InMux
    port map (
            O => \N__32041\,
            I => \N__32011\
        );

    \I__6882\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32006\
        );

    \I__6881\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32006\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__32036\,
            I => \N__31999\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__32033\,
            I => \N__31999\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__32028\,
            I => \N__31999\
        );

    \I__6877\ : InMux
    port map (
            O => \N__32027\,
            I => \N__31992\
        );

    \I__6876\ : InMux
    port map (
            O => \N__32026\,
            I => \N__31992\
        );

    \I__6875\ : InMux
    port map (
            O => \N__32025\,
            I => \N__31992\
        );

    \I__6874\ : Sp12to4
    port map (
            O => \N__32022\,
            I => \N__31987\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__32019\,
            I => \N__31987\
        );

    \I__6872\ : Span4Mux_v
    port map (
            O => \N__32016\,
            I => \N__31984\
        );

    \I__6871\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31979\
        );

    \I__6870\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31979\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__32011\,
            I => \aluOperand2_2_rep1\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__32006\,
            I => \aluOperand2_2_rep1\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__31999\,
            I => \aluOperand2_2_rep1\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__31992\,
            I => \aluOperand2_2_rep1\
        );

    \I__6865\ : Odrv12
    port map (
            O => \N__31987\,
            I => \aluOperand2_2_rep1\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__31984\,
            I => \aluOperand2_2_rep1\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__31979\,
            I => \aluOperand2_2_rep1\
        );

    \I__6862\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31960\
        );

    \I__6861\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31957\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31954\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__31957\,
            I => \ALU.bZ0Z_2\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__31954\,
            I => \ALU.bZ0Z_2\
        );

    \I__6857\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31946\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__31946\,
            I => \ALU.f_RNIESEJZ0Z_2\
        );

    \I__6855\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31940\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31937\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__31937\,
            I => \N__31934\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__31934\,
            I => \N__31930\
        );

    \I__6851\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31927\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__31930\,
            I => \ALU.gZ0Z_0\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__31927\,
            I => \ALU.gZ0Z_0\
        );

    \I__6848\ : CascadeMux
    port map (
            O => \N__31922\,
            I => \N__31918\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31915\
        );

    \I__6846\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31912\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__31915\,
            I => \N__31909\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__31912\,
            I => \N__31906\
        );

    \I__6843\ : Odrv4
    port map (
            O => \N__31909\,
            I => \ALU.gZ0Z_1\
        );

    \I__6842\ : Odrv12
    port map (
            O => \N__31906\,
            I => \ALU.gZ0Z_1\
        );

    \I__6841\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31898\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31895\
        );

    \I__6839\ : Span4Mux_h
    port map (
            O => \N__31895\,
            I => \N__31891\
        );

    \I__6838\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31888\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__31891\,
            I => \ALU.gZ0Z_2\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__31888\,
            I => \ALU.gZ0Z_2\
        );

    \I__6835\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31880\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31876\
        );

    \I__6833\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31873\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__31876\,
            I => \N__31870\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__31873\,
            I => \N__31867\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__31870\,
            I => \ALU.gZ0Z_3\
        );

    \I__6829\ : Odrv12
    port map (
            O => \N__31867\,
            I => \ALU.gZ0Z_3\
        );

    \I__6828\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31858\
        );

    \I__6827\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31855\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__31858\,
            I => \N__31852\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__31855\,
            I => \N__31849\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__31852\,
            I => \N__31846\
        );

    \I__6823\ : Span4Mux_v
    port map (
            O => \N__31849\,
            I => \N__31843\
        );

    \I__6822\ : Span4Mux_h
    port map (
            O => \N__31846\,
            I => \N__31840\
        );

    \I__6821\ : Odrv4
    port map (
            O => \N__31843\,
            I => \ALU.gZ0Z_4\
        );

    \I__6820\ : Odrv4
    port map (
            O => \N__31840\,
            I => \ALU.gZ0Z_4\
        );

    \I__6819\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31832\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__6817\ : Span4Mux_v
    port map (
            O => \N__31829\,
            I => \N__31826\
        );

    \I__6816\ : Span4Mux_h
    port map (
            O => \N__31826\,
            I => \N__31822\
        );

    \I__6815\ : InMux
    port map (
            O => \N__31825\,
            I => \N__31819\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__31822\,
            I => \ALU.gZ0Z_5\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__31819\,
            I => \ALU.gZ0Z_5\
        );

    \I__6812\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__31808\,
            I => \N__31804\
        );

    \I__6809\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31801\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__31804\,
            I => \N__31798\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31795\
        );

    \I__6806\ : Odrv4
    port map (
            O => \N__31798\,
            I => \ALU.gZ0Z_7\
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__31795\,
            I => \ALU.gZ0Z_7\
        );

    \I__6804\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31787\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__31787\,
            I => \N__31784\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__31784\,
            I => \N__31780\
        );

    \I__6801\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31777\
        );

    \I__6800\ : Odrv4
    port map (
            O => \N__31780\,
            I => \ALU.N_578\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__31777\,
            I => \ALU.N_578\
        );

    \I__6798\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31768\
        );

    \I__6797\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31764\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31761\
        );

    \I__6795\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31758\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__31764\,
            I => \ALU.N_477\
        );

    \I__6793\ : Odrv12
    port map (
            O => \N__31761\,
            I => \ALU.N_477\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__31758\,
            I => \ALU.N_477\
        );

    \I__6791\ : InMux
    port map (
            O => \N__31751\,
            I => \N__31748\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__31748\,
            I => \ALU.N_634\
        );

    \I__6789\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31742\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__31742\,
            I => \N__31738\
        );

    \I__6787\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31735\
        );

    \I__6786\ : Span4Mux_h
    port map (
            O => \N__31738\,
            I => \N__31732\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__31735\,
            I => \N__31729\
        );

    \I__6784\ : Odrv4
    port map (
            O => \N__31732\,
            I => \ALU.aZ0Z_15\
        );

    \I__6783\ : Odrv4
    port map (
            O => \N__31729\,
            I => \ALU.aZ0Z_15\
        );

    \I__6782\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31721\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__31721\,
            I => \N__31718\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__31718\,
            I => \N__31715\
        );

    \I__6779\ : Span4Mux_h
    port map (
            O => \N__31715\,
            I => \N__31712\
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__31712\,
            I => \ALU.f_RNI0P6LZ0Z_1\
        );

    \I__6777\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31706\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__31706\,
            I => \N__31703\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__31703\,
            I => \N__31700\
        );

    \I__6774\ : Span4Mux_h
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__6773\ : Odrv4
    port map (
            O => \N__31697\,
            I => \ALU.f_RNICQEJZ0Z_1\
        );

    \I__6772\ : InMux
    port map (
            O => \N__31694\,
            I => \N__31691\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__31691\,
            I => \N__31687\
        );

    \I__6770\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31684\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__31687\,
            I => \N__31681\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__31684\,
            I => \N__31678\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__31681\,
            I => \N__31673\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__31678\,
            I => \N__31673\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__31673\,
            I => \ALU.cZ0Z_7\
        );

    \I__6764\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31667\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31664\
        );

    \I__6762\ : Span4Mux_h
    port map (
            O => \N__31664\,
            I => \N__31661\
        );

    \I__6761\ : Span4Mux_h
    port map (
            O => \N__31661\,
            I => \N__31658\
        );

    \I__6760\ : Odrv4
    port map (
            O => \N__31658\,
            I => \ALU.g_RNIQCLLZ0Z_7\
        );

    \I__6759\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31652\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__31652\,
            I => \N__31649\
        );

    \I__6757\ : Odrv12
    port map (
            O => \N__31649\,
            I => \ALU.f_RNIL2FJZ0Z_5\
        );

    \I__6756\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31643\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__31643\,
            I => \N__31640\
        );

    \I__6754\ : Span4Mux_v
    port map (
            O => \N__31640\,
            I => \N__31637\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__31637\,
            I => \N__31634\
        );

    \I__6752\ : Span4Mux_v
    port map (
            O => \N__31634\,
            I => \N__31631\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__31631\,
            I => \ALU.m286_bmZ0\
        );

    \I__6750\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31625\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__6748\ : Span4Mux_v
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__6747\ : Span4Mux_h
    port map (
            O => \N__31619\,
            I => \N__31616\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__31616\,
            I => \N__31613\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__31613\,
            I => \N__31610\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__31610\,
            I => \ALU.m286_amZ0\
        );

    \I__6743\ : InMux
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__31604\,
            I => \N__31601\
        );

    \I__6741\ : Odrv12
    port map (
            O => \N__31601\,
            I => \ALU.f_RNIAOEJZ0Z_0\
        );

    \I__6740\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31594\
        );

    \I__6739\ : InMux
    port map (
            O => \N__31597\,
            I => \N__31590\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__31594\,
            I => \N__31587\
        );

    \I__6737\ : CascadeMux
    port map (
            O => \N__31593\,
            I => \N__31584\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__31590\,
            I => \N__31581\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__31587\,
            I => \N__31578\
        );

    \I__6734\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31574\
        );

    \I__6733\ : Span4Mux_h
    port map (
            O => \N__31581\,
            I => \N__31571\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__31578\,
            I => \N__31568\
        );

    \I__6731\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31565\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__31574\,
            I => \aluOperand2_fast_0\
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__31571\,
            I => \aluOperand2_fast_0\
        );

    \I__6728\ : Odrv4
    port map (
            O => \N__31568\,
            I => \aluOperand2_fast_0\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__31565\,
            I => \aluOperand2_fast_0\
        );

    \I__6726\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__6724\ : Span4Mux_h
    port map (
            O => \N__31550\,
            I => \N__31547\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__6722\ : Span4Mux_h
    port map (
            O => \N__31544\,
            I => \N__31540\
        );

    \I__6721\ : InMux
    port map (
            O => \N__31543\,
            I => \N__31537\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__31540\,
            I => \ALU.cZ0Z_14\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__31537\,
            I => \ALU.cZ0Z_14\
        );

    \I__6718\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31529\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__6716\ : Odrv12
    port map (
            O => \N__31526\,
            I => \ALU.c_RNIND49Z0Z_14\
        );

    \I__6715\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31519\
        );

    \I__6714\ : InMux
    port map (
            O => \N__31522\,
            I => \N__31516\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__31519\,
            I => \N__31513\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__31516\,
            I => \N__31510\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__31513\,
            I => \N__31507\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__31510\,
            I => \ALU.cZ0Z_15\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__31507\,
            I => \ALU.cZ0Z_15\
        );

    \I__6708\ : CEMux
    port map (
            O => \N__31502\,
            I => \N__31499\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__31499\,
            I => \N__31494\
        );

    \I__6706\ : CEMux
    port map (
            O => \N__31498\,
            I => \N__31491\
        );

    \I__6705\ : CEMux
    port map (
            O => \N__31497\,
            I => \N__31488\
        );

    \I__6704\ : Span4Mux_h
    port map (
            O => \N__31494\,
            I => \N__31485\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__31491\,
            I => \N__31482\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__31488\,
            I => \N__31479\
        );

    \I__6701\ : Span4Mux_v
    port map (
            O => \N__31485\,
            I => \N__31476\
        );

    \I__6700\ : Span4Mux_s1_v
    port map (
            O => \N__31482\,
            I => \N__31473\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__31479\,
            I => \N__31470\
        );

    \I__6698\ : Span4Mux_v
    port map (
            O => \N__31476\,
            I => \N__31467\
        );

    \I__6697\ : Span4Mux_v
    port map (
            O => \N__31473\,
            I => \N__31464\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__31470\,
            I => \N__31461\
        );

    \I__6695\ : Span4Mux_v
    port map (
            O => \N__31467\,
            I => \N__31458\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__31464\,
            I => \N__31455\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__31461\,
            I => \N__31452\
        );

    \I__6692\ : Span4Mux_h
    port map (
            O => \N__31458\,
            I => \N__31449\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__31455\,
            I => \ALU.c_cnvZ0Z_0\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__31452\,
            I => \ALU.c_cnvZ0Z_0\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__31449\,
            I => \ALU.c_cnvZ0Z_0\
        );

    \I__6688\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31436\
        );

    \I__6687\ : InMux
    port map (
            O => \N__31441\,
            I => \N__31436\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__31436\,
            I => \N__31433\
        );

    \I__6685\ : Span4Mux_v
    port map (
            O => \N__31433\,
            I => \N__31430\
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__31430\,
            I => \ALU.hZ0Z_1\
        );

    \I__6683\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31424\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31420\
        );

    \I__6681\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31417\
        );

    \I__6680\ : Span4Mux_h
    port map (
            O => \N__31420\,
            I => \N__31412\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__31417\,
            I => \N__31412\
        );

    \I__6678\ : Span4Mux_v
    port map (
            O => \N__31412\,
            I => \N__31409\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__31409\,
            I => \ALU.hZ0Z_2\
        );

    \I__6676\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31403\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__31403\,
            I => \N__31400\
        );

    \I__6674\ : Span4Mux_h
    port map (
            O => \N__31400\,
            I => \N__31397\
        );

    \I__6673\ : Span4Mux_v
    port map (
            O => \N__31397\,
            I => \N__31393\
        );

    \I__6672\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31390\
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__31393\,
            I => \ALU.hZ0Z_5\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__31390\,
            I => \ALU.hZ0Z_5\
        );

    \I__6669\ : InMux
    port map (
            O => \N__31385\,
            I => \N__31382\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__6667\ : Span4Mux_h
    port map (
            O => \N__31379\,
            I => \N__31375\
        );

    \I__6666\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31372\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__31375\,
            I => \N__31367\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__31372\,
            I => \N__31367\
        );

    \I__6663\ : Span4Mux_v
    port map (
            O => \N__31367\,
            I => \N__31364\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__31364\,
            I => \ALU.aZ0Z_14\
        );

    \I__6661\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31357\
        );

    \I__6660\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31354\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__31357\,
            I => \ALU.eZ0Z_15\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__31354\,
            I => \ALU.eZ0Z_15\
        );

    \I__6657\ : CascadeMux
    port map (
            O => \N__31349\,
            I => \ALU.a_RNILVBOZ0Z_15_cascade_\
        );

    \I__6656\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31343\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__31343\,
            I => \ALU.c_RNIPF49Z0Z_15\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__31340\,
            I => \ALU.operand2_7_ns_1_15_cascade_\
        );

    \I__6653\ : InMux
    port map (
            O => \N__31337\,
            I => \N__31334\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__31334\,
            I => \N__31331\
        );

    \I__6651\ : Span4Mux_v
    port map (
            O => \N__31331\,
            I => \N__31328\
        );

    \I__6650\ : Span4Mux_v
    port map (
            O => \N__31328\,
            I => \N__31325\
        );

    \I__6649\ : Odrv4
    port map (
            O => \N__31325\,
            I => \ALU.b_RNIORSD1Z0Z_15\
        );

    \I__6648\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31319\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__31319\,
            I => \N__31316\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__31316\,
            I => \N__31313\
        );

    \I__6645\ : Span4Mux_h
    port map (
            O => \N__31313\,
            I => \N__31310\
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__31310\,
            I => \ALU.operand2_15\
        );

    \I__6643\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31304\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__6641\ : Span4Mux_v
    port map (
            O => \N__31301\,
            I => \N__31297\
        );

    \I__6640\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31294\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__31297\,
            I => \N__31289\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__31294\,
            I => \N__31289\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__31289\,
            I => \ALU.cZ0Z_11\
        );

    \I__6636\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31283\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__31283\,
            I => \N__31279\
        );

    \I__6634\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31276\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__31279\,
            I => \N__31271\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31271\
        );

    \I__6631\ : Span4Mux_h
    port map (
            O => \N__31271\,
            I => \N__31268\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__31268\,
            I => \ALU.cZ0Z_12\
        );

    \I__6629\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31257\
        );

    \I__6628\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31254\
        );

    \I__6627\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31251\
        );

    \I__6626\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31246\
        );

    \I__6625\ : InMux
    port map (
            O => \N__31261\,
            I => \N__31243\
        );

    \I__6624\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31240\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__31257\,
            I => \N__31237\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31234\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31231\
        );

    \I__6620\ : CascadeMux
    port map (
            O => \N__31250\,
            I => \N__31228\
        );

    \I__6619\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31225\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31212\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__31243\,
            I => \N__31212\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__31240\,
            I => \N__31212\
        );

    \I__6615\ : Span4Mux_h
    port map (
            O => \N__31237\,
            I => \N__31212\
        );

    \I__6614\ : Span4Mux_v
    port map (
            O => \N__31234\,
            I => \N__31212\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__31231\,
            I => \N__31212\
        );

    \I__6612\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31209\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__31225\,
            I => \N__31206\
        );

    \I__6610\ : Span4Mux_v
    port map (
            O => \N__31212\,
            I => \N__31203\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31198\
        );

    \I__6608\ : Span12Mux_h
    port map (
            O => \N__31206\,
            I => \N__31198\
        );

    \I__6607\ : Odrv4
    port map (
            O => \N__31203\,
            I => \aluOperand2_0_rep1\
        );

    \I__6606\ : Odrv12
    port map (
            O => \N__31198\,
            I => \aluOperand2_0_rep1\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__31193\,
            I => \ALU.a_RNICNBOZ0Z_11_cascade_\
        );

    \I__6604\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \ALU.operand2_7_ns_1_11_cascade_\
        );

    \I__6603\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31184\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__31184\,
            I => \ALU.b_RNIGJSD1Z0Z_11\
        );

    \I__6601\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31177\
        );

    \I__6600\ : CascadeMux
    port map (
            O => \N__31180\,
            I => \N__31174\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__31177\,
            I => \N__31171\
        );

    \I__6598\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31168\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__31171\,
            I => \N__31165\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31162\
        );

    \I__6595\ : Odrv4
    port map (
            O => \N__31165\,
            I => \ALU.operand2_11\
        );

    \I__6594\ : Odrv12
    port map (
            O => \N__31162\,
            I => \ALU.operand2_11\
        );

    \I__6593\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31154\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__31154\,
            I => \N__31150\
        );

    \I__6591\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31147\
        );

    \I__6590\ : Odrv12
    port map (
            O => \N__31150\,
            I => \ALU.dZ0Z_11\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__31147\,
            I => \ALU.dZ0Z_11\
        );

    \I__6588\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__31139\,
            I => \ALU.d_RNIK3LUZ0Z_11\
        );

    \I__6586\ : InMux
    port map (
            O => \N__31136\,
            I => \N__31133\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__6584\ : Span4Mux_v
    port map (
            O => \N__31130\,
            I => \N__31126\
        );

    \I__6583\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31123\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__31126\,
            I => \ALU.hZ0Z_11\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__31123\,
            I => \ALU.hZ0Z_11\
        );

    \I__6580\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31115\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__31115\,
            I => \ALU.c_RNIG749Z0Z_11\
        );

    \I__6578\ : CascadeMux
    port map (
            O => \N__31112\,
            I => \ALU.a_RNIHRBOZ0Z_13_cascade_\
        );

    \I__6577\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31106\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__31106\,
            I => \ALU.c_RNILB49Z0Z_13\
        );

    \I__6575\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31100\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__31100\,
            I => \N__31097\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__31097\,
            I => \N__31093\
        );

    \I__6572\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__31090\,
            I => \ALU.operand2_7_ns_1_13\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__31087\,
            I => \ALU.operand2_7_ns_1_13\
        );

    \I__6568\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31076\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__6565\ : Span4Mux_h
    port map (
            O => \N__31073\,
            I => \N__31070\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__31070\,
            I => \ALU.un2_addsub_cry_7_c_RNIL8JHGZ0\
        );

    \I__6563\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31064\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__31064\,
            I => \N__31061\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__31061\,
            I => \N__31057\
        );

    \I__6560\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31054\
        );

    \I__6559\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31051\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__31054\,
            I => \ALU.aZ0Z_8\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__31051\,
            I => \ALU.aZ0Z_8\
        );

    \I__6556\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31038\
        );

    \I__6555\ : CascadeMux
    port map (
            O => \N__31045\,
            I => \N__31035\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__31044\,
            I => \N__31032\
        );

    \I__6553\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31029\
        );

    \I__6552\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31026\
        );

    \I__6551\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31023\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__31038\,
            I => \N__31020\
        );

    \I__6549\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31015\
        );

    \I__6548\ : InMux
    port map (
            O => \N__31032\,
            I => \N__31015\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__31029\,
            I => \N__31010\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__31026\,
            I => \N__31007\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__31023\,
            I => \N__31004\
        );

    \I__6544\ : Span4Mux_v
    port map (
            O => \N__31020\,
            I => \N__30999\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__31015\,
            I => \N__30999\
        );

    \I__6542\ : InMux
    port map (
            O => \N__31014\,
            I => \N__30994\
        );

    \I__6541\ : InMux
    port map (
            O => \N__31013\,
            I => \N__30994\
        );

    \I__6540\ : Span4Mux_v
    port map (
            O => \N__31010\,
            I => \N__30991\
        );

    \I__6539\ : Span4Mux_v
    port map (
            O => \N__31007\,
            I => \N__30988\
        );

    \I__6538\ : Span4Mux_h
    port map (
            O => \N__31004\,
            I => \N__30983\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__30999\,
            I => \N__30983\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__30994\,
            I => \aluOperand2_fast_1\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__30991\,
            I => \aluOperand2_fast_1\
        );

    \I__6534\ : Odrv4
    port map (
            O => \N__30988\,
            I => \aluOperand2_fast_1\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__30983\,
            I => \aluOperand2_fast_1\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__30974\,
            I => \N__30970\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__30973\,
            I => \N__30967\
        );

    \I__6530\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30964\
        );

    \I__6529\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30961\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__30964\,
            I => \N__30958\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30955\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__30958\,
            I => \N__30952\
        );

    \I__6525\ : Span4Mux_v
    port map (
            O => \N__30955\,
            I => \N__30949\
        );

    \I__6524\ : Span4Mux_h
    port map (
            O => \N__30952\,
            I => \N__30946\
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__30949\,
            I => \ALU.eZ0Z_8\
        );

    \I__6522\ : Odrv4
    port map (
            O => \N__30946\,
            I => \ALU.eZ0Z_8\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__6520\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30934\
        );

    \I__6519\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30931\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__30934\,
            I => \N__30928\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__30931\,
            I => \N__30925\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__30928\,
            I => \N__30922\
        );

    \I__6515\ : Span4Mux_v
    port map (
            O => \N__30925\,
            I => \N__30919\
        );

    \I__6514\ : Span4Mux_v
    port map (
            O => \N__30922\,
            I => \N__30916\
        );

    \I__6513\ : Sp12to4
    port map (
            O => \N__30919\,
            I => \N__30913\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__30916\,
            I => \ALU.gZ0Z_8\
        );

    \I__6511\ : Odrv12
    port map (
            O => \N__30913\,
            I => \ALU.gZ0Z_8\
        );

    \I__6510\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30905\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__30905\,
            I => \N__30902\
        );

    \I__6508\ : Span4Mux_h
    port map (
            O => \N__30902\,
            I => \N__30898\
        );

    \I__6507\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30895\
        );

    \I__6506\ : Span4Mux_v
    port map (
            O => \N__30898\,
            I => \N__30892\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30889\
        );

    \I__6504\ : Span4Mux_v
    port map (
            O => \N__30892\,
            I => \N__30886\
        );

    \I__6503\ : Span4Mux_v
    port map (
            O => \N__30889\,
            I => \N__30883\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__30886\,
            I => \ALU.cZ0Z_8\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__30883\,
            I => \ALU.cZ0Z_8\
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__30878\,
            I => \ALU.operand2_3_ns_1_8_cascade_\
        );

    \I__6499\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30872\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__30872\,
            I => \N__30869\
        );

    \I__6497\ : Span4Mux_s3_h
    port map (
            O => \N__30869\,
            I => \N__30866\
        );

    \I__6496\ : Span4Mux_h
    port map (
            O => \N__30866\,
            I => \N__30863\
        );

    \I__6495\ : Odrv4
    port map (
            O => \N__30863\,
            I => \ALU.N_819\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__30860\,
            I => \ALU.addsub_0_sqmuxa_cascade_\
        );

    \I__6493\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30854\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__30854\,
            I => \N__30851\
        );

    \I__6491\ : Span12Mux_h
    port map (
            O => \N__30851\,
            I => \N__30848\
        );

    \I__6490\ : Odrv12
    port map (
            O => \N__30848\,
            I => \ALU.un2_addsub_cry_8_c_RNIKR81JZ0\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__30845\,
            I => \ALU.un9_addsub_cry_8_c_RNIKTS9SZ0_cascade_\
        );

    \I__6488\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__30839\,
            I => \N__30836\
        );

    \I__6486\ : Odrv4
    port map (
            O => \N__30836\,
            I => \ALU.a_15_m5_9\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__30833\,
            I => \ALU.a_15_ns_1_9_cascade_\
        );

    \I__6484\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30827\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__30827\,
            I => \N__30823\
        );

    \I__6482\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30820\
        );

    \I__6481\ : Span4Mux_v
    port map (
            O => \N__30823\,
            I => \N__30817\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30814\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__30817\,
            I => \ALU.eZ0Z_11\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__30814\,
            I => \ALU.eZ0Z_11\
        );

    \I__6477\ : CascadeMux
    port map (
            O => \N__30809\,
            I => \N__30802\
        );

    \I__6476\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30797\
        );

    \I__6475\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30797\
        );

    \I__6474\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30794\
        );

    \I__6473\ : InMux
    port map (
            O => \N__30805\,
            I => \N__30789\
        );

    \I__6472\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30789\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__30797\,
            I => \N__30784\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30784\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__30789\,
            I => \N__30775\
        );

    \I__6468\ : Span4Mux_v
    port map (
            O => \N__30784\,
            I => \N__30775\
        );

    \I__6467\ : CascadeMux
    port map (
            O => \N__30783\,
            I => \N__30772\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__30782\,
            I => \N__30769\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__30781\,
            I => \N__30766\
        );

    \I__6464\ : CascadeMux
    port map (
            O => \N__30780\,
            I => \N__30763\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__30775\,
            I => \N__30760\
        );

    \I__6462\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30757\
        );

    \I__6461\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30750\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30750\
        );

    \I__6459\ : InMux
    port map (
            O => \N__30763\,
            I => \N__30750\
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__30760\,
            I => \testStateZ0Z_2\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__30757\,
            I => \testStateZ0Z_2\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__30750\,
            I => \testStateZ0Z_2\
        );

    \I__6455\ : IoInMux
    port map (
            O => \N__30743\,
            I => \N__30740\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__30740\,
            I => \N__30737\
        );

    \I__6453\ : Span12Mux_s0_h
    port map (
            O => \N__30737\,
            I => \N__30734\
        );

    \I__6452\ : Span12Mux_v
    port map (
            O => \N__30734\,
            I => \N__30731\
        );

    \I__6451\ : Odrv12
    port map (
            O => \N__30731\,
            I => \testState_i_2\
        );

    \I__6450\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30725\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30722\
        );

    \I__6448\ : Span4Mux_h
    port map (
            O => \N__30722\,
            I => \N__30718\
        );

    \I__6447\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30715\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__30718\,
            I => \N__30710\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30710\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__30710\,
            I => \N__30707\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__30707\,
            I => \ALU.eZ0Z_14\
        );

    \I__6442\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30701\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__30701\,
            I => \N__30698\
        );

    \I__6440\ : Span4Mux_v
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__6438\ : Span4Mux_h
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__30689\,
            I => \ALU.un2_addsub_cry_13_c_RNINVE5KZ0\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__30686\,
            I => \un2_addsub_cry_13_c_RNI2LH1U_cascade_\
        );

    \I__6435\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__30680\,
            I => \N__30677\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__30677\,
            I => \N__30674\
        );

    \I__6432\ : Span4Mux_h
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__30671\,
            I => \c_RNIFCGVL2_14\
        );

    \I__6430\ : CascadeMux
    port map (
            O => \N__30668\,
            I => \aluOperation_RNIR872K3_0_cascade_\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__6428\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30659\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__30659\,
            I => \ALU.a_RNIJTBOZ0Z_14\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__30656\,
            I => \ALU.operand2_7_ns_1_14_cascade_\
        );

    \I__6425\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30650\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__30650\,
            I => \ALU.b_RNIMPSD1Z0Z_14\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__30647\,
            I => \N__30643\
        );

    \I__6422\ : CascadeMux
    port map (
            O => \N__30646\,
            I => \N__30640\
        );

    \I__6421\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30635\
        );

    \I__6420\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30635\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__30635\,
            I => \N__30631\
        );

    \I__6418\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30628\
        );

    \I__6417\ : Span12Mux_s5_v
    port map (
            O => \N__30631\,
            I => \N__30623\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__30628\,
            I => \N__30623\
        );

    \I__6415\ : Odrv12
    port map (
            O => \N__30623\,
            I => \ALU.operand2_14\
        );

    \I__6414\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30617\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__30617\,
            I => \N__30614\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__30614\,
            I => \N__30611\
        );

    \I__6411\ : Span4Mux_s3_h
    port map (
            O => \N__30611\,
            I => \N__30607\
        );

    \I__6410\ : InMux
    port map (
            O => \N__30610\,
            I => \N__30604\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__30607\,
            I => \N__30601\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__30604\,
            I => \ALU.hZ0Z_14\
        );

    \I__6407\ : Odrv4
    port map (
            O => \N__30601\,
            I => \ALU.hZ0Z_14\
        );

    \I__6406\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__30593\,
            I => \N__30590\
        );

    \I__6404\ : Span4Mux_h
    port map (
            O => \N__30590\,
            I => \N__30586\
        );

    \I__6403\ : InMux
    port map (
            O => \N__30589\,
            I => \N__30583\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__30586\,
            I => \N__30580\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__30583\,
            I => \N__30577\
        );

    \I__6400\ : Span4Mux_v
    port map (
            O => \N__30580\,
            I => \N__30574\
        );

    \I__6399\ : Span4Mux_h
    port map (
            O => \N__30577\,
            I => \N__30571\
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__30574\,
            I => \ALU.dZ0Z_14\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__30571\,
            I => \ALU.dZ0Z_14\
        );

    \I__6396\ : InMux
    port map (
            O => \N__30566\,
            I => \N__30563\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__30563\,
            I => \ALU.d_RNIQ9LUZ0Z_14\
        );

    \I__6394\ : CascadeMux
    port map (
            O => \N__30560\,
            I => \ALU.c_RNI1OCN4Z0Z_15_cascade_\
        );

    \I__6393\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30553\
        );

    \I__6392\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30550\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__30553\,
            I => \N__30547\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__30550\,
            I => \N__30544\
        );

    \I__6389\ : Span12Mux_h
    port map (
            O => \N__30547\,
            I => \N__30539\
        );

    \I__6388\ : Span12Mux_s5_h
    port map (
            O => \N__30544\,
            I => \N__30539\
        );

    \I__6387\ : Odrv12
    port map (
            O => \N__30539\,
            I => \ALU.N_762\
        );

    \I__6386\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30532\
        );

    \I__6385\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30526\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30523\
        );

    \I__6382\ : Span4Mux_h
    port map (
            O => \N__30526\,
            I => \N__30520\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__30523\,
            I => \N__30517\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__30520\,
            I => \N__30514\
        );

    \I__6379\ : Span4Mux_v
    port map (
            O => \N__30517\,
            I => \N__30509\
        );

    \I__6378\ : Span4Mux_h
    port map (
            O => \N__30514\,
            I => \N__30509\
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__30509\,
            I => \ALU.N_714\
        );

    \I__6376\ : CascadeMux
    port map (
            O => \N__30506\,
            I => \ALU.N_621_1_cascade_\
        );

    \I__6375\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30499\
        );

    \I__6374\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30496\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__30499\,
            I => \N__30492\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30489\
        );

    \I__6371\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30486\
        );

    \I__6370\ : Odrv4
    port map (
            O => \N__30492\,
            I => \ALU.N_589\
        );

    \I__6369\ : Odrv4
    port map (
            O => \N__30489\,
            I => \ALU.N_589\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__30486\,
            I => \ALU.N_589\
        );

    \I__6367\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30472\
        );

    \I__6366\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30472\
        );

    \I__6365\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30466\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__30472\,
            I => \N__30463\
        );

    \I__6363\ : InMux
    port map (
            O => \N__30471\,
            I => \N__30460\
        );

    \I__6362\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30455\
        );

    \I__6361\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30455\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30452\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__30463\,
            I => \ALU.N_621_1\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__30460\,
            I => \ALU.N_621_1\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__30455\,
            I => \ALU.N_621_1\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__30452\,
            I => \ALU.N_621_1\
        );

    \I__6355\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30440\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__30440\,
            I => \ALU.c_RNI4JFV4_0Z0Z_15\
        );

    \I__6353\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30434\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__30434\,
            I => \N__30431\
        );

    \I__6351\ : Odrv12
    port map (
            O => \N__30431\,
            I => \ALU.N_274_0\
        );

    \I__6350\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__30425\,
            I => \ALU.d_RNI36KJ21Z0Z_9\
        );

    \I__6348\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30419\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__30419\,
            I => \N__30414\
        );

    \I__6346\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30411\
        );

    \I__6345\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30407\
        );

    \I__6344\ : Span4Mux_s2_v
    port map (
            O => \N__30414\,
            I => \N__30404\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30401\
        );

    \I__6342\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30398\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30395\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__30404\,
            I => \FTDI.TXready\
        );

    \I__6339\ : Odrv4
    port map (
            O => \N__30401\,
            I => \FTDI.TXready\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__30398\,
            I => \FTDI.TXready\
        );

    \I__6337\ : Odrv12
    port map (
            O => \N__30395\,
            I => \FTDI.TXready\
        );

    \I__6336\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30381\
        );

    \I__6335\ : InMux
    port map (
            O => \N__30385\,
            I => \N__30372\
        );

    \I__6334\ : InMux
    port map (
            O => \N__30384\,
            I => \N__30372\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__30381\,
            I => \N__30369\
        );

    \I__6332\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30366\
        );

    \I__6331\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30359\
        );

    \I__6330\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30359\
        );

    \I__6329\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30359\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__30372\,
            I => \N__30356\
        );

    \I__6327\ : Span4Mux_v
    port map (
            O => \N__30369\,
            I => \N__30349\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__30366\,
            I => \N__30349\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__30359\,
            I => \N__30349\
        );

    \I__6324\ : Span4Mux_h
    port map (
            O => \N__30356\,
            I => \N__30346\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__30349\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__30346\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__6321\ : InMux
    port map (
            O => \N__30341\,
            I => \N__30338\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30333\
        );

    \I__6319\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30328\
        );

    \I__6318\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30328\
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__30333\,
            I => \TXstartZ0\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__30328\,
            I => \TXstartZ0\
        );

    \I__6315\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30319\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__30322\,
            I => \N__30316\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__30319\,
            I => \N__30311\
        );

    \I__6312\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30306\
        );

    \I__6311\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30306\
        );

    \I__6310\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30303\
        );

    \I__6309\ : Span4Mux_v
    port map (
            O => \N__30311\,
            I => \N__30299\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__30306\,
            I => \N__30296\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__30303\,
            I => \N__30293\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__30302\,
            I => \N__30286\
        );

    \I__6305\ : Sp12to4
    port map (
            O => \N__30299\,
            I => \N__30282\
        );

    \I__6304\ : Span4Mux_v
    port map (
            O => \N__30296\,
            I => \N__30279\
        );

    \I__6303\ : Span4Mux_s2_v
    port map (
            O => \N__30293\,
            I => \N__30276\
        );

    \I__6302\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30269\
        );

    \I__6301\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30269\
        );

    \I__6300\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30269\
        );

    \I__6299\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30264\
        );

    \I__6298\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30264\
        );

    \I__6297\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30261\
        );

    \I__6296\ : Span12Mux_s6_h
    port map (
            O => \N__30282\,
            I => \N__30258\
        );

    \I__6295\ : Span4Mux_h
    port map (
            O => \N__30279\,
            I => \N__30253\
        );

    \I__6294\ : Span4Mux_h
    port map (
            O => \N__30276\,
            I => \N__30253\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__30269\,
            I => \N__30250\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__30264\,
            I => \testStateZ0Z_0\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__30261\,
            I => \testStateZ0Z_0\
        );

    \I__6290\ : Odrv12
    port map (
            O => \N__30258\,
            I => \testStateZ0Z_0\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__30253\,
            I => \testStateZ0Z_0\
        );

    \I__6288\ : Odrv12
    port map (
            O => \N__30250\,
            I => \testStateZ0Z_0\
        );

    \I__6287\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30235\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__30238\,
            I => \N__30231\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30228\
        );

    \I__6284\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30223\
        );

    \I__6283\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30223\
        );

    \I__6282\ : Odrv12
    port map (
            O => \N__30228\,
            I => \ctrlOut_13\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__30223\,
            I => \ctrlOut_13\
        );

    \I__6280\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30212\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__30217\,
            I => \N__30208\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__30216\,
            I => \N__30202\
        );

    \I__6277\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30197\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__30212\,
            I => \N__30189\
        );

    \I__6275\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30186\
        );

    \I__6274\ : InMux
    port map (
            O => \N__30208\,
            I => \N__30181\
        );

    \I__6273\ : InMux
    port map (
            O => \N__30207\,
            I => \N__30181\
        );

    \I__6272\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30176\
        );

    \I__6271\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30176\
        );

    \I__6270\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30173\
        );

    \I__6269\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30167\
        );

    \I__6268\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30164\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__30197\,
            I => \N__30161\
        );

    \I__6266\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30158\
        );

    \I__6265\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30153\
        );

    \I__6264\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30153\
        );

    \I__6263\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30148\
        );

    \I__6262\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30148\
        );

    \I__6261\ : Span4Mux_h
    port map (
            O => \N__30189\,
            I => \N__30143\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__30186\,
            I => \N__30143\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__30181\,
            I => \N__30140\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__30176\,
            I => \N__30137\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__30173\,
            I => \N__30132\
        );

    \I__6256\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30122\
        );

    \I__6255\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30122\
        );

    \I__6254\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30122\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__30167\,
            I => \N__30117\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__30164\,
            I => \N__30117\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__30161\,
            I => \N__30112\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__30158\,
            I => \N__30112\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__30153\,
            I => \N__30109\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__30148\,
            I => \N__30106\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__30143\,
            I => \N__30103\
        );

    \I__6246\ : Span4Mux_v
    port map (
            O => \N__30140\,
            I => \N__30098\
        );

    \I__6245\ : Span4Mux_s1_h
    port map (
            O => \N__30137\,
            I => \N__30098\
        );

    \I__6244\ : InMux
    port map (
            O => \N__30136\,
            I => \N__30093\
        );

    \I__6243\ : InMux
    port map (
            O => \N__30135\,
            I => \N__30093\
        );

    \I__6242\ : Span4Mux_v
    port map (
            O => \N__30132\,
            I => \N__30090\
        );

    \I__6241\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30083\
        );

    \I__6240\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30083\
        );

    \I__6239\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30083\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__30122\,
            I => \N__30074\
        );

    \I__6237\ : Span4Mux_h
    port map (
            O => \N__30117\,
            I => \N__30074\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__30112\,
            I => \N__30074\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__30109\,
            I => \N__30074\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__30106\,
            I => \busState_2\
        );

    \I__6233\ : Odrv4
    port map (
            O => \N__30103\,
            I => \busState_2\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__30098\,
            I => \busState_2\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__30093\,
            I => \busState_2\
        );

    \I__6230\ : Odrv4
    port map (
            O => \N__30090\,
            I => \busState_2\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__30083\,
            I => \busState_2\
        );

    \I__6228\ : Odrv4
    port map (
            O => \N__30074\,
            I => \busState_2\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__30059\,
            I => \N__30051\
        );

    \I__6226\ : CascadeMux
    port map (
            O => \N__30058\,
            I => \N__30046\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__30057\,
            I => \N__30042\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__30056\,
            I => \N__30039\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__30055\,
            I => \N__30036\
        );

    \I__6222\ : CascadeMux
    port map (
            O => \N__30054\,
            I => \N__30033\
        );

    \I__6221\ : InMux
    port map (
            O => \N__30051\,
            I => \N__30027\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__30050\,
            I => \N__30018\
        );

    \I__6219\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30015\
        );

    \I__6218\ : InMux
    port map (
            O => \N__30046\,
            I => \N__30007\
        );

    \I__6217\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30007\
        );

    \I__6216\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30002\
        );

    \I__6215\ : InMux
    port map (
            O => \N__30039\,
            I => \N__30002\
        );

    \I__6214\ : InMux
    port map (
            O => \N__30036\,
            I => \N__29995\
        );

    \I__6213\ : InMux
    port map (
            O => \N__30033\,
            I => \N__29995\
        );

    \I__6212\ : InMux
    port map (
            O => \N__30032\,
            I => \N__29995\
        );

    \I__6211\ : CascadeMux
    port map (
            O => \N__30031\,
            I => \N__29990\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__30030\,
            I => \N__29987\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__30027\,
            I => \N__29984\
        );

    \I__6208\ : InMux
    port map (
            O => \N__30026\,
            I => \N__29981\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__30025\,
            I => \N__29977\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__30024\,
            I => \N__29974\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__30023\,
            I => \N__29971\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__30022\,
            I => \N__29968\
        );

    \I__6203\ : InMux
    port map (
            O => \N__30021\,
            I => \N__29963\
        );

    \I__6202\ : InMux
    port map (
            O => \N__30018\,
            I => \N__29960\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__29957\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__29951\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__30013\,
            I => \N__29948\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__30012\,
            I => \N__29945\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__30007\,
            I => \N__29942\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29937\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__29995\,
            I => \N__29937\
        );

    \I__6194\ : CascadeMux
    port map (
            O => \N__29994\,
            I => \N__29934\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__29993\,
            I => \N__29931\
        );

    \I__6192\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29926\
        );

    \I__6191\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29926\
        );

    \I__6190\ : Span4Mux_v
    port map (
            O => \N__29984\,
            I => \N__29921\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__29981\,
            I => \N__29921\
        );

    \I__6188\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29918\
        );

    \I__6187\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29915\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29911\
        );

    \I__6185\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29908\
        );

    \I__6184\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29905\
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__29967\,
            I => \N__29902\
        );

    \I__6182\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29899\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__29963\,
            I => \N__29891\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__29960\,
            I => \N__29891\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__29957\,
            I => \N__29891\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__29956\,
            I => \N__29888\
        );

    \I__6177\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29883\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29883\
        );

    \I__6175\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29880\
        );

    \I__6174\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29875\
        );

    \I__6173\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29875\
        );

    \I__6172\ : Span4Mux_h
    port map (
            O => \N__29942\,
            I => \N__29870\
        );

    \I__6171\ : Span4Mux_v
    port map (
            O => \N__29937\,
            I => \N__29870\
        );

    \I__6170\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29865\
        );

    \I__6169\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29865\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__29926\,
            I => \N__29860\
        );

    \I__6167\ : Span4Mux_v
    port map (
            O => \N__29921\,
            I => \N__29860\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__29918\,
            I => \N__29857\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__29915\,
            I => \N__29854\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__29914\,
            I => \N__29851\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29844\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__29908\,
            I => \N__29844\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__29905\,
            I => \N__29844\
        );

    \I__6160\ : InMux
    port map (
            O => \N__29902\,
            I => \N__29841\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__29899\,
            I => \N__29838\
        );

    \I__6158\ : CascadeMux
    port map (
            O => \N__29898\,
            I => \N__29833\
        );

    \I__6157\ : Span4Mux_h
    port map (
            O => \N__29891\,
            I => \N__29830\
        );

    \I__6156\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29827\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29818\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29818\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__29875\,
            I => \N__29818\
        );

    \I__6152\ : Span4Mux_v
    port map (
            O => \N__29870\,
            I => \N__29818\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__29865\,
            I => \N__29815\
        );

    \I__6150\ : Span4Mux_h
    port map (
            O => \N__29860\,
            I => \N__29810\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__29857\,
            I => \N__29810\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__29854\,
            I => \N__29807\
        );

    \I__6147\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29804\
        );

    \I__6146\ : Span4Mux_v
    port map (
            O => \N__29844\,
            I => \N__29801\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__29841\,
            I => \N__29798\
        );

    \I__6144\ : Span12Mux_v
    port map (
            O => \N__29838\,
            I => \N__29795\
        );

    \I__6143\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29788\
        );

    \I__6142\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29788\
        );

    \I__6141\ : InMux
    port map (
            O => \N__29833\,
            I => \N__29788\
        );

    \I__6140\ : Span4Mux_v
    port map (
            O => \N__29830\,
            I => \N__29785\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__29827\,
            I => \N__29780\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__29818\,
            I => \N__29780\
        );

    \I__6137\ : Span4Mux_v
    port map (
            O => \N__29815\,
            I => \N__29773\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__29810\,
            I => \N__29773\
        );

    \I__6135\ : Span4Mux_h
    port map (
            O => \N__29807\,
            I => \N__29773\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__29804\,
            I => \aluReadBus_rep2\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__29801\,
            I => \aluReadBus_rep2\
        );

    \I__6132\ : Odrv12
    port map (
            O => \N__29798\,
            I => \aluReadBus_rep2\
        );

    \I__6131\ : Odrv12
    port map (
            O => \N__29795\,
            I => \aluReadBus_rep2\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__29788\,
            I => \aluReadBus_rep2\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__29785\,
            I => \aluReadBus_rep2\
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__29780\,
            I => \aluReadBus_rep2\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__29773\,
            I => \aluReadBus_rep2\
        );

    \I__6126\ : CascadeMux
    port map (
            O => \N__29756\,
            I => \N__29750\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__29755\,
            I => \N__29747\
        );

    \I__6124\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29742\
        );

    \I__6123\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29736\
        );

    \I__6122\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29730\
        );

    \I__6121\ : InMux
    port map (
            O => \N__29747\,
            I => \N__29730\
        );

    \I__6120\ : InMux
    port map (
            O => \N__29746\,
            I => \N__29723\
        );

    \I__6119\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29723\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__29742\,
            I => \N__29720\
        );

    \I__6117\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29717\
        );

    \I__6116\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29714\
        );

    \I__6115\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29711\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__29736\,
            I => \N__29708\
        );

    \I__6113\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29705\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29698\
        );

    \I__6111\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29693\
        );

    \I__6110\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29693\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29688\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__29720\,
            I => \N__29683\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__29717\,
            I => \N__29683\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29673\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29673\
        );

    \I__6104\ : Span4Mux_v
    port map (
            O => \N__29708\,
            I => \N__29668\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29668\
        );

    \I__6102\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29659\
        );

    \I__6101\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29659\
        );

    \I__6100\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29659\
        );

    \I__6099\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29659\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__29698\,
            I => \N__29654\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29654\
        );

    \I__6096\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29649\
        );

    \I__6095\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29649\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__29688\,
            I => \N__29644\
        );

    \I__6093\ : Span4Mux_h
    port map (
            O => \N__29683\,
            I => \N__29644\
        );

    \I__6092\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29639\
        );

    \I__6091\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29639\
        );

    \I__6090\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29632\
        );

    \I__6089\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29632\
        );

    \I__6088\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29632\
        );

    \I__6087\ : Span4Mux_h
    port map (
            O => \N__29673\,
            I => \N__29623\
        );

    \I__6086\ : Span4Mux_v
    port map (
            O => \N__29668\,
            I => \N__29623\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__29659\,
            I => \N__29623\
        );

    \I__6084\ : Span4Mux_h
    port map (
            O => \N__29654\,
            I => \N__29623\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__29649\,
            I => \busState_0\
        );

    \I__6082\ : Odrv4
    port map (
            O => \N__29644\,
            I => \busState_0\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__29639\,
            I => \busState_0\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__29632\,
            I => \busState_0\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__29623\,
            I => \busState_0\
        );

    \I__6078\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29609\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29606\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__29606\,
            I => \N__29603\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__29603\,
            I => \ALU.N_9_1\
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__29600\,
            I => \FTDI.N_217_0_cascade_\
        );

    \I__6073\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29594\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__29594\,
            I => \FTDI.N_216_0\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__29591\,
            I => \FTDI.TXready_cascade_\
        );

    \I__6070\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29583\
        );

    \I__6069\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29580\
        );

    \I__6068\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29577\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__29583\,
            I => \FTDI.baudAccZ0Z_0\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__29580\,
            I => \FTDI.baudAccZ0Z_0\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__29577\,
            I => \FTDI.baudAccZ0Z_0\
        );

    \I__6064\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29564\
        );

    \I__6062\ : Span4Mux_h
    port map (
            O => \N__29564\,
            I => \N__29560\
        );

    \I__6061\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29557\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__29560\,
            I => \FTDI.baudAccZ0Z_1\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__29557\,
            I => \FTDI.baudAccZ0Z_1\
        );

    \I__6058\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__29549\,
            I => \N__29546\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__29546\,
            I => \N__29543\
        );

    \I__6055\ : Span4Mux_h
    port map (
            O => \N__29543\,
            I => \N__29540\
        );

    \I__6054\ : Span4Mux_h
    port map (
            O => \N__29540\,
            I => \N__29537\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__29537\,
            I => \ALU.N_290_0\
        );

    \I__6052\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29531\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__29531\,
            I => \ALU.rshift_5\
        );

    \I__6050\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29525\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__29525\,
            I => \ALU.a_15_m3_5\
        );

    \I__6048\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29514\
        );

    \I__6047\ : InMux
    port map (
            O => \N__29521\,
            I => \N__29507\
        );

    \I__6046\ : InMux
    port map (
            O => \N__29520\,
            I => \N__29507\
        );

    \I__6045\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29507\
        );

    \I__6044\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29502\
        );

    \I__6043\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29502\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__29514\,
            I => \FTDI.TXstateZ1Z_0\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__29507\,
            I => \FTDI.TXstateZ1Z_0\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__29502\,
            I => \FTDI.TXstateZ1Z_0\
        );

    \I__6039\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29483\
        );

    \I__6038\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29483\
        );

    \I__6037\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29483\
        );

    \I__6036\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29480\
        );

    \I__6035\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29475\
        );

    \I__6034\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29475\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__29483\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__29480\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__29475\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__6030\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29464\
        );

    \I__6029\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29461\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__29464\,
            I => \FTDI.N_170_0\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__29461\,
            I => \FTDI.N_170_0\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__29456\,
            I => \FTDI.TXstate_e_1_3_cascade_\
        );

    \I__6025\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29450\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29447\
        );

    \I__6023\ : Span4Mux_h
    port map (
            O => \N__29447\,
            I => \N__29444\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__29444\,
            I => \N__29441\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__29441\,
            I => \ALU.N_11_0\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__29438\,
            I => \N__29430\
        );

    \I__6019\ : InMux
    port map (
            O => \N__29437\,
            I => \N__29427\
        );

    \I__6018\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29423\
        );

    \I__6017\ : InMux
    port map (
            O => \N__29435\,
            I => \N__29420\
        );

    \I__6016\ : CascadeMux
    port map (
            O => \N__29434\,
            I => \N__29417\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__29433\,
            I => \N__29414\
        );

    \I__6014\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29409\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29406\
        );

    \I__6012\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29399\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29394\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29394\
        );

    \I__6009\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29387\
        );

    \I__6008\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29387\
        );

    \I__6007\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29387\
        );

    \I__6006\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29384\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29381\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__29406\,
            I => \N__29374\
        );

    \I__6003\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29371\
        );

    \I__6002\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29368\
        );

    \I__6001\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29362\
        );

    \I__6000\ : InMux
    port map (
            O => \N__29402\,
            I => \N__29362\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__29399\,
            I => \N__29355\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__29394\,
            I => \N__29355\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__29387\,
            I => \N__29355\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__29384\,
            I => \N__29352\
        );

    \I__5995\ : Span4Mux_h
    port map (
            O => \N__29381\,
            I => \N__29349\
        );

    \I__5994\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29342\
        );

    \I__5993\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29342\
        );

    \I__5992\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29342\
        );

    \I__5991\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29339\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__29374\,
            I => \N__29334\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__29371\,
            I => \N__29334\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__29368\,
            I => \N__29331\
        );

    \I__5987\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29328\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29325\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__29355\,
            I => \N__29316\
        );

    \I__5984\ : Span4Mux_h
    port map (
            O => \N__29352\,
            I => \N__29316\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__29349\,
            I => \N__29316\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__29342\,
            I => \N__29316\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29311\
        );

    \I__5980\ : Span4Mux_h
    port map (
            O => \N__29334\,
            I => \N__29311\
        );

    \I__5979\ : Span4Mux_v
    port map (
            O => \N__29331\,
            I => \N__29306\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__29328\,
            I => \N__29299\
        );

    \I__5977\ : Span4Mux_v
    port map (
            O => \N__29325\,
            I => \N__29299\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__29316\,
            I => \N__29299\
        );

    \I__5975\ : Sp12to4
    port map (
            O => \N__29311\,
            I => \N__29296\
        );

    \I__5974\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29293\
        );

    \I__5973\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29289\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__29306\,
            I => \N__29284\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__29299\,
            I => \N__29284\
        );

    \I__5970\ : Span12Mux_s6_v
    port map (
            O => \N__29296\,
            I => \N__29279\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__29293\,
            I => \N__29279\
        );

    \I__5968\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29276\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__29289\,
            I => \ALU.N_5_0\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__29284\,
            I => \ALU.N_5_0\
        );

    \I__5965\ : Odrv12
    port map (
            O => \N__29279\,
            I => \ALU.N_5_0\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__29276\,
            I => \ALU.N_5_0\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__29267\,
            I => \N__29263\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__29266\,
            I => \N__29258\
        );

    \I__5961\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29251\
        );

    \I__5960\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29251\
        );

    \I__5959\ : InMux
    port map (
            O => \N__29261\,
            I => \N__29251\
        );

    \I__5958\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29246\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29243\
        );

    \I__5956\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29238\
        );

    \I__5955\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29238\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29235\
        );

    \I__5953\ : Span4Mux_v
    port map (
            O => \N__29243\,
            I => \N__29230\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__29238\,
            I => \N__29230\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__29235\,
            I => \N__29227\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__29230\,
            I => \N__29224\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__29227\,
            I => \FTDI.gapZ0Z_2\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__29224\,
            I => \FTDI.gapZ0Z_2\
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__29219\,
            I => \N__29216\
        );

    \I__5946\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29210\
        );

    \I__5945\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29210\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29207\
        );

    \I__5943\ : Span4Mux_s1_v
    port map (
            O => \N__29207\,
            I => \N__29203\
        );

    \I__5942\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29200\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__29203\,
            I => \FTDI.gapZ0Z_0\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__29200\,
            I => \FTDI.gapZ0Z_0\
        );

    \I__5939\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29190\
        );

    \I__5938\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29185\
        );

    \I__5937\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29185\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__29190\,
            I => \N__29182\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29179\
        );

    \I__5934\ : IoSpan4Mux
    port map (
            O => \N__29182\,
            I => \N__29176\
        );

    \I__5933\ : Span4Mux_h
    port map (
            O => \N__29179\,
            I => \N__29171\
        );

    \I__5932\ : Span4Mux_s0_v
    port map (
            O => \N__29176\,
            I => \N__29171\
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__29171\,
            I => \FTDI.gap8\
        );

    \I__5930\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29162\
        );

    \I__5929\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29162\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__29162\,
            I => \FTDI.gapZ0Z_1\
        );

    \I__5927\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29156\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__29156\,
            I => \FTDI.TXstate_e_1_0\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__29153\,
            I => \FTDI.N_169_0_cascade_\
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__5923\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__29144\,
            I => \FTDI.N_169_0\
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__29141\,
            I => \FTDI.TXstate_cnst_0_0_2_cascade_\
        );

    \I__5920\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29135\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__29135\,
            I => \N__29131\
        );

    \I__5918\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29128\
        );

    \I__5917\ : Span4Mux_h
    port map (
            O => \N__29131\,
            I => \N__29125\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__29128\,
            I => \N__29122\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__29125\,
            I => \ALU.cZ0Z_0\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__29122\,
            I => \ALU.cZ0Z_0\
        );

    \I__5913\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29114\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29111\
        );

    \I__5911\ : Span4Mux_v
    port map (
            O => \N__29111\,
            I => \N__29107\
        );

    \I__5910\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29104\
        );

    \I__5909\ : Span4Mux_h
    port map (
            O => \N__29107\,
            I => \N__29101\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__29104\,
            I => \ALU.cZ0Z_1\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__29101\,
            I => \ALU.cZ0Z_1\
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__29096\,
            I => \N__29093\
        );

    \I__5905\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__29090\,
            I => \N__29086\
        );

    \I__5903\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29083\
        );

    \I__5902\ : Span4Mux_v
    port map (
            O => \N__29086\,
            I => \N__29080\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29077\
        );

    \I__5900\ : Odrv4
    port map (
            O => \N__29080\,
            I => \ALU.cZ0Z_2\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__29077\,
            I => \ALU.cZ0Z_2\
        );

    \I__5898\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29068\
        );

    \I__5897\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29062\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29059\
        );

    \I__5894\ : Span4Mux_h
    port map (
            O => \N__29062\,
            I => \N__29056\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__29059\,
            I => \ALU.cZ0Z_3\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__29056\,
            I => \ALU.cZ0Z_3\
        );

    \I__5891\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29048\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__29048\,
            I => \N__29044\
        );

    \I__5889\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29041\
        );

    \I__5888\ : Span4Mux_v
    port map (
            O => \N__29044\,
            I => \N__29036\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__29041\,
            I => \N__29036\
        );

    \I__5886\ : Span4Mux_h
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__29033\,
            I => \ALU.cZ0Z_4\
        );

    \I__5884\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29027\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__29027\,
            I => \N__29023\
        );

    \I__5882\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29020\
        );

    \I__5881\ : Odrv12
    port map (
            O => \N__29023\,
            I => \ALU.cZ0Z_5\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__29020\,
            I => \ALU.cZ0Z_5\
        );

    \I__5879\ : InMux
    port map (
            O => \N__29015\,
            I => \N__29012\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__29012\,
            I => \N__29008\
        );

    \I__5877\ : InMux
    port map (
            O => \N__29011\,
            I => \N__29005\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__29008\,
            I => \N__29002\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__29005\,
            I => \ALU.cZ0Z_6\
        );

    \I__5874\ : Odrv4
    port map (
            O => \N__29002\,
            I => \ALU.cZ0Z_6\
        );

    \I__5873\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28994\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__5871\ : Span4Mux_h
    port map (
            O => \N__28991\,
            I => \N__28987\
        );

    \I__5870\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28984\
        );

    \I__5869\ : Span4Mux_v
    port map (
            O => \N__28987\,
            I => \N__28979\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__28984\,
            I => \N__28979\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__28979\,
            I => \ALU.dZ0Z_4\
        );

    \I__5866\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28972\
        );

    \I__5865\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28969\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28966\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__28969\,
            I => \N__28963\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__28966\,
            I => \N__28960\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__28963\,
            I => \N__28957\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__28960\,
            I => \ALU.gZ0Z_6\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__28957\,
            I => \ALU.gZ0Z_6\
        );

    \I__5858\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28949\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__28949\,
            I => \N__28945\
        );

    \I__5856\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28942\
        );

    \I__5855\ : Odrv12
    port map (
            O => \N__28945\,
            I => \ALU.eZ0Z_0\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__28942\,
            I => \ALU.eZ0Z_0\
        );

    \I__5853\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28930\
        );

    \I__5851\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28927\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__28930\,
            I => \N__28923\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28920\
        );

    \I__5848\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28917\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__28923\,
            I => \N__28914\
        );

    \I__5846\ : Span4Mux_v
    port map (
            O => \N__28920\,
            I => \N__28909\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__28917\,
            I => \N__28909\
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__28914\,
            I => a_0
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__28909\,
            I => a_0
        );

    \I__5842\ : CascadeMux
    port map (
            O => \N__28904\,
            I => \N__28901\
        );

    \I__5841\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28898\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__28898\,
            I => \N__28895\
        );

    \I__5839\ : Odrv12
    port map (
            O => \N__28895\,
            I => \ALU.e_RNINIVJZ0Z_0\
        );

    \I__5838\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28889\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__28889\,
            I => \ALU.g_RNIM8LLZ0Z_5\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__28886\,
            I => \ALU.e_RNI1TVJZ0Z_5_cascade_\
        );

    \I__5835\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28880\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__28880\,
            I => \N__28877\
        );

    \I__5833\ : Span4Mux_v
    port map (
            O => \N__28877\,
            I => \N__28874\
        );

    \I__5832\ : Span4Mux_h
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__28871\,
            I => \ALU.operand2_7_ns_1_5\
        );

    \I__5830\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28865\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__28865\,
            I => \N__28862\
        );

    \I__5828\ : Span4Mux_h
    port map (
            O => \N__28862\,
            I => \N__28858\
        );

    \I__5827\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28855\
        );

    \I__5826\ : Odrv4
    port map (
            O => \N__28858\,
            I => \ALU.eZ0Z_5\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__28855\,
            I => \ALU.eZ0Z_5\
        );

    \I__5824\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28847\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__28841\,
            I => \ALU.g_RNIRUBOZ0Z_0\
        );

    \I__5820\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28835\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28832\
        );

    \I__5818\ : Span4Mux_h
    port map (
            O => \N__28832\,
            I => \N__28829\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__28829\,
            I => \ALU.d_RNIG6R7Z0Z_1\
        );

    \I__5816\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28820\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__28820\,
            I => \N__28817\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__28814\,
            I => \ALU.d_RNI45J9Z0Z_1\
        );

    \I__5811\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28808\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__28808\,
            I => \ALU.d_RNII8R7Z0Z_2\
        );

    \I__5809\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28802\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__5807\ : Span4Mux_h
    port map (
            O => \N__28799\,
            I => \N__28795\
        );

    \I__5806\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28792\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__28795\,
            I => \N__28789\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28786\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__28789\,
            I => \ALU.eZ0Z_7\
        );

    \I__5802\ : Odrv12
    port map (
            O => \N__28786\,
            I => \ALU.eZ0Z_7\
        );

    \I__5801\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28777\
        );

    \I__5800\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28774\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__28777\,
            I => \ALU.eZ0Z_2\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__28774\,
            I => \ALU.eZ0Z_2\
        );

    \I__5797\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__28763\,
            I => \N__28760\
        );

    \I__5794\ : Span4Mux_v
    port map (
            O => \N__28760\,
            I => \N__28755\
        );

    \I__5793\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28752\
        );

    \I__5792\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28749\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__28755\,
            I => a_2
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__28752\,
            I => a_2
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__28749\,
            I => a_2
        );

    \I__5788\ : CascadeMux
    port map (
            O => \N__28742\,
            I => \ALU.g_RNIV2COZ0Z_2_cascade_\
        );

    \I__5787\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28736\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__28736\,
            I => \ALU.e_RNIRMVJZ0Z_2\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__28733\,
            I => \ALU.operand2_7_ns_1_2_cascade_\
        );

    \I__5784\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28727\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28723\
        );

    \I__5782\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28720\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__28723\,
            I => \N__28717\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__28720\,
            I => \N__28714\
        );

    \I__5779\ : Span4Mux_h
    port map (
            O => \N__28717\,
            I => \N__28711\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__28714\,
            I => \N__28708\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__28711\,
            I => \N__28703\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__28708\,
            I => \N__28703\
        );

    \I__5775\ : Odrv4
    port map (
            O => \N__28703\,
            I => \ALU.operand2_2\
        );

    \I__5774\ : InMux
    port map (
            O => \N__28700\,
            I => \N__28697\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__28697\,
            I => \N__28694\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__28694\,
            I => \N__28691\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__28691\,
            I => \ALU.un2_addsub_cry_12_c_RNIUL1GKZ0\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__28688\,
            I => \un2_addsub_cry_12_c_RNIG3PMU_cascade_\
        );

    \I__5769\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28682\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28679\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__5765\ : Odrv4
    port map (
            O => \N__28673\,
            I => \c_RNI88B4N2_13\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__28670\,
            I => \aluOperation_RNI2J9SL3_0_cascade_\
        );

    \I__5763\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28664\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__28664\,
            I => \N__28661\
        );

    \I__5761\ : Span4Mux_v
    port map (
            O => \N__28661\,
            I => \N__28658\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__28658\,
            I => \ALU.mult_2\
        );

    \I__5759\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__28652\,
            I => \N__28649\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__28649\,
            I => \N__28646\
        );

    \I__5756\ : Span4Mux_v
    port map (
            O => \N__28646\,
            I => \N__28643\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__28643\,
            I => \ALU.a_15_m5_2\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__28640\,
            I => \ALU.d_RNIIFMN04Z0Z_2_cascade_\
        );

    \I__5753\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28631\
        );

    \I__5752\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28631\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__28631\,
            I => \N__28628\
        );

    \I__5750\ : Span4Mux_h
    port map (
            O => \N__28628\,
            I => \N__28625\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__28625\,
            I => \ALU.eZ0Z_3\
        );

    \I__5748\ : InMux
    port map (
            O => \N__28622\,
            I => \N__28618\
        );

    \I__5747\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28615\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28612\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__28615\,
            I => \N__28609\
        );

    \I__5744\ : Span4Mux_h
    port map (
            O => \N__28612\,
            I => \N__28606\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__28609\,
            I => \ALU.eZ0Z_6\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__28606\,
            I => \ALU.eZ0Z_6\
        );

    \I__5741\ : InMux
    port map (
            O => \N__28601\,
            I => \N__28597\
        );

    \I__5740\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28594\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__28597\,
            I => \N__28590\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__28594\,
            I => \N__28587\
        );

    \I__5737\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28584\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__28590\,
            I => \N__28581\
        );

    \I__5735\ : Span4Mux_v
    port map (
            O => \N__28587\,
            I => \N__28576\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28576\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__28581\,
            I => \N__28573\
        );

    \I__5732\ : Span4Mux_h
    port map (
            O => \N__28576\,
            I => \N__28570\
        );

    \I__5731\ : Odrv4
    port map (
            O => \N__28573\,
            I => \ALU.eZ0Z_10\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__28570\,
            I => \ALU.eZ0Z_10\
        );

    \I__5729\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28562\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__28562\,
            I => \N__28558\
        );

    \I__5727\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28555\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__28558\,
            I => \N__28552\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__28555\,
            I => \N__28549\
        );

    \I__5724\ : Span4Mux_h
    port map (
            O => \N__28552\,
            I => \N__28544\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__28549\,
            I => \N__28544\
        );

    \I__5722\ : Odrv4
    port map (
            O => \N__28544\,
            I => \ALU.eZ0Z_12\
        );

    \I__5721\ : InMux
    port map (
            O => \N__28541\,
            I => \N__28538\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__28535\,
            I => \N__28532\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__28532\,
            I => \N__28529\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__28529\,
            I => \ALU.d_RNIPER7Z0Z_5\
        );

    \I__5716\ : InMux
    port map (
            O => \N__28526\,
            I => \N__28522\
        );

    \I__5715\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28519\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28515\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28512\
        );

    \I__5712\ : InMux
    port map (
            O => \N__28518\,
            I => \N__28509\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__28515\,
            I => \N__28506\
        );

    \I__5710\ : Span4Mux_h
    port map (
            O => \N__28512\,
            I => \N__28503\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__28509\,
            I => \ALU.bZ0Z_10\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__28506\,
            I => \ALU.bZ0Z_10\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__28503\,
            I => \ALU.bZ0Z_10\
        );

    \I__5706\ : InMux
    port map (
            O => \N__28496\,
            I => \N__28492\
        );

    \I__5705\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28489\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28484\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__28489\,
            I => \N__28484\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__28481\,
            I => \N__28478\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__28478\,
            I => \ALU.bZ0Z_15\
        );

    \I__5699\ : InMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__5697\ : Span4Mux_h
    port map (
            O => \N__28469\,
            I => \N__28465\
        );

    \I__5696\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28462\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__28465\,
            I => \ALU.fZ0Z_11\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__28462\,
            I => \ALU.fZ0Z_11\
        );

    \I__5693\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28454\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__28454\,
            I => \N__28451\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__28451\,
            I => \N__28447\
        );

    \I__5690\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28444\
        );

    \I__5689\ : Odrv4
    port map (
            O => \N__28447\,
            I => \ALU.bZ0Z_11\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__28444\,
            I => \ALU.bZ0Z_11\
        );

    \I__5687\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28436\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__28430\,
            I => \ALU.b_RNIKNSD1Z0Z_13\
        );

    \I__5683\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28423\
        );

    \I__5682\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28419\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28416\
        );

    \I__5680\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28413\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__28419\,
            I => \N__28408\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__28416\,
            I => \N__28408\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__28413\,
            I => \N__28405\
        );

    \I__5676\ : Span4Mux_v
    port map (
            O => \N__28408\,
            I => \N__28402\
        );

    \I__5675\ : Span4Mux_h
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__28402\,
            I => \ALU.dZ0Z_10\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__28399\,
            I => \ALU.dZ0Z_10\
        );

    \I__5672\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28391\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__28391\,
            I => \N__28387\
        );

    \I__5670\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28384\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__28387\,
            I => \N__28381\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__5667\ : Span4Mux_h
    port map (
            O => \N__28381\,
            I => \N__28373\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__28378\,
            I => \N__28373\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__28373\,
            I => \ALU.dZ0Z_12\
        );

    \I__5664\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28367\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__28367\,
            I => \N__28364\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__28364\,
            I => \N__28360\
        );

    \I__5661\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28357\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__28360\,
            I => \N__28354\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__28357\,
            I => \ALU.bZ0Z_12\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__28354\,
            I => \ALU.bZ0Z_12\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__28349\,
            I => \N__28346\
        );

    \I__5656\ : InMux
    port map (
            O => \N__28346\,
            I => \N__28343\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__28343\,
            I => \N__28339\
        );

    \I__5654\ : InMux
    port map (
            O => \N__28342\,
            I => \N__28336\
        );

    \I__5653\ : Span12Mux_s8_h
    port map (
            O => \N__28339\,
            I => \N__28333\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__28336\,
            I => \ALU.fZ0Z_12\
        );

    \I__5651\ : Odrv12
    port map (
            O => \N__28333\,
            I => \ALU.fZ0Z_12\
        );

    \I__5650\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__28325\,
            I => \ALU.b_RNIILSD1Z0Z_12\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__28322\,
            I => \N__28319\
        );

    \I__5647\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28316\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__28313\,
            I => \N__28310\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__28310\,
            I => \N__28306\
        );

    \I__5643\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28303\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__28306\,
            I => \ALU.fZ0Z_14\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__28303\,
            I => \ALU.fZ0Z_14\
        );

    \I__5640\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__28292\,
            I => \N__28289\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__28289\,
            I => \N__28285\
        );

    \I__5636\ : InMux
    port map (
            O => \N__28288\,
            I => \N__28282\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__28285\,
            I => \ALU.bZ0Z_14\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__28282\,
            I => \ALU.bZ0Z_14\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__28277\,
            I => \ALU.g0_3_1_cascade_\
        );

    \I__5632\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__28271\,
            I => \N__28268\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__28265\,
            I => \N__28262\
        );

    \I__5628\ : Span4Mux_h
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__28259\,
            I => \ALU.N_703_0_0\
        );

    \I__5626\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28253\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__28253\,
            I => \ALU.N_4\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__28250\,
            I => \N__28247\
        );

    \I__5623\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28244\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__28244\,
            I => \N__28241\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__28241\,
            I => \ALU.N_5\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__28238\,
            I => \ALU.a_15_m4_12_cascade_\
        );

    \I__5619\ : InMux
    port map (
            O => \N__28235\,
            I => \N__28232\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__28232\,
            I => \N__28229\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__28226\,
            I => \ALU.un2_addsub_cry_11_c_RNII7OFZ0Z9\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__28223\,
            I => \un2_addsub_cry_11_c_RNIQ9LMU_cascade_\
        );

    \I__5614\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28217\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__28217\,
            I => \c_RNIC8RDN2_12\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__28214\,
            I => \aluOperation_RNIGPL5M3_0_cascade_\
        );

    \I__5611\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28208\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__28208\,
            I => \N__28204\
        );

    \I__5609\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28201\
        );

    \I__5608\ : Odrv12
    port map (
            O => \N__28204\,
            I => \ALU.aZ0Z_12\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__28201\,
            I => \ALU.aZ0Z_12\
        );

    \I__5606\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28193\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__5604\ : Odrv12
    port map (
            O => \N__28190\,
            I => \ALU.N_271_0\
        );

    \I__5603\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__28184\,
            I => \ALU.a_15_m3_12\
        );

    \I__5601\ : InMux
    port map (
            O => \N__28181\,
            I => \N__28178\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__5599\ : Span4Mux_v
    port map (
            O => \N__28175\,
            I => \N__28172\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__28169\,
            I => \ALU.N_314\
        );

    \I__5596\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28163\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__28163\,
            I => \ALU.lshift_12\
        );

    \I__5594\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28155\
        );

    \I__5593\ : CascadeMux
    port map (
            O => \N__28159\,
            I => \N__28152\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__28158\,
            I => \N__28149\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__28155\,
            I => \N__28146\
        );

    \I__5590\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28141\
        );

    \I__5589\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28141\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__28146\,
            I => \N__28138\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__28141\,
            I => \ALU.fZ0Z_9\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__28138\,
            I => \ALU.fZ0Z_9\
        );

    \I__5585\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28130\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__28130\,
            I => \N__28127\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__28127\,
            I => \N__28122\
        );

    \I__5582\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28117\
        );

    \I__5581\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28117\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__28122\,
            I => \N__28114\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__28117\,
            I => \ALU.bZ0Z_9\
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__28114\,
            I => \ALU.bZ0Z_9\
        );

    \I__5577\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28106\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__28106\,
            I => \N__28103\
        );

    \I__5575\ : Odrv12
    port map (
            O => \N__28103\,
            I => \ALU.f_RNIUUJ01Z0Z_9\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__28100\,
            I => \ALU.a_15_m2_ns_1Z0Z_5_cascade_\
        );

    \I__5573\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__5571\ : Span4Mux_v
    port map (
            O => \N__28091\,
            I => \N__28081\
        );

    \I__5570\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28078\
        );

    \I__5569\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28075\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__28088\,
            I => \N__28072\
        );

    \I__5567\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28065\
        );

    \I__5566\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28060\
        );

    \I__5565\ : InMux
    port map (
            O => \N__28085\,
            I => \N__28060\
        );

    \I__5564\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28057\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__28081\,
            I => \N__28050\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__28078\,
            I => \N__28050\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__28075\,
            I => \N__28050\
        );

    \I__5560\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28047\
        );

    \I__5559\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28044\
        );

    \I__5558\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28041\
        );

    \I__5557\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28036\
        );

    \I__5556\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28036\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__28065\,
            I => \N__28031\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28028\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28020\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__28050\,
            I => \N__28020\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__28047\,
            I => \N__28015\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__28044\,
            I => \N__28015\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__28041\,
            I => \N__28010\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__28010\
        );

    \I__5547\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28007\
        );

    \I__5546\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28004\
        );

    \I__5545\ : Span4Mux_v
    port map (
            O => \N__28031\,
            I => \N__27999\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__28028\,
            I => \N__27999\
        );

    \I__5543\ : InMux
    port map (
            O => \N__28027\,
            I => \N__27996\
        );

    \I__5542\ : InMux
    port map (
            O => \N__28026\,
            I => \N__27991\
        );

    \I__5541\ : InMux
    port map (
            O => \N__28025\,
            I => \N__27991\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__28020\,
            I => \N__27988\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__28015\,
            I => \N__27983\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__27983\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__28007\,
            I => \ALU.N_225_0\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__28004\,
            I => \ALU.N_225_0\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__27999\,
            I => \ALU.N_225_0\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__27996\,
            I => \ALU.N_225_0\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__27991\,
            I => \ALU.N_225_0\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__27988\,
            I => \ALU.N_225_0\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__27983\,
            I => \ALU.N_225_0\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__27968\,
            I => \ALU.a_15_m2_5_cascade_\
        );

    \I__5529\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__27959\,
            I => \N__27955\
        );

    \I__5526\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27952\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__27955\,
            I => \ALU.N_420\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__27952\,
            I => \ALU.N_420\
        );

    \I__5523\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27944\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__27944\,
            I => \ALU.a_15_m4_5\
        );

    \I__5521\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27937\
        );

    \I__5520\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27934\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27931\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__27934\,
            I => \N__27928\
        );

    \I__5517\ : Span4Mux_h
    port map (
            O => \N__27931\,
            I => \N__27925\
        );

    \I__5516\ : Span12Mux_h
    port map (
            O => \N__27928\,
            I => \N__27921\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__27925\,
            I => \N__27918\
        );

    \I__5514\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27915\
        );

    \I__5513\ : Odrv12
    port map (
            O => \N__27921\,
            I => a_4
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__27918\,
            I => a_4
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__27915\,
            I => a_4
        );

    \I__5510\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27905\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__27905\,
            I => \N__27902\
        );

    \I__5508\ : Span4Mux_v
    port map (
            O => \N__27902\,
            I => \N__27899\
        );

    \I__5507\ : Sp12to4
    port map (
            O => \N__27899\,
            I => \N__27894\
        );

    \I__5506\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27891\
        );

    \I__5505\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27888\
        );

    \I__5504\ : Span12Mux_s8_h
    port map (
            O => \N__27894\,
            I => \N__27883\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__27891\,
            I => \N__27883\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__27888\,
            I => \N__27880\
        );

    \I__5501\ : Odrv12
    port map (
            O => \N__27883\,
            I => a_6
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__27880\,
            I => a_6
        );

    \I__5499\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27871\
        );

    \I__5498\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27867\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__27871\,
            I => \N__27864\
        );

    \I__5496\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27861\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__27867\,
            I => \N__27858\
        );

    \I__5494\ : Span4Mux_h
    port map (
            O => \N__27864\,
            I => \N__27855\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__27861\,
            I => \N__27852\
        );

    \I__5492\ : Span12Mux_v
    port map (
            O => \N__27858\,
            I => \N__27849\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__27855\,
            I => \N__27846\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__27852\,
            I => \N__27843\
        );

    \I__5489\ : Odrv12
    port map (
            O => \N__27849\,
            I => a_7
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__27846\,
            I => a_7
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__27843\,
            I => a_7
        );

    \I__5486\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27833\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__27833\,
            I => \N__27830\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__27830\,
            I => \ALU.a_15_m2_12\
        );

    \I__5483\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27824\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__27824\,
            I => \ALU.rshift_15_ns_1_7\
        );

    \I__5481\ : CascadeMux
    port map (
            O => \N__27821\,
            I => \ALU.rshift_3_ns_1_3_cascade_\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__27818\,
            I => \ALU.N_471_cascade_\
        );

    \I__5479\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__27812\,
            I => \ALU.N_475\
        );

    \I__5477\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27806\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__27806\,
            I => \ALU.rshift_3_ns_1_7\
        );

    \I__5475\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27797\
        );

    \I__5474\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27797\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__27797\,
            I => \ALU.N_576\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__27794\,
            I => \ALU.a_15_m5_5_cascade_\
        );

    \I__5471\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27788\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__27788\,
            I => \N__27785\
        );

    \I__5469\ : Span4Mux_h
    port map (
            O => \N__27785\,
            I => \N__27782\
        );

    \I__5468\ : Span4Mux_v
    port map (
            O => \N__27782\,
            I => \N__27779\
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__27779\,
            I => \ALU.mult_5\
        );

    \I__5466\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27773\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__27773\,
            I => \N__27770\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__27770\,
            I => \ALU.d_RNIPFIBI1Z0Z_9\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__27767\,
            I => \ALU.dout_3_ns_1_6_cascade_\
        );

    \I__5462\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27761\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__27761\,
            I => \ALU.N_705\
        );

    \I__5460\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27752\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__27752\,
            I => \N__27749\
        );

    \I__5457\ : Span4Mux_v
    port map (
            O => \N__27749\,
            I => \N__27746\
        );

    \I__5456\ : Span4Mux_v
    port map (
            O => \N__27746\,
            I => \N__27742\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__27745\,
            I => \N__27739\
        );

    \I__5454\ : Sp12to4
    port map (
            O => \N__27742\,
            I => \N__27736\
        );

    \I__5453\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27733\
        );

    \I__5452\ : Odrv12
    port map (
            O => \N__27736\,
            I => \testWordZ0Z_7\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__27733\,
            I => \testWordZ0Z_7\
        );

    \I__5450\ : CEMux
    port map (
            O => \N__27728\,
            I => \N__27724\
        );

    \I__5449\ : CEMux
    port map (
            O => \N__27727\,
            I => \N__27720\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27716\
        );

    \I__5447\ : CEMux
    port map (
            O => \N__27723\,
            I => \N__27713\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__27720\,
            I => \N__27710\
        );

    \I__5445\ : CEMux
    port map (
            O => \N__27719\,
            I => \N__27707\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__27716\,
            I => \N__27704\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27701\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__27710\,
            I => \N__27698\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27694\
        );

    \I__5440\ : Span4Mux_h
    port map (
            O => \N__27704\,
            I => \N__27691\
        );

    \I__5439\ : Span4Mux_h
    port map (
            O => \N__27701\,
            I => \N__27688\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__27698\,
            I => \N__27685\
        );

    \I__5437\ : CEMux
    port map (
            O => \N__27697\,
            I => \N__27682\
        );

    \I__5436\ : Span4Mux_h
    port map (
            O => \N__27694\,
            I => \N__27679\
        );

    \I__5435\ : Span4Mux_v
    port map (
            O => \N__27691\,
            I => \N__27674\
        );

    \I__5434\ : Span4Mux_h
    port map (
            O => \N__27688\,
            I => \N__27674\
        );

    \I__5433\ : IoSpan4Mux
    port map (
            O => \N__27685\,
            I => \N__27671\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__27682\,
            I => \N__27668\
        );

    \I__5431\ : Span4Mux_h
    port map (
            O => \N__27679\,
            I => \N__27665\
        );

    \I__5430\ : Span4Mux_v
    port map (
            O => \N__27674\,
            I => \N__27662\
        );

    \I__5429\ : IoSpan4Mux
    port map (
            O => \N__27671\,
            I => \N__27659\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__27668\,
            I => \N__27656\
        );

    \I__5427\ : Span4Mux_s2_h
    port map (
            O => \N__27665\,
            I => \N__27653\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__27662\,
            I => \N__27650\
        );

    \I__5425\ : IoSpan4Mux
    port map (
            O => \N__27659\,
            I => \N__27645\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__27656\,
            I => \N__27645\
        );

    \I__5423\ : Span4Mux_v
    port map (
            O => \N__27653\,
            I => \N__27642\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__27650\,
            I => \N__27639\
        );

    \I__5421\ : Span4Mux_s3_h
    port map (
            O => \N__27645\,
            I => \N__27636\
        );

    \I__5420\ : Span4Mux_v
    port map (
            O => \N__27642\,
            I => \N__27633\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__27639\,
            I => \N__27630\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__27636\,
            I => \N__27627\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__27633\,
            I => \CONTROL.operand1_cnvZ0Z_0\
        );

    \I__5416\ : Odrv4
    port map (
            O => \N__27630\,
            I => \CONTROL.operand1_cnvZ0Z_0\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__27627\,
            I => \CONTROL.operand1_cnvZ0Z_0\
        );

    \I__5414\ : CascadeMux
    port map (
            O => \N__27620\,
            I => \ALU.c_RNI72MICZ0Z_15_cascade_\
        );

    \I__5413\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27614\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__5411\ : Odrv4
    port map (
            O => \N__27611\,
            I => \ALU.d_RNI4HG101Z0Z_7\
        );

    \I__5410\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27604\
        );

    \I__5409\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27590\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27583\
        );

    \I__5407\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27580\
        );

    \I__5406\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27577\
        );

    \I__5405\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27570\
        );

    \I__5404\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27570\
        );

    \I__5403\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27570\
        );

    \I__5402\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27567\
        );

    \I__5401\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27559\
        );

    \I__5400\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27559\
        );

    \I__5399\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27559\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__27594\,
            I => \N__27555\
        );

    \I__5397\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27551\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__27590\,
            I => \N__27547\
        );

    \I__5395\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27544\
        );

    \I__5394\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27541\
        );

    \I__5393\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27536\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__27586\,
            I => \N__27531\
        );

    \I__5391\ : Span4Mux_s3_v
    port map (
            O => \N__27583\,
            I => \N__27526\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27526\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__27577\,
            I => \N__27521\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__27570\,
            I => \N__27521\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__27567\,
            I => \N__27518\
        );

    \I__5386\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27515\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27512\
        );

    \I__5384\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27508\
        );

    \I__5383\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27503\
        );

    \I__5382\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27503\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__27551\,
            I => \N__27500\
        );

    \I__5380\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27496\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__27547\,
            I => \N__27493\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27488\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__27541\,
            I => \N__27488\
        );

    \I__5376\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27485\
        );

    \I__5375\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27482\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__27536\,
            I => \N__27479\
        );

    \I__5373\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27472\
        );

    \I__5372\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27472\
        );

    \I__5371\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27472\
        );

    \I__5370\ : Span4Mux_v
    port map (
            O => \N__27526\,
            I => \N__27469\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__27521\,
            I => \N__27466\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__27518\,
            I => \N__27463\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__27515\,
            I => \N__27460\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__27512\,
            I => \N__27457\
        );

    \I__5365\ : InMux
    port map (
            O => \N__27511\,
            I => \N__27454\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__27508\,
            I => \N__27451\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__27503\,
            I => \N__27446\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__27500\,
            I => \N__27446\
        );

    \I__5361\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27443\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__27496\,
            I => \N__27436\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__27493\,
            I => \N__27436\
        );

    \I__5358\ : Span4Mux_v
    port map (
            O => \N__27488\,
            I => \N__27436\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__27485\,
            I => \N__27431\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__27482\,
            I => \N__27431\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__27479\,
            I => \N__27428\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__27472\,
            I => \N__27425\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__27469\,
            I => \N__27414\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__27466\,
            I => \N__27414\
        );

    \I__5351\ : Span4Mux_v
    port map (
            O => \N__27463\,
            I => \N__27414\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__27460\,
            I => \N__27414\
        );

    \I__5349\ : Span4Mux_h
    port map (
            O => \N__27457\,
            I => \N__27414\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27405\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__27451\,
            I => \N__27405\
        );

    \I__5346\ : Span4Mux_h
    port map (
            O => \N__27446\,
            I => \N__27405\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__27443\,
            I => \N__27405\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__27436\,
            I => \N__27400\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__27431\,
            I => \N__27400\
        );

    \I__5342\ : Span4Mux_v
    port map (
            O => \N__27428\,
            I => \N__27395\
        );

    \I__5341\ : Span4Mux_s3_h
    port map (
            O => \N__27425\,
            I => \N__27395\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__27414\,
            I => \ALU.aluOut_10\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__27405\,
            I => \ALU.aluOut_10\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__27400\,
            I => \ALU.aluOut_10\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__27395\,
            I => \ALU.aluOut_10\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__27386\,
            I => \ALU.N_475_cascade_\
        );

    \I__5335\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__27380\,
            I => \ALU.rshift_7\
        );

    \I__5333\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27374\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__27374\,
            I => \N__27371\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__5330\ : Odrv4
    port map (
            O => \N__27368\,
            I => \ALU.g_RNI0MJNZ0Z_1\
        );

    \I__5329\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__5327\ : Span4Mux_h
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__5326\ : Odrv4
    port map (
            O => \N__27356\,
            I => \ALU.dout_6_ns_1_3\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__5324\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27345\
        );

    \I__5323\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27342\
        );

    \I__5322\ : CascadeMux
    port map (
            O => \N__27348\,
            I => \N__27339\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27331\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27331\
        );

    \I__5319\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27326\
        );

    \I__5318\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27326\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__27337\,
            I => \N__27322\
        );

    \I__5316\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27318\
        );

    \I__5315\ : Span4Mux_v
    port map (
            O => \N__27331\,
            I => \N__27315\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27312\
        );

    \I__5313\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27309\
        );

    \I__5312\ : InMux
    port map (
            O => \N__27322\,
            I => \N__27304\
        );

    \I__5311\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27304\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__27318\,
            I => \N__27299\
        );

    \I__5309\ : Sp12to4
    port map (
            O => \N__27315\,
            I => \N__27299\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__27312\,
            I => \N__27296\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__27309\,
            I => \aluOperand1_2_rep1\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__27304\,
            I => \aluOperand1_2_rep1\
        );

    \I__5305\ : Odrv12
    port map (
            O => \N__27299\,
            I => \aluOperand1_2_rep1\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__27296\,
            I => \aluOperand1_2_rep1\
        );

    \I__5303\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27284\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__27284\,
            I => \N__27281\
        );

    \I__5301\ : Span4Mux_h
    port map (
            O => \N__27281\,
            I => \N__27278\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__27278\,
            I => \ALU.dout_6_ns_1_4\
        );

    \I__5299\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__27272\,
            I => \N__27269\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__27269\,
            I => \N__27266\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__27266\,
            I => \ALU.N_747\
        );

    \I__5295\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27260\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27257\
        );

    \I__5293\ : Span4Mux_v
    port map (
            O => \N__27257\,
            I => \N__27253\
        );

    \I__5292\ : InMux
    port map (
            O => \N__27256\,
            I => \N__27250\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__27253\,
            I => \ALU.N_699\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__27250\,
            I => \ALU.N_699\
        );

    \I__5289\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__27236\,
            I => \N__27232\
        );

    \I__5285\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__27232\,
            I => \N__27226\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27223\
        );

    \I__5282\ : Span4Mux_h
    port map (
            O => \N__27226\,
            I => \N__27220\
        );

    \I__5281\ : Span12Mux_s10_v
    port map (
            O => \N__27223\,
            I => \N__27217\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__27220\,
            I => \ALU.N_404_1\
        );

    \I__5279\ : Odrv12
    port map (
            O => \N__27217\,
            I => \ALU.N_404_1\
        );

    \I__5278\ : CascadeMux
    port map (
            O => \N__27212\,
            I => \N__27209\
        );

    \I__5277\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27206\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__27206\,
            I => \N__27203\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__27203\,
            I => \ALU.dout_6_ns_1_6\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__27200\,
            I => \ALU.N_753_cascade_\
        );

    \I__5273\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27192\
        );

    \I__5272\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27189\
        );

    \I__5271\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27186\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27182\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__27189\,
            I => \N__27177\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__27186\,
            I => \N__27177\
        );

    \I__5267\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27174\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__27182\,
            I => \N__27171\
        );

    \I__5265\ : Span4Mux_v
    port map (
            O => \N__27177\,
            I => \N__27168\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27165\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__27171\,
            I => \N__27162\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__27168\,
            I => \N__27159\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__27165\,
            I => \N__27156\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__27162\,
            I => \N__27148\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__27159\,
            I => \N__27148\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__27156\,
            I => \N__27148\
        );

    \I__5257\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27145\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__27148\,
            I => \N__27142\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__27145\,
            I => \N__27139\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__27142\,
            I => \testWordZ0Z_9\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__27139\,
            I => \testWordZ0Z_9\
        );

    \I__5252\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27121\
        );

    \I__5251\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27117\
        );

    \I__5250\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27114\
        );

    \I__5249\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27109\
        );

    \I__5248\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27109\
        );

    \I__5247\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27103\
        );

    \I__5246\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27103\
        );

    \I__5245\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27100\
        );

    \I__5244\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27097\
        );

    \I__5243\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27092\
        );

    \I__5242\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27092\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__27121\,
            I => \N__27089\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__27120\,
            I => \N__27086\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27083\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__27114\,
            I => \N__27078\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__27109\,
            I => \N__27078\
        );

    \I__5236\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27075\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__27103\,
            I => \N__27072\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27069\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__27097\,
            I => \N__27062\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__27092\,
            I => \N__27062\
        );

    \I__5231\ : Span4Mux_v
    port map (
            O => \N__27089\,
            I => \N__27062\
        );

    \I__5230\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27059\
        );

    \I__5229\ : Span4Mux_v
    port map (
            O => \N__27083\,
            I => \N__27054\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__27078\,
            I => \N__27054\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__27075\,
            I => \aluOperand1_fast_1\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__27072\,
            I => \aluOperand1_fast_1\
        );

    \I__5225\ : Odrv12
    port map (
            O => \N__27069\,
            I => \aluOperand1_fast_1\
        );

    \I__5224\ : Odrv4
    port map (
            O => \N__27062\,
            I => \aluOperand1_fast_1\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__27059\,
            I => \aluOperand1_fast_1\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__27054\,
            I => \aluOperand1_fast_1\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__27041\,
            I => \N__27036\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__27040\,
            I => \N__27033\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__27039\,
            I => \N__27030\
        );

    \I__5218\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27021\
        );

    \I__5217\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27021\
        );

    \I__5216\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27018\
        );

    \I__5215\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27015\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__27028\,
            I => \N__27012\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__27027\,
            I => \N__27008\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__27026\,
            I => \N__27005\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__27021\,
            I => \N__27002\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__26997\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__27015\,
            I => \N__26997\
        );

    \I__5208\ : InMux
    port map (
            O => \N__27012\,
            I => \N__26990\
        );

    \I__5207\ : InMux
    port map (
            O => \N__27011\,
            I => \N__26990\
        );

    \I__5206\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26990\
        );

    \I__5205\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26987\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__27002\,
            I => \N__26984\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__26997\,
            I => \aluOperand1_fast_2\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__26990\,
            I => \aluOperand1_fast_2\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__26987\,
            I => \aluOperand1_fast_2\
        );

    \I__5200\ : Odrv4
    port map (
            O => \N__26984\,
            I => \aluOperand1_fast_2\
        );

    \I__5199\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26972\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__26972\,
            I => \N__26969\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__26969\,
            I => \N__26966\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__26966\,
            I => \ALU.dout_3_ns_1_4\
        );

    \I__5195\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26960\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__26960\,
            I => \N__26956\
        );

    \I__5193\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26953\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__26956\,
            I => \N__26950\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__26953\,
            I => \ALU.eZ0Z_4\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__26950\,
            I => \ALU.eZ0Z_4\
        );

    \I__5189\ : InMux
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__26942\,
            I => \N__26939\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__26939\,
            I => \N__26936\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__26936\,
            I => \ALU.e_RNIS97JZ0Z_1\
        );

    \I__5185\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26929\
        );

    \I__5184\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26926\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__26929\,
            I => \N__26923\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__26926\,
            I => \ALU.eZ0Z_1\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__26923\,
            I => \ALU.eZ0Z_1\
        );

    \I__5180\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__26915\,
            I => \ALU.N_701\
        );

    \I__5178\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__26909\,
            I => \ALU.dout_3_ns_1_2\
        );

    \I__5176\ : InMux
    port map (
            O => \N__26906\,
            I => \N__26903\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__26903\,
            I => \N__26900\
        );

    \I__5174\ : Odrv12
    port map (
            O => \N__26900\,
            I => \ALU.dout_6_ns_1_7\
        );

    \I__5173\ : InMux
    port map (
            O => \N__26897\,
            I => \N__26894\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__26894\,
            I => \N__26891\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__26891\,
            I => \N__26888\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__26885\,
            I => \ALU.f_RNIQQJ01Z0Z_7\
        );

    \I__5168\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26874\
        );

    \I__5167\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26874\
        );

    \I__5166\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26869\
        );

    \I__5165\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26869\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__26874\,
            I => \N__26866\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26863\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__26866\,
            I => \N__26860\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__26863\,
            I => \N__26857\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__5159\ : Sp12to4
    port map (
            O => \N__26857\,
            I => \N__26851\
        );

    \I__5158\ : Span4Mux_v
    port map (
            O => \N__26854\,
            I => \N__26848\
        );

    \I__5157\ : Span12Mux_v
    port map (
            O => \N__26851\,
            I => \N__26845\
        );

    \I__5156\ : Span4Mux_v
    port map (
            O => \N__26848\,
            I => \N__26841\
        );

    \I__5155\ : Span12Mux_h
    port map (
            O => \N__26845\,
            I => \N__26838\
        );

    \I__5154\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26835\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__26841\,
            I => \testWordZ0Z_8\
        );

    \I__5152\ : Odrv12
    port map (
            O => \N__26838\,
            I => \testWordZ0Z_8\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__26835\,
            I => \testWordZ0Z_8\
        );

    \I__5150\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26823\
        );

    \I__5149\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26820\
        );

    \I__5148\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26817\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__26823\,
            I => \N__26812\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26812\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__26817\,
            I => \N__26809\
        );

    \I__5144\ : Span4Mux_v
    port map (
            O => \N__26812\,
            I => \N__26806\
        );

    \I__5143\ : Odrv12
    port map (
            O => \N__26809\,
            I => \ALU.fZ0Z_10\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__26806\,
            I => \ALU.fZ0Z_10\
        );

    \I__5141\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__26798\,
            I => \N__26795\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__26795\,
            I => \N__26792\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__26792\,
            I => \N__26789\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__26789\,
            I => \ALU.b_RNIEHSD1Z0Z_10\
        );

    \I__5136\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26780\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__5133\ : Span4Mux_h
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__26774\,
            I => \ALU.madd_cry_13_ma\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__26771\,
            I => \N__26768\
        );

    \I__5130\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__5128\ : Span4Mux_h
    port map (
            O => \N__26762\,
            I => \N__26759\
        );

    \I__5127\ : Span4Mux_h
    port map (
            O => \N__26759\,
            I => \N__26756\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__26756\,
            I => \ALU.madd_axb_13_l_ofx\
        );

    \I__5125\ : InMux
    port map (
            O => \N__26753\,
            I => \ALU.madd_cry_12\
        );

    \I__5124\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26747\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__26747\,
            I => \N__26744\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__26744\,
            I => \N__26741\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__26738\,
            I => \ALU.madd_axb_14\
        );

    \I__5119\ : InMux
    port map (
            O => \N__26735\,
            I => \ALU.madd_cry_13\
        );

    \I__5118\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26722\
        );

    \I__5117\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26722\
        );

    \I__5116\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26717\
        );

    \I__5115\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26717\
        );

    \I__5114\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26712\
        );

    \I__5113\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26708\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__26722\,
            I => \N__26705\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26702\
        );

    \I__5110\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26697\
        );

    \I__5109\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26697\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__26712\,
            I => \N__26694\
        );

    \I__5107\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26691\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__26708\,
            I => \N__26686\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__26705\,
            I => \N__26683\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__26702\,
            I => \N__26678\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__26697\,
            I => \N__26678\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__26694\,
            I => \N__26673\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26673\
        );

    \I__5100\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26668\
        );

    \I__5099\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26668\
        );

    \I__5098\ : Span12Mux_s6_h
    port map (
            O => \N__26686\,
            I => \N__26665\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__26683\,
            I => \N__26660\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__26678\,
            I => \N__26660\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__26673\,
            I => \ALU.operand2_6\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__26668\,
            I => \ALU.operand2_6\
        );

    \I__5093\ : Odrv12
    port map (
            O => \N__26665\,
            I => \ALU.operand2_6\
        );

    \I__5092\ : Odrv4
    port map (
            O => \N__26660\,
            I => \ALU.operand2_6\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__26651\,
            I => \N__26646\
        );

    \I__5090\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26643\
        );

    \I__5089\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26638\
        );

    \I__5088\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26634\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26631\
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__26642\,
            I => \N__26628\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__26641\,
            I => \N__26623\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__26638\,
            I => \N__26620\
        );

    \I__5083\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26617\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__26634\,
            I => \N__26612\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__26631\,
            I => \N__26612\
        );

    \I__5080\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26609\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__26627\,
            I => \N__26606\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__26626\,
            I => \N__26592\
        );

    \I__5077\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26589\
        );

    \I__5076\ : Span4Mux_s1_v
    port map (
            O => \N__26620\,
            I => \N__26583\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26583\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__26612\,
            I => \N__26578\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__26609\,
            I => \N__26578\
        );

    \I__5072\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26572\
        );

    \I__5071\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26569\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__26604\,
            I => \N__26565\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__26603\,
            I => \N__26561\
        );

    \I__5068\ : CascadeMux
    port map (
            O => \N__26602\,
            I => \N__26558\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__26601\,
            I => \N__26555\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__26600\,
            I => \N__26550\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__26599\,
            I => \N__26546\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__26598\,
            I => \N__26543\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__26597\,
            I => \N__26540\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__26596\,
            I => \N__26537\
        );

    \I__5061\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26530\
        );

    \I__5060\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26530\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__26589\,
            I => \N__26527\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__26588\,
            I => \N__26524\
        );

    \I__5057\ : Span4Mux_v
    port map (
            O => \N__26583\,
            I => \N__26518\
        );

    \I__5056\ : Span4Mux_v
    port map (
            O => \N__26578\,
            I => \N__26518\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__26577\,
            I => \N__26515\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__26576\,
            I => \N__26511\
        );

    \I__5053\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26508\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__26572\,
            I => \N__26503\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__26569\,
            I => \N__26503\
        );

    \I__5050\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26500\
        );

    \I__5049\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26487\
        );

    \I__5048\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26487\
        );

    \I__5047\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26487\
        );

    \I__5046\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26484\
        );

    \I__5045\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26477\
        );

    \I__5044\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26477\
        );

    \I__5043\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26477\
        );

    \I__5042\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26468\
        );

    \I__5041\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26468\
        );

    \I__5040\ : InMux
    port map (
            O => \N__26546\,
            I => \N__26468\
        );

    \I__5039\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26468\
        );

    \I__5038\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26463\
        );

    \I__5037\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26463\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \N__26460\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__26535\,
            I => \N__26457\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__26530\,
            I => \N__26452\
        );

    \I__5033\ : Span4Mux_v
    port map (
            O => \N__26527\,
            I => \N__26452\
        );

    \I__5032\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26449\
        );

    \I__5031\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26446\
        );

    \I__5030\ : Span4Mux_h
    port map (
            O => \N__26518\,
            I => \N__26442\
        );

    \I__5029\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26439\
        );

    \I__5028\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26436\
        );

    \I__5027\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26433\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__26508\,
            I => \N__26428\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__26503\,
            I => \N__26428\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__26500\,
            I => \N__26425\
        );

    \I__5023\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26418\
        );

    \I__5022\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26418\
        );

    \I__5021\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26418\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__26496\,
            I => \N__26415\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__26495\,
            I => \N__26412\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__26494\,
            I => \N__26409\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__26487\,
            I => \N__26404\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__26484\,
            I => \N__26404\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26401\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26398\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26395\
        );

    \I__5012\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26390\
        );

    \I__5011\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26390\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__26452\,
            I => \N__26387\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26384\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__26446\,
            I => \N__26381\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__26445\,
            I => \N__26376\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__26442\,
            I => \N__26370\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__26439\,
            I => \N__26370\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__26436\,
            I => \N__26363\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__26433\,
            I => \N__26363\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__26428\,
            I => \N__26363\
        );

    \I__5001\ : Span4Mux_s1_h
    port map (
            O => \N__26425\,
            I => \N__26358\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__26418\,
            I => \N__26358\
        );

    \I__4999\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26355\
        );

    \I__4998\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26352\
        );

    \I__4997\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26349\
        );

    \I__4996\ : Sp12to4
    port map (
            O => \N__26404\,
            I => \N__26346\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__26401\,
            I => \N__26341\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__26398\,
            I => \N__26341\
        );

    \I__4993\ : Span4Mux_h
    port map (
            O => \N__26395\,
            I => \N__26334\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26334\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__26387\,
            I => \N__26334\
        );

    \I__4990\ : Span4Mux_v
    port map (
            O => \N__26384\,
            I => \N__26329\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__26381\,
            I => \N__26329\
        );

    \I__4988\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26320\
        );

    \I__4987\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26320\
        );

    \I__4986\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26320\
        );

    \I__4985\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26320\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__26370\,
            I => \N__26317\
        );

    \I__4983\ : Span4Mux_v
    port map (
            O => \N__26363\,
            I => \N__26314\
        );

    \I__4982\ : Sp12to4
    port map (
            O => \N__26358\,
            I => \N__26303\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__26355\,
            I => \N__26303\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__26352\,
            I => \N__26303\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__26349\,
            I => \N__26303\
        );

    \I__4978\ : Span12Mux_h
    port map (
            O => \N__26346\,
            I => \N__26303\
        );

    \I__4977\ : Span4Mux_h
    port map (
            O => \N__26341\,
            I => \N__26298\
        );

    \I__4976\ : Span4Mux_v
    port map (
            O => \N__26334\,
            I => \N__26298\
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__26329\,
            I => \aluReadBus\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__26320\,
            I => \aluReadBus\
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__26317\,
            I => \aluReadBus\
        );

    \I__4972\ : Odrv4
    port map (
            O => \N__26314\,
            I => \aluReadBus\
        );

    \I__4971\ : Odrv12
    port map (
            O => \N__26303\,
            I => \aluReadBus\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__26298\,
            I => \aluReadBus\
        );

    \I__4969\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26271\
        );

    \I__4968\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26271\
        );

    \I__4967\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26268\
        );

    \I__4966\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26265\
        );

    \I__4965\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26262\
        );

    \I__4964\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26259\
        );

    \I__4963\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26254\
        );

    \I__4962\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26254\
        );

    \I__4961\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26248\
        );

    \I__4960\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26248\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__26271\,
            I => \N__26245\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__26268\,
            I => \N__26242\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__26265\,
            I => \N__26237\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26237\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__26259\,
            I => \N__26232\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26232\
        );

    \I__4953\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26229\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__26248\,
            I => \N__26226\
        );

    \I__4951\ : Span4Mux_h
    port map (
            O => \N__26245\,
            I => \N__26223\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__26242\,
            I => \N__26220\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__26237\,
            I => \N__26215\
        );

    \I__4948\ : Span4Mux_h
    port map (
            O => \N__26232\,
            I => \N__26215\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__26229\,
            I => \N__26212\
        );

    \I__4946\ : Span4Mux_h
    port map (
            O => \N__26226\,
            I => \N__26209\
        );

    \I__4945\ : Span4Mux_s0_h
    port map (
            O => \N__26223\,
            I => \N__26206\
        );

    \I__4944\ : Span4Mux_v
    port map (
            O => \N__26220\,
            I => \N__26201\
        );

    \I__4943\ : Span4Mux_h
    port map (
            O => \N__26215\,
            I => \N__26201\
        );

    \I__4942\ : Odrv12
    port map (
            O => \N__26212\,
            I => \ALU.N_217_0\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__26209\,
            I => \ALU.N_217_0\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__26206\,
            I => \ALU.N_217_0\
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__26201\,
            I => \ALU.N_217_0\
        );

    \I__4938\ : CascadeMux
    port map (
            O => \N__26192\,
            I => \ALU.dout_3_ns_1_15_cascade_\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__26189\,
            I => \ALU.dout_6_ns_1_2_cascade_\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__26186\,
            I => \ALU.N_749_cascade_\
        );

    \I__4935\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26176\
        );

    \I__4933\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26173\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__26176\,
            I => \N__26170\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__26173\,
            I => \N__26167\
        );

    \I__4930\ : Sp12to4
    port map (
            O => \N__26170\,
            I => \N__26162\
        );

    \I__4929\ : Span12Mux_h
    port map (
            O => \N__26167\,
            I => \N__26162\
        );

    \I__4928\ : Odrv12
    port map (
            O => \N__26162\,
            I => \ALU.madd_52\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__4926\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26153\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__26153\,
            I => \N__26150\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__26150\,
            I => \N__26147\
        );

    \I__4923\ : Span4Mux_h
    port map (
            O => \N__26147\,
            I => \N__26144\
        );

    \I__4922\ : Span4Mux_v
    port map (
            O => \N__26144\,
            I => \N__26141\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__26141\,
            I => \ALU.madd_axb_5_l_fx\
        );

    \I__4920\ : InMux
    port map (
            O => \N__26138\,
            I => \ALU.madd_cry_4\
        );

    \I__4919\ : InMux
    port map (
            O => \N__26135\,
            I => \ALU.madd_cry_5\
        );

    \I__4918\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26129\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__26129\,
            I => \N__26125\
        );

    \I__4916\ : InMux
    port map (
            O => \N__26128\,
            I => \N__26122\
        );

    \I__4915\ : Span4Mux_v
    port map (
            O => \N__26125\,
            I => \N__26117\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__26122\,
            I => \N__26117\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__26117\,
            I => \N__26114\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__26114\,
            I => \N__26111\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__26111\,
            I => \ALU.madd_axb_7\
        );

    \I__4910\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__26102\,
            I => \ALU.madd_cry_6_THRU_CO\
        );

    \I__4907\ : InMux
    port map (
            O => \N__26099\,
            I => \ALU.madd_cry_6\
        );

    \I__4906\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__4903\ : Span4Mux_h
    port map (
            O => \N__26087\,
            I => \N__26084\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__26081\,
            I => \ALU.madd_axb_8_l_fx\
        );

    \I__4900\ : CascadeMux
    port map (
            O => \N__26078\,
            I => \N__26075\
        );

    \I__4899\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__26072\,
            I => \N__26069\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__26069\,
            I => \N__26065\
        );

    \I__4896\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26062\
        );

    \I__4895\ : Span4Mux_h
    port map (
            O => \N__26065\,
            I => \N__26059\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__26062\,
            I => \ALU.madd_159\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__26059\,
            I => \ALU.madd_159\
        );

    \I__4892\ : InMux
    port map (
            O => \N__26054\,
            I => \bfn_9_10_0_\
        );

    \I__4891\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__26048\,
            I => \N__26045\
        );

    \I__4889\ : Span12Mux_h
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__4888\ : Odrv12
    port map (
            O => \N__26042\,
            I => \ALU.madd_cry_9_ma\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__4886\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26033\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__4884\ : Span4Mux_h
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__4883\ : Span4Mux_v
    port map (
            O => \N__26027\,
            I => \N__26024\
        );

    \I__4882\ : Span4Mux_h
    port map (
            O => \N__26024\,
            I => \N__26021\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__26021\,
            I => \ALU.madd_axb_9_l_ofx\
        );

    \I__4880\ : InMux
    port map (
            O => \N__26018\,
            I => \ALU.madd_cry_8\
        );

    \I__4879\ : InMux
    port map (
            O => \N__26015\,
            I => \N__26012\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__4876\ : Span4Mux_h
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__4875\ : Span4Mux_h
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__26000\,
            I => \ALU.madd_cry_10_ma\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__4872\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__4870\ : Span12Mux_h
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__4869\ : Odrv12
    port map (
            O => \N__25985\,
            I => \ALU.madd_axb_10_l_ofx\
        );

    \I__4868\ : InMux
    port map (
            O => \N__25982\,
            I => \ALU.madd_cry_9\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__4866\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25973\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__25973\,
            I => \N__25970\
        );

    \I__4864\ : Span12Mux_h
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__4863\ : Odrv12
    port map (
            O => \N__25967\,
            I => \ALU.madd_axb_11\
        );

    \I__4862\ : InMux
    port map (
            O => \N__25964\,
            I => \ALU.madd_cry_10\
        );

    \I__4861\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__25958\,
            I => \N__25955\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__25955\,
            I => \N__25952\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__4857\ : Span4Mux_s1_h
    port map (
            O => \N__25949\,
            I => \N__25946\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__25946\,
            I => \ALU.madd_axb_12_l_fx\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__4854\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25937\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__25937\,
            I => \N__25934\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__25934\,
            I => \N__25930\
        );

    \I__4851\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25927\
        );

    \I__4850\ : Span4Mux_h
    port map (
            O => \N__25930\,
            I => \N__25924\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__25927\,
            I => \ALU.madd_360\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__25924\,
            I => \ALU.madd_360\
        );

    \I__4847\ : InMux
    port map (
            O => \N__25919\,
            I => \ALU.madd_cry_11\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__4845\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25909\
        );

    \I__4844\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25906\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__25909\,
            I => \N__25901\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__25906\,
            I => \N__25901\
        );

    \I__4841\ : Span4Mux_v
    port map (
            O => \N__25901\,
            I => \N__25898\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__25895\,
            I => \ALU.fZ0Z_15\
        );

    \I__4838\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25889\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__4835\ : Span4Mux_v
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__25880\,
            I => \ALU.madd_cry_0_ma\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__4832\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25871\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__25871\,
            I => \N__25868\
        );

    \I__4830\ : Span4Mux_h
    port map (
            O => \N__25868\,
            I => \N__25865\
        );

    \I__4829\ : Span4Mux_h
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__4828\ : Span4Mux_v
    port map (
            O => \N__25862\,
            I => \N__25859\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__25859\,
            I => \ALU.madd_cry_1_ma\
        );

    \I__4826\ : InMux
    port map (
            O => \N__25856\,
            I => \ALU.madd_cry_0\
        );

    \I__4825\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25850\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__25850\,
            I => \N__25847\
        );

    \I__4823\ : Span4Mux_h
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__4822\ : Span4Mux_v
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__25841\,
            I => \ALU.madd_axb_2_l_fx\
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__4819\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__25832\,
            I => \N__25828\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__25831\,
            I => \N__25825\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__25828\,
            I => \N__25822\
        );

    \I__4815\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25819\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__25822\,
            I => \N__25816\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__25819\,
            I => \N__25813\
        );

    \I__4812\ : Span4Mux_v
    port map (
            O => \N__25816\,
            I => \N__25810\
        );

    \I__4811\ : Span4Mux_v
    port map (
            O => \N__25813\,
            I => \N__25807\
        );

    \I__4810\ : Sp12to4
    port map (
            O => \N__25810\,
            I => \N__25804\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__25807\,
            I => \N__25801\
        );

    \I__4808\ : Odrv12
    port map (
            O => \N__25804\,
            I => \ALU.madd_6\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__25801\,
            I => \ALU.madd_6\
        );

    \I__4806\ : InMux
    port map (
            O => \N__25796\,
            I => \ALU.madd_cry_1\
        );

    \I__4805\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25790\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__4803\ : Span4Mux_h
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__25784\,
            I => \ALU.madd_13\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__4800\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__25772\,
            I => \N__25769\
        );

    \I__4797\ : Span4Mux_v
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__25763\,
            I => \ALU.madd_18\
        );

    \I__4794\ : InMux
    port map (
            O => \N__25760\,
            I => \ALU.madd_cry_2\
        );

    \I__4793\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__4791\ : Span4Mux_h
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__25745\,
            I => \ALU.madd_axb_4_l_fx\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__25742\,
            I => \N__25738\
        );

    \I__4787\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25735\
        );

    \I__4786\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25732\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__25735\,
            I => \N__25729\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25726\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__25729\,
            I => \N__25721\
        );

    \I__4782\ : Span4Mux_v
    port map (
            O => \N__25726\,
            I => \N__25721\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__25718\,
            I => \ALU.madd_30\
        );

    \I__4779\ : InMux
    port map (
            O => \N__25715\,
            I => \ALU.madd_cry_3\
        );

    \I__4778\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25709\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25706\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__25706\,
            I => \N__25703\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__25700\,
            I => \ALU.d_RNICJE9BZ0Z_8\
        );

    \I__4773\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__25688\,
            I => \ALU.d_RNIEUKR11Z0Z_0\
        );

    \I__4769\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25682\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__4767\ : Span4Mux_v
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__4766\ : Span4Mux_h
    port map (
            O => \N__25676\,
            I => \N__25673\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__25673\,
            I => \N__25670\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__25670\,
            I => \ALU.a_15_m3_8\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__25667\,
            I => \ALU.a_15_m4_8_cascade_\
        );

    \I__4762\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25661\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__25661\,
            I => \ALU.a_15_m5_8\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__25658\,
            I => \N__25655\
        );

    \I__4759\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25651\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__25654\,
            I => \N__25648\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__25651\,
            I => \N__25645\
        );

    \I__4756\ : InMux
    port map (
            O => \N__25648\,
            I => \N__25642\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__25645\,
            I => \N__25639\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__25642\,
            I => \N__25636\
        );

    \I__4753\ : Span4Mux_h
    port map (
            O => \N__25639\,
            I => \N__25631\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__25636\,
            I => \N__25631\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__25631\,
            I => \ALU.fZ0Z_8\
        );

    \I__4750\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25624\
        );

    \I__4749\ : InMux
    port map (
            O => \N__25627\,
            I => \N__25621\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__25624\,
            I => \N__25618\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25615\
        );

    \I__4746\ : Span12Mux_v
    port map (
            O => \N__25618\,
            I => \N__25612\
        );

    \I__4745\ : Odrv12
    port map (
            O => \N__25615\,
            I => \ALU.dZ0Z_8\
        );

    \I__4744\ : Odrv12
    port map (
            O => \N__25612\,
            I => \ALU.dZ0Z_8\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__25607\,
            I => \ALU.operand2_6_ns_1_8_cascade_\
        );

    \I__4742\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25601\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__25601\,
            I => \N__25598\
        );

    \I__4740\ : Odrv12
    port map (
            O => \N__25598\,
            I => \ALU.N_867\
        );

    \I__4739\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25592\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__25589\,
            I => \N__25586\
        );

    \I__4736\ : Span4Mux_h
    port map (
            O => \N__25586\,
            I => \N__25582\
        );

    \I__4735\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25579\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__25582\,
            I => \ALU.hZ0Z_8\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__25579\,
            I => \ALU.hZ0Z_8\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__25574\,
            I => \ALU.N_186_0_i_cascade_\
        );

    \I__4731\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__25559\,
            I => \ALU.c_RNIA7OEEZ0Z_11\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__4725\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__25547\,
            I => \N__25542\
        );

    \I__4722\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25539\
        );

    \I__4721\ : CascadeMux
    port map (
            O => \N__25545\,
            I => \N__25535\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__25542\,
            I => \N__25531\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__25539\,
            I => \N__25528\
        );

    \I__4718\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25525\
        );

    \I__4717\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25522\
        );

    \I__4716\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25519\
        );

    \I__4715\ : Span4Mux_h
    port map (
            O => \N__25531\,
            I => \N__25516\
        );

    \I__4714\ : Span4Mux_s1_v
    port map (
            O => \N__25528\,
            I => \N__25513\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__25525\,
            I => \N__25506\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__25522\,
            I => \N__25506\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__25519\,
            I => \N__25506\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__25516\,
            I => \RXbuffer_5\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__25513\,
            I => \RXbuffer_5\
        );

    \I__4708\ : Odrv12
    port map (
            O => \N__25506\,
            I => \RXbuffer_5\
        );

    \I__4707\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25496\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__25496\,
            I => \N__25493\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__25493\,
            I => \N__25489\
        );

    \I__4704\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25486\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__25489\,
            I => \ALU.hZ0Z_12\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__25486\,
            I => \ALU.hZ0Z_12\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__25481\,
            I => \ALU.c_RNIJ949Z0Z_12_cascade_\
        );

    \I__4700\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25475\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__25475\,
            I => \ALU.a_RNIFPBOZ0Z_12\
        );

    \I__4698\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25469\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__25469\,
            I => \ALU.d_RNIM5LUZ0Z_12\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__25466\,
            I => \ALU.operand2_7_ns_1_12_cascade_\
        );

    \I__4695\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25454\
        );

    \I__4694\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25454\
        );

    \I__4693\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25454\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__25454\,
            I => \N__25449\
        );

    \I__4691\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25446\
        );

    \I__4690\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25443\
        );

    \I__4689\ : Span4Mux_h
    port map (
            O => \N__25449\,
            I => \N__25439\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__25446\,
            I => \N__25434\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25434\
        );

    \I__4686\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25431\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__25439\,
            I => \N__25428\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__25434\,
            I => \N__25423\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25423\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__25428\,
            I => \ALU.operand2_12\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__25423\,
            I => \ALU.operand2_12\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__25418\,
            I => \ALU.N_636_cascade_\
        );

    \I__4679\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__4677\ : Span4Mux_h
    port map (
            O => \N__25409\,
            I => \N__25406\
        );

    \I__4676\ : Span4Mux_h
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__4674\ : Span4Mux_v
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__25397\,
            I => \ALU.N_272_0\
        );

    \I__4672\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__4670\ : Span4Mux_h
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__25382\,
            I => \ALU.N_264_0\
        );

    \I__4667\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25374\
        );

    \I__4666\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25367\
        );

    \I__4665\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25364\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N__25361\
        );

    \I__4663\ : InMux
    port map (
            O => \N__25373\,
            I => \N__25356\
        );

    \I__4662\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25356\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__25371\,
            I => \N__25349\
        );

    \I__4660\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25345\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__25367\,
            I => \N__25335\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__25364\,
            I => \N__25335\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__25361\,
            I => \N__25330\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__25356\,
            I => \N__25330\
        );

    \I__4655\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25327\
        );

    \I__4654\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25323\
        );

    \I__4653\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25316\
        );

    \I__4652\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25316\
        );

    \I__4651\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25316\
        );

    \I__4650\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25313\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__25345\,
            I => \N__25310\
        );

    \I__4648\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25301\
        );

    \I__4647\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25301\
        );

    \I__4646\ : InMux
    port map (
            O => \N__25342\,
            I => \N__25301\
        );

    \I__4645\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25301\
        );

    \I__4644\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25298\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__25335\,
            I => \N__25295\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__25330\,
            I => \N__25290\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__25327\,
            I => \N__25290\
        );

    \I__4640\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25285\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__25323\,
            I => \N__25282\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__25316\,
            I => \N__25279\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__25313\,
            I => \N__25274\
        );

    \I__4636\ : Span4Mux_v
    port map (
            O => \N__25310\,
            I => \N__25274\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25269\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__25298\,
            I => \N__25269\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__25295\,
            I => \N__25264\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__25290\,
            I => \N__25264\
        );

    \I__4631\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25259\
        );

    \I__4630\ : InMux
    port map (
            O => \N__25288\,
            I => \N__25259\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__25285\,
            I => \N__25252\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__25282\,
            I => \N__25252\
        );

    \I__4627\ : Span4Mux_s3_h
    port map (
            O => \N__25279\,
            I => \N__25252\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__25274\,
            I => \ALU.aluOut_12\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__25269\,
            I => \ALU.aluOut_12\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__25264\,
            I => \ALU.aluOut_12\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__25259\,
            I => \ALU.aluOut_12\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__25252\,
            I => \ALU.aluOut_12\
        );

    \I__4621\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25238\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__25238\,
            I => \ALU.N_462\
        );

    \I__4619\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__25232\,
            I => \ALU.N_270_0\
        );

    \I__4617\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__25226\,
            I => \N__25222\
        );

    \I__4615\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25217\
        );

    \I__4614\ : Span4Mux_v
    port map (
            O => \N__25222\,
            I => \N__25210\
        );

    \I__4613\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25207\
        );

    \I__4612\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25201\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__25217\,
            I => \N__25198\
        );

    \I__4610\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25195\
        );

    \I__4609\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25192\
        );

    \I__4608\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25189\
        );

    \I__4607\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25186\
        );

    \I__4606\ : Span4Mux_s1_h
    port map (
            O => \N__25210\,
            I => \N__25183\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25180\
        );

    \I__4604\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25177\
        );

    \I__4603\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25174\
        );

    \I__4602\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25171\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25166\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__25198\,
            I => \N__25159\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__25195\,
            I => \N__25159\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__25192\,
            I => \N__25156\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__25189\,
            I => \N__25151\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__25186\,
            I => \N__25151\
        );

    \I__4595\ : Sp12to4
    port map (
            O => \N__25183\,
            I => \N__25148\
        );

    \I__4594\ : Span4Mux_h
    port map (
            O => \N__25180\,
            I => \N__25145\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25140\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__25174\,
            I => \N__25140\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__25171\,
            I => \N__25136\
        );

    \I__4590\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25133\
        );

    \I__4589\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25130\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__25166\,
            I => \N__25127\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__25165\,
            I => \N__25124\
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__25164\,
            I => \N__25119\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__25159\,
            I => \N__25111\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__25156\,
            I => \N__25111\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__25151\,
            I => \N__25111\
        );

    \I__4582\ : Span12Mux_s4_h
    port map (
            O => \N__25148\,
            I => \N__25108\
        );

    \I__4581\ : Span4Mux_v
    port map (
            O => \N__25145\,
            I => \N__25103\
        );

    \I__4580\ : Span4Mux_h
    port map (
            O => \N__25140\,
            I => \N__25103\
        );

    \I__4579\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25100\
        );

    \I__4578\ : Span12Mux_h
    port map (
            O => \N__25136\,
            I => \N__25091\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25091\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__25130\,
            I => \N__25091\
        );

    \I__4575\ : Sp12to4
    port map (
            O => \N__25127\,
            I => \N__25091\
        );

    \I__4574\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25084\
        );

    \I__4573\ : InMux
    port map (
            O => \N__25123\,
            I => \N__25084\
        );

    \I__4572\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25084\
        );

    \I__4571\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25079\
        );

    \I__4570\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25079\
        );

    \I__4569\ : Span4Mux_v
    port map (
            O => \N__25111\,
            I => \N__25076\
        );

    \I__4568\ : Odrv12
    port map (
            O => \N__25108\,
            I => \aluReadBus_fast\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__25103\,
            I => \aluReadBus_fast\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__25100\,
            I => \aluReadBus_fast\
        );

    \I__4565\ : Odrv12
    port map (
            O => \N__25091\,
            I => \aluReadBus_fast\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__25084\,
            I => \aluReadBus_fast\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__25079\,
            I => \aluReadBus_fast\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__25076\,
            I => \aluReadBus_fast\
        );

    \I__4561\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25057\
        );

    \I__4560\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25054\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__25057\,
            I => \N__25049\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__25054\,
            I => \N__25046\
        );

    \I__4557\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25043\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__25052\,
            I => \N__25040\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__25049\,
            I => \N__25036\
        );

    \I__4554\ : Span4Mux_h
    port map (
            O => \N__25046\,
            I => \N__25031\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__25043\,
            I => \N__25031\
        );

    \I__4552\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25026\
        );

    \I__4551\ : InMux
    port map (
            O => \N__25039\,
            I => \N__25026\
        );

    \I__4550\ : Span4Mux_v
    port map (
            O => \N__25036\,
            I => \N__25023\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__25031\,
            I => \N__25020\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__25026\,
            I => \ALU.N_175_0\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__25023\,
            I => \ALU.N_175_0\
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__25020\,
            I => \ALU.N_175_0\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__25013\,
            I => \ALU.N_175_0_cascade_\
        );

    \I__4544\ : InMux
    port map (
            O => \N__25010\,
            I => \N__25003\
        );

    \I__4543\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__4542\ : InMux
    port map (
            O => \N__25008\,
            I => \N__25000\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__24996\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__25000\,
            I => \N__24993\
        );

    \I__4539\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24990\
        );

    \I__4538\ : Span4Mux_h
    port map (
            O => \N__24996\,
            I => \N__24985\
        );

    \I__4537\ : Span4Mux_h
    port map (
            O => \N__24993\,
            I => \N__24985\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__24990\,
            I => \ALU.operand2_13\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__24985\,
            I => \ALU.operand2_13\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__24980\,
            I => \ALU.un2_addsub_axb_13_cascade_\
        );

    \I__4533\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24974\,
            I => \N__24970\
        );

    \I__4531\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24966\
        );

    \I__4530\ : Span4Mux_v
    port map (
            O => \N__24970\,
            I => \N__24963\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24960\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__24966\,
            I => \N__24957\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__24963\,
            I => \N__24954\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__24960\,
            I => \ALU.N_177_0\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__24957\,
            I => \ALU.N_177_0\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__24954\,
            I => \ALU.N_177_0\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__24947\,
            I => \N__24944\
        );

    \I__4522\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24941\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__24941\,
            I => \N__24938\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__24938\,
            I => \N__24935\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__24935\,
            I => \N__24932\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__24932\,
            I => \N__24929\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__24929\,
            I => \ALU.d_RNI9FOTEZ0Z_13\
        );

    \I__4516\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24923\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__24923\,
            I => \N__24919\
        );

    \I__4514\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24916\
        );

    \I__4513\ : Span4Mux_v
    port map (
            O => \N__24919\,
            I => \N__24913\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__24916\,
            I => \N__24910\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__24913\,
            I => \N__24906\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__24910\,
            I => \N__24902\
        );

    \I__4509\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24899\
        );

    \I__4508\ : Span4Mux_h
    port map (
            O => \N__24906\,
            I => \N__24896\
        );

    \I__4507\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24893\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__24902\,
            I => \N__24889\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__24899\,
            I => \N__24886\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__24896\,
            I => \N__24883\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__24893\,
            I => \N__24880\
        );

    \I__4502\ : CascadeMux
    port map (
            O => \N__24892\,
            I => \N__24877\
        );

    \I__4501\ : Span4Mux_v
    port map (
            O => \N__24889\,
            I => \N__24872\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__24886\,
            I => \N__24872\
        );

    \I__4499\ : Span4Mux_s1_h
    port map (
            O => \N__24883\,
            I => \N__24867\
        );

    \I__4498\ : Span4Mux_h
    port map (
            O => \N__24880\,
            I => \N__24867\
        );

    \I__4497\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24864\
        );

    \I__4496\ : Span4Mux_v
    port map (
            O => \N__24872\,
            I => \N__24861\
        );

    \I__4495\ : Span4Mux_h
    port map (
            O => \N__24867\,
            I => \N__24858\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24853\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__24861\,
            I => \N__24853\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__24858\,
            I => \ctrlOut_11\
        );

    \I__4491\ : Odrv4
    port map (
            O => \N__24853\,
            I => \ctrlOut_11\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__4489\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__4487\ : Span12Mux_s8_h
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__4486\ : Odrv12
    port map (
            O => \N__24836\,
            I => \ALU.N_186_0_i\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__24833\,
            I => \ALU.a_15_m4_bm_1Z0Z_2_cascade_\
        );

    \I__4484\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__24827\,
            I => \N__24824\
        );

    \I__4482\ : Odrv4
    port map (
            O => \N__24824\,
            I => \ALU.d_RNIII58AZ0Z_2\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__24821\,
            I => \ALU.rshift_3_ns_1_2_cascade_\
        );

    \I__4480\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__24812\,
            I => \ALU.N_470\
        );

    \I__4477\ : InMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__24800\,
            I => \ALU.N_376\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__24797\,
            I => \ALU.N_589_cascade_\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__24794\,
            I => \ALU.rshift_1_13_cascade_\
        );

    \I__4471\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__4469\ : Span4Mux_h
    port map (
            O => \N__24785\,
            I => \N__24782\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__24782\,
            I => \ALU.a_15_m3_13\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__24779\,
            I => \ALU.N_576_cascade_\
        );

    \I__4466\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24769\
        );

    \I__4464\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24763\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__24769\,
            I => \N__24760\
        );

    \I__4462\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24753\
        );

    \I__4461\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24753\
        );

    \I__4460\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24753\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__24763\,
            I => \FTDI.RXstateZ0Z_2\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__24760\,
            I => \FTDI.RXstateZ0Z_2\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__24753\,
            I => \FTDI.RXstateZ0Z_2\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__24746\,
            I => \FTDI.N_23_cascade_\
        );

    \I__4455\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24733\
        );

    \I__4454\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24733\
        );

    \I__4453\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24733\
        );

    \I__4452\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24730\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__24733\,
            I => \N__24727\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__24730\,
            I => \N__24724\
        );

    \I__4449\ : Span4Mux_s1_v
    port map (
            O => \N__24727\,
            I => \N__24719\
        );

    \I__4448\ : Span4Mux_s1_v
    port map (
            O => \N__24724\,
            I => \N__24716\
        );

    \I__4447\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24711\
        );

    \I__4446\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24711\
        );

    \I__4445\ : Span4Mux_h
    port map (
            O => \N__24719\,
            I => \N__24708\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__24716\,
            I => \FTDI.RXstateZ0Z_1\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__24711\,
            I => \FTDI.RXstateZ0Z_1\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__24708\,
            I => \FTDI.RXstateZ0Z_1\
        );

    \I__4441\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__24692\,
            I => \FTDI.m13_ns_1\
        );

    \I__4437\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24683\
        );

    \I__4436\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24683\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__24683\,
            I => \N__24677\
        );

    \I__4434\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24670\
        );

    \I__4433\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24670\
        );

    \I__4432\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24670\
        );

    \I__4431\ : Span4Mux_s1_v
    port map (
            O => \N__24677\,
            I => \N__24667\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__24670\,
            I => \FTDI.RXstateZ0Z_0\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__24667\,
            I => \FTDI.RXstateZ0Z_0\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__24662\,
            I => \N__24656\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__24661\,
            I => \N__24653\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__24660\,
            I => \N__24649\
        );

    \I__4425\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24646\
        );

    \I__4424\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24636\
        );

    \I__4423\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24636\
        );

    \I__4422\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24636\
        );

    \I__4421\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24636\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24633\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__24645\,
            I => \N__24628\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__24636\,
            I => \N__24624\
        );

    \I__4417\ : Span4Mux_s1_v
    port map (
            O => \N__24633\,
            I => \N__24621\
        );

    \I__4416\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24612\
        );

    \I__4415\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24612\
        );

    \I__4414\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24612\
        );

    \I__4413\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24612\
        );

    \I__4412\ : Span4Mux_s1_v
    port map (
            O => \N__24624\,
            I => \N__24609\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__24621\,
            I => \FTDI.RXstateZ0Z_3\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__24612\,
            I => \FTDI.RXstateZ0Z_3\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__24609\,
            I => \FTDI.RXstateZ0Z_3\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__24602\,
            I => \ALU.a_15_sm0_cascade_\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__24599\,
            I => \ALU.a_15_m2_ns_1Z0Z_12_cascade_\
        );

    \I__4406\ : InMux
    port map (
            O => \N__24596\,
            I => \N__24589\
        );

    \I__4405\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24589\
        );

    \I__4404\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24584\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__24589\,
            I => \N__24581\
        );

    \I__4402\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24574\
        );

    \I__4401\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24574\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24571\
        );

    \I__4399\ : Span4Mux_s2_v
    port map (
            O => \N__24581\,
            I => \N__24568\
        );

    \I__4398\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24563\
        );

    \I__4397\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24563\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24558\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__24571\,
            I => \N__24558\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__24568\,
            I => \N__24555\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__24563\,
            I => \N__24552\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__24558\,
            I => \ALU.log_2_sqmuxa\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__24555\,
            I => \ALU.log_2_sqmuxa\
        );

    \I__4390\ : Odrv12
    port map (
            O => \N__24552\,
            I => \ALU.log_2_sqmuxa\
        );

    \I__4389\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24542\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__24536\,
            I => \ALU.a7_b_0\
        );

    \I__4385\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__24527\,
            I => \N__24523\
        );

    \I__4382\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24520\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__24523\,
            I => \ALU.a5_b_2\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__24520\,
            I => \ALU.a5_b_2\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__4378\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24506\
        );

    \I__4377\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24506\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24503\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__24503\,
            I => \ALU.madd_63\
        );

    \I__4374\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24497\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24494\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__24494\,
            I => \N__24491\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__24491\,
            I => \ALU.a2_b_1\
        );

    \I__4370\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24485\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__4368\ : Span4Mux_h
    port map (
            O => \N__24482\,
            I => \N__24478\
        );

    \I__4367\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24475\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__24478\,
            I => \ALU.a3_b_0\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__24475\,
            I => \ALU.a3_b_0\
        );

    \I__4364\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__4361\ : Span4Mux_h
    port map (
            O => \N__24461\,
            I => \N__24457\
        );

    \I__4360\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24454\
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__24457\,
            I => \ALU.a1_b_2\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__24454\,
            I => \ALU.a1_b_2\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__4356\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24443\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24440\
        );

    \I__4354\ : Span4Mux_v
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__24437\,
            I => \N__24434\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__24434\,
            I => \ALU.d_RNI2B0LZ0Z_9\
        );

    \I__4351\ : InMux
    port map (
            O => \N__24431\,
            I => \N__24428\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__24428\,
            I => \N__24424\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__24427\,
            I => \N__24420\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__24424\,
            I => \N__24417\
        );

    \I__4347\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24414\
        );

    \I__4346\ : InMux
    port map (
            O => \N__24420\,
            I => \N__24411\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__24417\,
            I => \ALU.hZ0Z_10\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__24414\,
            I => \ALU.hZ0Z_10\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__24411\,
            I => \ALU.hZ0Z_10\
        );

    \I__4342\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__4339\ : Span4Mux_v
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__24392\,
            I => \ALU.d_RNII1LUZ0Z_10\
        );

    \I__4337\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__24380\,
            I => \ALU.d_RNIO00LZ0Z_4\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__24377\,
            I => \N__24372\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__24376\,
            I => \N__24369\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__24375\,
            I => \N__24366\
        );

    \I__4330\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24361\
        );

    \I__4329\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24361\
        );

    \I__4328\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24358\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__24361\,
            I => \N__24355\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24352\
        );

    \I__4325\ : Span4Mux_v
    port map (
            O => \N__24355\,
            I => \N__24349\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__24352\,
            I => \N__24346\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__24349\,
            I => \ALU.a3_b_3\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__24346\,
            I => \ALU.a3_b_3\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__24341\,
            I => \N__24337\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__24340\,
            I => \N__24334\
        );

    \I__4319\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24329\
        );

    \I__4318\ : InMux
    port map (
            O => \N__24334\,
            I => \N__24329\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24326\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__24326\,
            I => \N__24322\
        );

    \I__4315\ : InMux
    port map (
            O => \N__24325\,
            I => \N__24319\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__24322\,
            I => \N__24308\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__24319\,
            I => \N__24305\
        );

    \I__4312\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24302\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__24317\,
            I => \N__24299\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__24316\,
            I => \N__24294\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__24315\,
            I => \N__24291\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \N__24287\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__24313\,
            I => \N__24284\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__24312\,
            I => \N__24280\
        );

    \I__4305\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24277\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__24308\,
            I => \N__24270\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__24305\,
            I => \N__24270\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24270\
        );

    \I__4301\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24267\
        );

    \I__4300\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24264\
        );

    \I__4299\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24260\
        );

    \I__4298\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24257\
        );

    \I__4297\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24254\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__24290\,
            I => \N__24250\
        );

    \I__4295\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24246\
        );

    \I__4294\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24243\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__24283\,
            I => \N__24239\
        );

    \I__4292\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24236\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__24277\,
            I => \N__24226\
        );

    \I__4290\ : Span4Mux_v
    port map (
            O => \N__24270\,
            I => \N__24226\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24223\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__24264\,
            I => \N__24220\
        );

    \I__4287\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24217\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__24260\,
            I => \N__24214\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__24257\,
            I => \N__24209\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24209\
        );

    \I__4283\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24202\
        );

    \I__4282\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24202\
        );

    \I__4281\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24202\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__24246\,
            I => \N__24197\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__24243\,
            I => \N__24197\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__24242\,
            I => \N__24194\
        );

    \I__4277\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24190\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24187\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \N__24184\
        );

    \I__4274\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24181\
        );

    \I__4273\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24176\
        );

    \I__4272\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24176\
        );

    \I__4271\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24173\
        );

    \I__4270\ : IoSpan4Mux
    port map (
            O => \N__24226\,
            I => \N__24170\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__24223\,
            I => \N__24161\
        );

    \I__4268\ : Span4Mux_s3_h
    port map (
            O => \N__24220\,
            I => \N__24161\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__24217\,
            I => \N__24161\
        );

    \I__4266\ : Span4Mux_s3_h
    port map (
            O => \N__24214\,
            I => \N__24161\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__24209\,
            I => \N__24154\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24154\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__24197\,
            I => \N__24154\
        );

    \I__4262\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24150\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__24193\,
            I => \N__24145\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24141\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__24187\,
            I => \N__24138\
        );

    \I__4258\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24135\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__24181\,
            I => \N__24131\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24128\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__24173\,
            I => \N__24121\
        );

    \I__4254\ : Span4Mux_s3_h
    port map (
            O => \N__24170\,
            I => \N__24121\
        );

    \I__4253\ : Span4Mux_v
    port map (
            O => \N__24161\,
            I => \N__24121\
        );

    \I__4252\ : Span4Mux_v
    port map (
            O => \N__24154\,
            I => \N__24118\
        );

    \I__4251\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24115\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__24150\,
            I => \N__24112\
        );

    \I__4249\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24107\
        );

    \I__4248\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24107\
        );

    \I__4247\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24104\
        );

    \I__4246\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24101\
        );

    \I__4245\ : Span12Mux_s4_h
    port map (
            O => \N__24141\,
            I => \N__24094\
        );

    \I__4244\ : Sp12to4
    port map (
            O => \N__24138\,
            I => \N__24094\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__24135\,
            I => \N__24094\
        );

    \I__4242\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24091\
        );

    \I__4241\ : Span4Mux_v
    port map (
            O => \N__24131\,
            I => \N__24082\
        );

    \I__4240\ : Span4Mux_s3_h
    port map (
            O => \N__24128\,
            I => \N__24082\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__24121\,
            I => \N__24082\
        );

    \I__4238\ : Span4Mux_h
    port map (
            O => \N__24118\,
            I => \N__24082\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__24115\,
            I => \aluReadBus_rep1\
        );

    \I__4236\ : Odrv12
    port map (
            O => \N__24112\,
            I => \aluReadBus_rep1\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__24107\,
            I => \aluReadBus_rep1\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__24104\,
            I => \aluReadBus_rep1\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__24101\,
            I => \aluReadBus_rep1\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__24094\,
            I => \aluReadBus_rep1\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__24091\,
            I => \aluReadBus_rep1\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__24082\,
            I => \aluReadBus_rep1\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__24065\,
            I => \N__24061\
        );

    \I__4228\ : InMux
    port map (
            O => \N__24064\,
            I => \N__24056\
        );

    \I__4227\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24056\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__4225\ : Span4Mux_h
    port map (
            O => \N__24053\,
            I => \N__24050\
        );

    \I__4224\ : Span4Mux_h
    port map (
            O => \N__24050\,
            I => \N__24047\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__24047\,
            I => \ALU.a2_b_3\
        );

    \I__4222\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24039\
        );

    \I__4221\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24034\
        );

    \I__4220\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24034\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__24039\,
            I => \N__24031\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__24034\,
            I => \N__24026\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__24031\,
            I => \N__24023\
        );

    \I__4216\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24019\
        );

    \I__4215\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24016\
        );

    \I__4214\ : Span4Mux_v
    port map (
            O => \N__24026\,
            I => \N__24010\
        );

    \I__4213\ : Span4Mux_v
    port map (
            O => \N__24023\,
            I => \N__24007\
        );

    \I__4212\ : InMux
    port map (
            O => \N__24022\,
            I => \N__24004\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__24019\,
            I => \N__24001\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__24016\,
            I => \N__23998\
        );

    \I__4209\ : InMux
    port map (
            O => \N__24015\,
            I => \N__23991\
        );

    \I__4208\ : InMux
    port map (
            O => \N__24014\,
            I => \N__23991\
        );

    \I__4207\ : InMux
    port map (
            O => \N__24013\,
            I => \N__23991\
        );

    \I__4206\ : Span4Mux_v
    port map (
            O => \N__24010\,
            I => \N__23988\
        );

    \I__4205\ : Sp12to4
    port map (
            O => \N__24007\,
            I => \N__23983\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__24004\,
            I => \N__23983\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__24001\,
            I => \N__23980\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__23998\,
            I => \N__23975\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23975\
        );

    \I__4200\ : Sp12to4
    port map (
            O => \N__23988\,
            I => \N__23969\
        );

    \I__4199\ : Span12Mux_s6_h
    port map (
            O => \N__23983\,
            I => \N__23964\
        );

    \I__4198\ : Sp12to4
    port map (
            O => \N__23980\,
            I => \N__23964\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__23975\,
            I => \N__23961\
        );

    \I__4196\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23954\
        );

    \I__4195\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23954\
        );

    \I__4194\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23954\
        );

    \I__4193\ : Odrv12
    port map (
            O => \N__23969\,
            I => \ALU.operand2_3\
        );

    \I__4192\ : Odrv12
    port map (
            O => \N__23964\,
            I => \ALU.operand2_3\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__23961\,
            I => \ALU.operand2_3\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__23954\,
            I => \ALU.operand2_3\
        );

    \I__4189\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23941\
        );

    \I__4188\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23934\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__23941\,
            I => \N__23931\
        );

    \I__4186\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23922\
        );

    \I__4185\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23922\
        );

    \I__4184\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23922\
        );

    \I__4183\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23922\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__23934\,
            I => \N__23913\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__23931\,
            I => \N__23910\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23907\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__23921\,
            I => \N__23904\
        );

    \I__4178\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23901\
        );

    \I__4177\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23894\
        );

    \I__4176\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23894\
        );

    \I__4175\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23894\
        );

    \I__4174\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23891\
        );

    \I__4173\ : Span4Mux_v
    port map (
            O => \N__23913\,
            I => \N__23888\
        );

    \I__4172\ : Span4Mux_s3_h
    port map (
            O => \N__23910\,
            I => \N__23885\
        );

    \I__4171\ : Span4Mux_v
    port map (
            O => \N__23907\,
            I => \N__23882\
        );

    \I__4170\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23879\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__23901\,
            I => \N__23876\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23873\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23868\
        );

    \I__4166\ : Span4Mux_v
    port map (
            O => \N__23888\,
            I => \N__23868\
        );

    \I__4165\ : Span4Mux_v
    port map (
            O => \N__23885\,
            I => \N__23863\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__23882\,
            I => \N__23863\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__23879\,
            I => \ALU.N_235_0\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__23876\,
            I => \ALU.N_235_0\
        );

    \I__4161\ : Odrv12
    port map (
            O => \N__23873\,
            I => \ALU.N_235_0\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__23868\,
            I => \ALU.N_235_0\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__23863\,
            I => \ALU.N_235_0\
        );

    \I__4158\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__23849\,
            I => \ALU.un2_addsub_axb_3\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__4155\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23840\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__23840\,
            I => \N__23837\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__4152\ : Span4Mux_v
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__23831\,
            I => \ALU.d_RNIDK21BZ0Z_3\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__23828\,
            I => \ALU.dout_3_ns_1_3_cascade_\
        );

    \I__4149\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23822\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__23822\,
            I => \ALU.N_702\
        );

    \I__4147\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23816\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__23816\,
            I => \ALU.g_RNII4LLZ0Z_3\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \ALU.e_RNITOVJZ0Z_3_cascade_\
        );

    \I__4144\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__23807\,
            I => \ALU.operand2_7_ns_1_3\
        );

    \I__4142\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__4140\ : Span12Mux_v
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__23795\,
            I => \ALU.un2_addsub_cry_6_c_RNIL4LMIZ0\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__23792\,
            I => \ALU.operand2_3_ns_1_6_cascade_\
        );

    \I__4137\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23786\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__23786\,
            I => \ALU.N_817\
        );

    \I__4135\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23776\
        );

    \I__4133\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23772\
        );

    \I__4132\ : Span4Mux_s2_h
    port map (
            O => \N__23776\,
            I => \N__23769\
        );

    \I__4131\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23766\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23761\
        );

    \I__4129\ : Span4Mux_v
    port map (
            O => \N__23769\,
            I => \N__23761\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__23766\,
            I => \N__23758\
        );

    \I__4127\ : Span4Mux_h
    port map (
            O => \N__23761\,
            I => \N__23755\
        );

    \I__4126\ : Odrv12
    port map (
            O => \N__23758\,
            I => \ALU.a6_b_6\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__23755\,
            I => \ALU.a6_b_6\
        );

    \I__4124\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23746\
        );

    \I__4123\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23743\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__23746\,
            I => \N__23740\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__23743\,
            I => \N__23737\
        );

    \I__4120\ : Span4Mux_s3_h
    port map (
            O => \N__23740\,
            I => \N__23734\
        );

    \I__4119\ : Span4Mux_s3_h
    port map (
            O => \N__23737\,
            I => \N__23731\
        );

    \I__4118\ : Span4Mux_v
    port map (
            O => \N__23734\,
            I => \N__23728\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__23731\,
            I => \N__23723\
        );

    \I__4116\ : Span4Mux_h
    port map (
            O => \N__23728\,
            I => \N__23723\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__23723\,
            I => \ALU.a3_b_6\
        );

    \I__4114\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__23717\,
            I => \ALU.operand2_6_ns_1_6\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__23714\,
            I => \ALU.N_750_cascade_\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__23711\,
            I => \ALU.operand2_3_cascade_\
        );

    \I__4110\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23703\
        );

    \I__4109\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23700\
        );

    \I__4108\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23697\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__23703\,
            I => \N__23694\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23691\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__23697\,
            I => \N__23688\
        );

    \I__4104\ : Span4Mux_h
    port map (
            O => \N__23694\,
            I => \N__23685\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__23691\,
            I => \ALU.aZ0Z_10\
        );

    \I__4102\ : Odrv12
    port map (
            O => \N__23688\,
            I => \ALU.aZ0Z_10\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__23685\,
            I => \ALU.aZ0Z_10\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__23678\,
            I => \ALU.dout_3_ns_1_10_cascade_\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__23675\,
            I => \ALU.dout_6_ns_1_10_cascade_\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__23672\,
            I => \ALU.N_757_cascade_\
        );

    \I__4097\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__23666\,
            I => \ALU.N_709\
        );

    \I__4095\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__4093\ : Span4Mux_h
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__23654\,
            I => \ALU.dout_6_ns_1_5\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__23651\,
            I => \ALU.N_865_cascade_\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__23648\,
            I => \ALU.d_RNI61SHAZ0Z_1_cascade_\
        );

    \I__4089\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__23642\,
            I => \ALU.d_RNIJM067Z0Z_1\
        );

    \I__4087\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__4085\ : Span12Mux_s4_v
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__4084\ : Odrv12
    port map (
            O => \N__23630\,
            I => \ALU.a_15_m2_1\
        );

    \I__4083\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \ALU.g_RNIK6LLZ0Z_4_cascade_\
        );

    \I__4082\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__23621\,
            I => \ALU.e_RNIGQ8HZ0Z_4\
        );

    \I__4080\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23612\
        );

    \I__4079\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23612\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__4077\ : Odrv12
    port map (
            O => \N__23609\,
            I => \ALU.a1_b_4\
        );

    \I__4076\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23602\
        );

    \I__4075\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23599\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__23602\,
            I => \N__23596\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__23599\,
            I => \N__23593\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__23596\,
            I => \N__23590\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__23593\,
            I => \N__23587\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__23590\,
            I => \N__23584\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__23587\,
            I => \ALU.a2_b_4\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__23584\,
            I => \ALU.a2_b_4\
        );

    \I__4067\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__23576\,
            I => \ALU.operand2_7_ns_1_4\
        );

    \I__4065\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23563\
        );

    \I__4063\ : InMux
    port map (
            O => \N__23569\,
            I => \N__23560\
        );

    \I__4062\ : InMux
    port map (
            O => \N__23568\,
            I => \N__23555\
        );

    \I__4061\ : InMux
    port map (
            O => \N__23567\,
            I => \N__23552\
        );

    \I__4060\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23549\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__23563\,
            I => \N__23544\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__23560\,
            I => \N__23544\
        );

    \I__4057\ : InMux
    port map (
            O => \N__23559\,
            I => \N__23539\
        );

    \I__4056\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23539\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__23555\,
            I => \N__23534\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__23552\,
            I => \N__23534\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23531\
        );

    \I__4052\ : Span4Mux_v
    port map (
            O => \N__23544\,
            I => \N__23528\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__23539\,
            I => \N__23525\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__23534\,
            I => \N__23520\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__23531\,
            I => \N__23513\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__23528\,
            I => \N__23513\
        );

    \I__4047\ : Span4Mux_v
    port map (
            O => \N__23525\,
            I => \N__23513\
        );

    \I__4046\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23508\
        );

    \I__4045\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23508\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__23520\,
            I => \ALU.operand2_4\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__23513\,
            I => \ALU.operand2_4\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__23508\,
            I => \ALU.operand2_4\
        );

    \I__4041\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23497\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__23500\,
            I => \N__23494\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__23497\,
            I => \N__23490\
        );

    \I__4038\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23480\
        );

    \I__4037\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23480\
        );

    \I__4036\ : Span4Mux_s2_h
    port map (
            O => \N__23490\,
            I => \N__23477\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__23489\,
            I => \N__23474\
        );

    \I__4034\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23469\
        );

    \I__4033\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23469\
        );

    \I__4032\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23465\
        );

    \I__4031\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23462\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__23480\,
            I => \N__23457\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__23477\,
            I => \N__23457\
        );

    \I__4028\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23453\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23450\
        );

    \I__4026\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23447\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23443\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__23462\,
            I => \N__23440\
        );

    \I__4023\ : Sp12to4
    port map (
            O => \N__23457\,
            I => \N__23437\
        );

    \I__4022\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23434\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23429\
        );

    \I__4020\ : Span4Mux_h
    port map (
            O => \N__23450\,
            I => \N__23429\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__23447\,
            I => \N__23426\
        );

    \I__4018\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23423\
        );

    \I__4017\ : Span12Mux_s3_h
    port map (
            O => \N__23443\,
            I => \N__23420\
        );

    \I__4016\ : Span4Mux_v
    port map (
            O => \N__23440\,
            I => \N__23417\
        );

    \I__4015\ : Span12Mux_v
    port map (
            O => \N__23437\,
            I => \N__23414\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N__23409\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__23429\,
            I => \N__23409\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__23426\,
            I => \ALU.N_229_0\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__23423\,
            I => \ALU.N_229_0\
        );

    \I__4010\ : Odrv12
    port map (
            O => \N__23420\,
            I => \ALU.N_229_0\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__23417\,
            I => \ALU.N_229_0\
        );

    \I__4008\ : Odrv12
    port map (
            O => \N__23414\,
            I => \ALU.N_229_0\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__23409\,
            I => \ALU.N_229_0\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \ALU.operand2_4_cascade_\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__23393\,
            I => \ALU.N_231_0_cascade_\
        );

    \I__4004\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__23381\,
            I => \ALU.madd_93_0\
        );

    \I__4000\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__23375\,
            I => \ALU.N_758\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__23372\,
            I => \ALU.N_710_cascade_\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__23369\,
            I => \ALU.aluOut_11_cascade_\
        );

    \I__3996\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__3994\ : Span4Mux_h
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__23357\,
            I => \ALU.madd_484_6\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__23354\,
            I => \ALU.un2_addsub_axb_1_cascade_\
        );

    \I__3991\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__23348\,
            I => \ALU.d_RNIC4AT9Z0Z_1\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \ALU.dout_7_ns_1_1_cascade_\
        );

    \I__3988\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23333\
        );

    \I__3986\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23330\
        );

    \I__3985\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23327\
        );

    \I__3984\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23324\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__23333\,
            I => \N__23321\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23316\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23316\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__23324\,
            I => \N__23313\
        );

    \I__3979\ : Sp12to4
    port map (
            O => \N__23321\,
            I => \N__23308\
        );

    \I__3978\ : Span12Mux_h
    port map (
            O => \N__23316\,
            I => \N__23308\
        );

    \I__3977\ : Sp12to4
    port map (
            O => \N__23313\,
            I => \N__23305\
        );

    \I__3976\ : Odrv12
    port map (
            O => \N__23308\,
            I => \ALU.N_247_0\
        );

    \I__3975\ : Odrv12
    port map (
            O => \N__23305\,
            I => \ALU.N_247_0\
        );

    \I__3974\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23294\
        );

    \I__3973\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23294\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3971\ : Span4Mux_h
    port map (
            O => \N__23291\,
            I => \N__23287\
        );

    \I__3970\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23284\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__23287\,
            I => \ALU.operand2_1\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__23284\,
            I => \ALU.operand2_1\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__23279\,
            I => \N__23275\
        );

    \I__3966\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23272\
        );

    \I__3965\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__23269\,
            I => \ALU.N_249_0\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__23266\,
            I => \ALU.N_249_0\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__23261\,
            I => \ALU.N_249_0_cascade_\
        );

    \I__3960\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__23255\,
            I => \ALU.a_15_m2_10\
        );

    \I__3958\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23249\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__23249\,
            I => \ALU.a_15_m2_ns_1Z0Z_10\
        );

    \I__3956\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__23240\,
            I => \ALU.un2_addsub_cry_9_c_RNIVCOFAZ0\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__23237\,
            I => \un9_addsub_cry_9_c_RNI8H83V_cascade_\
        );

    \I__3952\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__23231\,
            I => \c_RNI5V90O2_10\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \aluOperation_RNINNN4N3_0_cascade_\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__23225\,
            I => \ALU.dout_6_ns_1_11_cascade_\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__23222\,
            I => \ALU.dout_3_ns_1_11_cascade_\
        );

    \I__3947\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__23210\,
            I => \N__23206\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__23209\,
            I => \N__23203\
        );

    \I__3942\ : Sp12to4
    port map (
            O => \N__23206\,
            I => \N__23200\
        );

    \I__3941\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23197\
        );

    \I__3940\ : Odrv12
    port map (
            O => \N__23200\,
            I => \ALU.a0_b_4\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__23197\,
            I => \ALU.a0_b_4\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__23192\,
            I => \ALU.a1_b_3_cascade_\
        );

    \I__3937\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23185\
        );

    \I__3936\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23182\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23179\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__3933\ : Span4Mux_h
    port map (
            O => \N__23179\,
            I => \N__23173\
        );

    \I__3932\ : Span4Mux_v
    port map (
            O => \N__23176\,
            I => \N__23170\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__23173\,
            I => \ALU.madd_0\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__23170\,
            I => \ALU.madd_0\
        );

    \I__3929\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__23159\,
            I => \N__23155\
        );

    \I__3926\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23152\
        );

    \I__3925\ : Span4Mux_h
    port map (
            O => \N__23155\,
            I => \N__23149\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__23152\,
            I => \ALU.a0_b_3\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__23149\,
            I => \ALU.a0_b_3\
        );

    \I__3922\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23138\
        );

    \I__3921\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23134\
        );

    \I__3920\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23129\
        );

    \I__3919\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23129\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__23138\,
            I => \N__23126\
        );

    \I__3917\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23123\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__23134\,
            I => \N__23118\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__23129\,
            I => \N__23118\
        );

    \I__3914\ : Odrv12
    port map (
            O => \N__23126\,
            I => \ALU.N_375\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__23123\,
            I => \ALU.N_375\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__23118\,
            I => \ALU.N_375\
        );

    \I__3911\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23108\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__23108\,
            I => \ALU.rshift_3_ns_1_0\
        );

    \I__3909\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23101\
        );

    \I__3908\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23098\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23093\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23093\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__23093\,
            I => \ALU.N_249\
        );

    \I__3904\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23086\
        );

    \I__3903\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23083\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__23086\,
            I => \ALU.N_245\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__23083\,
            I => \ALU.N_245\
        );

    \I__3900\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__23072\,
            I => \ALU.lshift_10\
        );

    \I__3897\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__23060\,
            I => \ALU.a_15_m3_10\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__23057\,
            I => \ALU.a_15_m4_10_cascade_\
        );

    \I__3892\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23049\
        );

    \I__3891\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23044\
        );

    \I__3890\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23044\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__23040\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23037\
        );

    \I__3887\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23034\
        );

    \I__3886\ : Odrv12
    port map (
            O => \N__23040\,
            I => \ALU.N_377\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__23037\,
            I => \ALU.N_377\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__23034\,
            I => \ALU.N_377\
        );

    \I__3883\ : CascadeMux
    port map (
            O => \N__23027\,
            I => \ALU.N_377_cascade_\
        );

    \I__3882\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23021\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__23021\,
            I => \ALU.N_216\
        );

    \I__3880\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__23015\,
            I => \ALU.N_404\
        );

    \I__3878\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23005\
        );

    \I__3876\ : InMux
    port map (
            O => \N__23008\,
            I => \N__23002\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__23005\,
            I => \ALU.N_246\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__23002\,
            I => \ALU.N_246\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__22997\,
            I => \ALU.N_376_cascade_\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \ALU.d_RNIEBMRAZ0Z_0_cascade_\
        );

    \I__3871\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22988\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__22988\,
            I => \ALU.d_RNI1GH4VZ0Z_7\
        );

    \I__3869\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22982\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__22979\,
            I => \N__22976\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__22973\,
            I => \ALU.N_468\
        );

    \I__3864\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__22967\,
            I => \N__22964\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__22958\,
            I => \ALU.a1_b_3\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__22955\,
            I => \ALU.d_RNIA28GU1Z0Z_1_cascade_\
        );

    \I__3858\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__22949\,
            I => \ALU.d_RNIJ1PCQZ0Z_1\
        );

    \I__3856\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22943\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__3854\ : Span4Mux_v
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__22937\,
            I => \ALU.N_225\
        );

    \I__3852\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22930\
        );

    \I__3851\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22927\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22924\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__22927\,
            I => \ALU.N_223\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__22924\,
            I => \ALU.N_223\
        );

    \I__3847\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22912\
        );

    \I__3845\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22909\
        );

    \I__3844\ : Span4Mux_h
    port map (
            O => \N__22912\,
            I => \N__22906\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22903\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__22906\,
            I => \ALU.N_221\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__22903\,
            I => \ALU.N_221\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__22898\,
            I => \ALU.lshift_7_ns_1_13_cascade_\
        );

    \I__3839\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22888\
        );

    \I__3838\ : InMux
    port map (
            O => \N__22894\,
            I => \N__22888\
        );

    \I__3837\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22885\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22882\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__3834\ : Span4Mux_h
    port map (
            O => \N__22882\,
            I => \N__22876\
        );

    \I__3833\ : Odrv12
    port map (
            O => \N__22879\,
            I => \ALU.N_219\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__22876\,
            I => \ALU.N_219\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__22871\,
            I => \ALU.N_315_cascade_\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__22868\,
            I => \ALU.lshift_13_cascade_\
        );

    \I__3829\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22862\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__22859\,
            I => \ALU.a_15_m2_13\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__22856\,
            I => \ALU.a_15_m4_13_cascade_\
        );

    \I__3825\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__22850\,
            I => \ALU.N_247\
        );

    \I__3823\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22844\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__22844\,
            I => \ALU.lshift_15_ns_1_15\
        );

    \I__3821\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22835\
        );

    \I__3820\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22835\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__22835\,
            I => \ALU.N_416\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__22832\,
            I => \ALU.rshift_3_ns_1_9_cascade_\
        );

    \I__3817\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__22826\,
            I => \ALU.rshift_3_ns_1_1\
        );

    \I__3815\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22817\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__22817\,
            I => \ALU.d_RNINEO9E_0Z0Z_1\
        );

    \I__3812\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__22811\,
            I => \N__22807\
        );

    \I__3810\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22804\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__22807\,
            I => \N__22800\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__22804\,
            I => \N__22797\
        );

    \I__3807\ : InMux
    port map (
            O => \N__22803\,
            I => \N__22794\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__22800\,
            I => \ALU.N_217\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__22797\,
            I => \ALU.N_217\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__22794\,
            I => \ALU.N_217\
        );

    \I__3803\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__22784\,
            I => \ALU.lshift_7_ns_1_9\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__22781\,
            I => \ALU.N_311_cascade_\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__22778\,
            I => \ALU.lshift_9_cascade_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__3797\ : Span4Mux_h
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__22766\,
            I => \ALU.a_15_m2_9\
        );

    \I__3795\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__3793\ : Span4Mux_h
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__22754\,
            I => \ALU.N_292_0\
        );

    \I__3791\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__22748\,
            I => \ALU.rshift_1\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__22745\,
            I => \ALU.N_473_cascade_\
        );

    \I__3788\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__22739\,
            I => \ALU.m42_nsZ0Z_1\
        );

    \I__3786\ : CascadeMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__3785\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22726\
        );

    \I__3783\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22716\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__22726\,
            I => \N__22712\
        );

    \I__3781\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22707\
        );

    \I__3780\ : InMux
    port map (
            O => \N__22724\,
            I => \N__22707\
        );

    \I__3779\ : InMux
    port map (
            O => \N__22723\,
            I => \N__22700\
        );

    \I__3778\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22700\
        );

    \I__3777\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22700\
        );

    \I__3776\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22693\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__22719\,
            I => \N__22688\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22681\
        );

    \I__3773\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22678\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__22712\,
            I => \N__22669\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__22707\,
            I => \N__22669\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__22700\,
            I => \N__22666\
        );

    \I__3769\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22657\
        );

    \I__3768\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22657\
        );

    \I__3767\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22657\
        );

    \I__3766\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22657\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__22693\,
            I => \N__22654\
        );

    \I__3764\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22645\
        );

    \I__3763\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22645\
        );

    \I__3762\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22645\
        );

    \I__3761\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22645\
        );

    \I__3760\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22638\
        );

    \I__3759\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22638\
        );

    \I__3758\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22638\
        );

    \I__3757\ : Span4Mux_s1_v
    port map (
            O => \N__22681\,
            I => \N__22635\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22632\
        );

    \I__3755\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22623\
        );

    \I__3754\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22623\
        );

    \I__3753\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22623\
        );

    \I__3752\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22623\
        );

    \I__3751\ : Span4Mux_s1_v
    port map (
            O => \N__22669\,
            I => \N__22618\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__22666\,
            I => \N__22618\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__22657\,
            I => \testWordZ0Z_1\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__22654\,
            I => \testWordZ0Z_1\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__22645\,
            I => \testWordZ0Z_1\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__22638\,
            I => \testWordZ0Z_1\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__22635\,
            I => \testWordZ0Z_1\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__22632\,
            I => \testWordZ0Z_1\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__22623\,
            I => \testWordZ0Z_1\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__22618\,
            I => \testWordZ0Z_1\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__22601\,
            I => \N__22591\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__22600\,
            I => \N__22588\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__22599\,
            I => \N__22585\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__22598\,
            I => \N__22578\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__22597\,
            I => \N__22575\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__22596\,
            I => \N__22570\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__22595\,
            I => \N__22566\
        );

    \I__3734\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22559\
        );

    \I__3733\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22559\
        );

    \I__3732\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22559\
        );

    \I__3731\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22556\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__22584\,
            I => \N__22552\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__22583\,
            I => \N__22549\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__22582\,
            I => \N__22546\
        );

    \I__3727\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22537\
        );

    \I__3726\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22537\
        );

    \I__3725\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22537\
        );

    \I__3724\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22537\
        );

    \I__3723\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22530\
        );

    \I__3722\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22530\
        );

    \I__3721\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22530\
        );

    \I__3720\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22527\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22520\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22520\
        );

    \I__3717\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22511\
        );

    \I__3716\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22511\
        );

    \I__3715\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22511\
        );

    \I__3714\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22511\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__22537\,
            I => \N__22508\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__22530\,
            I => \N__22505\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__22527\,
            I => \N__22501\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__22526\,
            I => \N__22498\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__22525\,
            I => \N__22494\
        );

    \I__3708\ : Span4Mux_s3_v
    port map (
            O => \N__22520\,
            I => \N__22489\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22482\
        );

    \I__3706\ : Span4Mux_h
    port map (
            O => \N__22508\,
            I => \N__22482\
        );

    \I__3705\ : Span4Mux_s1_v
    port map (
            O => \N__22505\,
            I => \N__22482\
        );

    \I__3704\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22479\
        );

    \I__3703\ : Span4Mux_h
    port map (
            O => \N__22501\,
            I => \N__22476\
        );

    \I__3702\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22473\
        );

    \I__3701\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22468\
        );

    \I__3700\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22468\
        );

    \I__3699\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22463\
        );

    \I__3698\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22463\
        );

    \I__3697\ : Span4Mux_h
    port map (
            O => \N__22489\,
            I => \N__22460\
        );

    \I__3696\ : Span4Mux_h
    port map (
            O => \N__22482\,
            I => \N__22457\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__22479\,
            I => \testWordZ0Z_4\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__22476\,
            I => \testWordZ0Z_4\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__22473\,
            I => \testWordZ0Z_4\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__22468\,
            I => \testWordZ0Z_4\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__22463\,
            I => \testWordZ0Z_4\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__22460\,
            I => \testWordZ0Z_4\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__22457\,
            I => \testWordZ0Z_4\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__22442\,
            I => \N__22433\
        );

    \I__3687\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22423\
        );

    \I__3686\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22423\
        );

    \I__3685\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22423\
        );

    \I__3684\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22420\
        );

    \I__3683\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22410\
        );

    \I__3682\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22410\
        );

    \I__3681\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22410\
        );

    \I__3680\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22410\
        );

    \I__3679\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22397\
        );

    \I__3678\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22397\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__22423\,
            I => \N__22392\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22392\
        );

    \I__3675\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22389\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22382\
        );

    \I__3673\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22379\
        );

    \I__3672\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22376\
        );

    \I__3671\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22373\
        );

    \I__3670\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22366\
        );

    \I__3669\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22366\
        );

    \I__3668\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22366\
        );

    \I__3667\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22361\
        );

    \I__3666\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22361\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22354\
        );

    \I__3664\ : Span4Mux_h
    port map (
            O => \N__22392\,
            I => \N__22354\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__22389\,
            I => \N__22354\
        );

    \I__3662\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22345\
        );

    \I__3661\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22345\
        );

    \I__3660\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22345\
        );

    \I__3659\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22345\
        );

    \I__3658\ : Span12Mux_s1_v
    port map (
            O => \N__22382\,
            I => \N__22342\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__22379\,
            I => \testWordZ0Z_2\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__22376\,
            I => \testWordZ0Z_2\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__22373\,
            I => \testWordZ0Z_2\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__22366\,
            I => \testWordZ0Z_2\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__22361\,
            I => \testWordZ0Z_2\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__22354\,
            I => \testWordZ0Z_2\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__22345\,
            I => \testWordZ0Z_2\
        );

    \I__3650\ : Odrv12
    port map (
            O => \N__22342\,
            I => \testWordZ0Z_2\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__22325\,
            I => \N__22316\
        );

    \I__3648\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22307\
        );

    \I__3647\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22307\
        );

    \I__3646\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22307\
        );

    \I__3645\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22307\
        );

    \I__3644\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22300\
        );

    \I__3643\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22300\
        );

    \I__3642\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22300\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22286\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__22300\,
            I => \N__22286\
        );

    \I__3639\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22282\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__22298\,
            I => \N__22277\
        );

    \I__3637\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22267\
        );

    \I__3636\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22267\
        );

    \I__3635\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22267\
        );

    \I__3634\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22258\
        );

    \I__3633\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22258\
        );

    \I__3632\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22258\
        );

    \I__3631\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22258\
        );

    \I__3630\ : Span4Mux_s3_v
    port map (
            O => \N__22286\,
            I => \N__22252\
        );

    \I__3629\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22249\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__22282\,
            I => \N__22246\
        );

    \I__3627\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22241\
        );

    \I__3626\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22241\
        );

    \I__3625\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22232\
        );

    \I__3624\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22232\
        );

    \I__3623\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22232\
        );

    \I__3622\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22232\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__22267\,
            I => \N__22229\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__22258\,
            I => \N__22226\
        );

    \I__3619\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22219\
        );

    \I__3618\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22219\
        );

    \I__3617\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22219\
        );

    \I__3616\ : IoSpan4Mux
    port map (
            O => \N__22252\,
            I => \N__22216\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__22249\,
            I => \N__22213\
        );

    \I__3614\ : Span4Mux_s1_v
    port map (
            O => \N__22246\,
            I => \N__22204\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__22241\,
            I => \N__22204\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__22232\,
            I => \N__22204\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__22229\,
            I => \N__22204\
        );

    \I__3610\ : Span4Mux_v
    port map (
            O => \N__22226\,
            I => \N__22200\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__22219\,
            I => \N__22197\
        );

    \I__3608\ : Span4Mux_s0_h
    port map (
            O => \N__22216\,
            I => \N__22192\
        );

    \I__3607\ : Span4Mux_h
    port map (
            O => \N__22213\,
            I => \N__22192\
        );

    \I__3606\ : Span4Mux_h
    port map (
            O => \N__22204\,
            I => \N__22189\
        );

    \I__3605\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22186\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__22200\,
            I => \N__22181\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__22197\,
            I => \N__22181\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__22192\,
            I => \N__22178\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__22189\,
            I => \N__22175\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__22186\,
            I => \testWordZ0Z_3\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__22181\,
            I => \testWordZ0Z_3\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__22178\,
            I => \testWordZ0Z_3\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__22175\,
            I => \testWordZ0Z_3\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__22166\,
            I => \ALU.N_469_cascade_\
        );

    \I__3595\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__22160\,
            I => \ALU.N_473\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__22157\,
            I => \ALU.rshift_15_ns_1_1_cascade_\
        );

    \I__3592\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22151\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__22142\,
            I => \N_305_0\
        );

    \I__3587\ : CEMux
    port map (
            O => \N__22139\,
            I => \N__22134\
        );

    \I__3586\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22131\
        );

    \I__3585\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22128\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__22134\,
            I => \N__22125\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__22131\,
            I => \N__22121\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22118\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__22125\,
            I => \N__22115\
        );

    \I__3580\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22112\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__22121\,
            I => \N__22107\
        );

    \I__3578\ : Span4Mux_s2_v
    port map (
            O => \N__22118\,
            I => \N__22107\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__22115\,
            I => \CONTROL.aluParams_cnvZ0Z_0\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__22112\,
            I => \CONTROL.aluParams_cnvZ0Z_0\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__22107\,
            I => \CONTROL.aluParams_cnvZ0Z_0\
        );

    \I__3574\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__22097\,
            I => \ALU.a4_b_4\
        );

    \I__3572\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__22091\,
            I => \ALU.a3_b_5\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__22088\,
            I => \ALU.a4_b_4_cascade_\
        );

    \I__3569\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__22076\,
            I => \ALU.madd_98\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__22073\,
            I => \N__22069\
        );

    \I__3564\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22061\
        );

    \I__3563\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22058\
        );

    \I__3562\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22054\
        );

    \I__3561\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22049\
        );

    \I__3560\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22049\
        );

    \I__3559\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22044\
        );

    \I__3558\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22041\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22036\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22036\
        );

    \I__3555\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22033\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__22054\,
            I => \N__22030\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22027\
        );

    \I__3552\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22022\
        );

    \I__3551\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22022\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__22044\,
            I => \N__22019\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__22014\
        );

    \I__3548\ : Span4Mux_v
    port map (
            O => \N__22036\,
            I => \N__22014\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__22033\,
            I => \N__22007\
        );

    \I__3546\ : Span4Mux_v
    port map (
            O => \N__22030\,
            I => \N__22007\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__22027\,
            I => \N__22007\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__22022\,
            I => \N__22004\
        );

    \I__3543\ : Span4Mux_v
    port map (
            O => \N__22019\,
            I => \N__21997\
        );

    \I__3542\ : Span4Mux_v
    port map (
            O => \N__22014\,
            I => \N__21997\
        );

    \I__3541\ : Span4Mux_v
    port map (
            O => \N__22007\,
            I => \N__21992\
        );

    \I__3540\ : Span4Mux_h
    port map (
            O => \N__22004\,
            I => \N__21992\
        );

    \I__3539\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21987\
        );

    \I__3538\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21987\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__21997\,
            I => \ALU.N_207_0\
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__21992\,
            I => \ALU.N_207_0\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__21987\,
            I => \ALU.N_207_0\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__21980\,
            I => \ALU.madd_98_cascade_\
        );

    \I__3533\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21970\
        );

    \I__3531\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21967\
        );

    \I__3530\ : Span4Mux_s3_h
    port map (
            O => \N__21970\,
            I => \N__21964\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__21967\,
            I => \N__21961\
        );

    \I__3528\ : Sp12to4
    port map (
            O => \N__21964\,
            I => \N__21958\
        );

    \I__3527\ : Span4Mux_h
    port map (
            O => \N__21961\,
            I => \N__21955\
        );

    \I__3526\ : Odrv12
    port map (
            O => \N__21958\,
            I => \ALU.madd_93\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__21955\,
            I => \ALU.madd_93\
        );

    \I__3524\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21941\
        );

    \I__3523\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21941\
        );

    \I__3522\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21941\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__21941\,
            I => \ALU.madd_139\
        );

    \I__3520\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21931\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__21934\,
            I => \N__21928\
        );

    \I__3517\ : Span4Mux_v
    port map (
            O => \N__21931\,
            I => \N__21925\
        );

    \I__3516\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21922\
        );

    \I__3515\ : Span4Mux_h
    port map (
            O => \N__21925\,
            I => \N__21917\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__21922\,
            I => \N__21917\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__3512\ : Span4Mux_h
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__3510\ : Span4Mux_h
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__21905\,
            I => \RX_c\
        );

    \I__3508\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__3506\ : Span4Mux_v
    port map (
            O => \N__21896\,
            I => \N__21892\
        );

    \I__3505\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21889\
        );

    \I__3504\ : Span4Mux_v
    port map (
            O => \N__21892\,
            I => \N__21884\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21880\
        );

    \I__3502\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21875\
        );

    \I__3501\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21875\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__21884\,
            I => \N__21872\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21869\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__21880\,
            I => \RXready\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__21875\,
            I => \RXready\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__21872\,
            I => \RXready\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__21869\,
            I => \RXready\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__21860\,
            I => \N__21856\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__21859\,
            I => \N__21853\
        );

    \I__3492\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21850\
        );

    \I__3491\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21847\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21843\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21840\
        );

    \I__3488\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21837\
        );

    \I__3487\ : Span12Mux_s3_v
    port map (
            O => \N__21843\,
            I => \N__21834\
        );

    \I__3486\ : Span4Mux_h
    port map (
            O => \N__21840\,
            I => \N__21831\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__21837\,
            I => \ctrlOut_1\
        );

    \I__3484\ : Odrv12
    port map (
            O => \N__21834\,
            I => \ctrlOut_1\
        );

    \I__3483\ : Odrv4
    port map (
            O => \N__21831\,
            I => \ctrlOut_1\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__21824\,
            I => \ALU.N_41_0_0_cascade_\
        );

    \I__3481\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__21818\,
            I => \ALU.rshift_3_ns_1_5\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__21815\,
            I => \ALU.N_752_cascade_\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__21812\,
            I => \ALU.dout_3_ns_1_5_cascade_\
        );

    \I__3477\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__21806\,
            I => \ALU.N_704\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__21803\,
            I => \ALU.un2_addsub_axb_4_cascade_\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__3473\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__3471\ : Odrv12
    port map (
            O => \N__21791\,
            I => \ALU.d_RNI312TBZ0Z_4\
        );

    \I__3470\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21781\
        );

    \I__3469\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21776\
        );

    \I__3468\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21776\
        );

    \I__3467\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21773\
        );

    \I__3466\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21770\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__21781\,
            I => \N__21767\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21762\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21759\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__21770\,
            I => \N__21754\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__21767\,
            I => \N__21754\
        );

    \I__3460\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21749\
        );

    \I__3459\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21749\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__21762\,
            I => \N__21746\
        );

    \I__3457\ : Span4Mux_h
    port map (
            O => \N__21759\,
            I => \N__21739\
        );

    \I__3456\ : Span4Mux_h
    port map (
            O => \N__21754\,
            I => \N__21739\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21739\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__21746\,
            I => \N__21736\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__21739\,
            I => \N__21733\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__21736\,
            I => \ALU.N_223_0\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__21733\,
            I => \ALU.N_223_0\
        );

    \I__3450\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21718\
        );

    \I__3448\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21715\
        );

    \I__3447\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21710\
        );

    \I__3446\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21710\
        );

    \I__3445\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21707\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__21718\,
            I => \N__21704\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21701\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21696\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__21707\,
            I => \N__21693\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__21704\,
            I => \N__21688\
        );

    \I__3439\ : Span4Mux_v
    port map (
            O => \N__21701\,
            I => \N__21688\
        );

    \I__3438\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21683\
        );

    \I__3437\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21683\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__21696\,
            I => \ALU.operand2_5\
        );

    \I__3435\ : Odrv12
    port map (
            O => \N__21693\,
            I => \ALU.operand2_5\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__21688\,
            I => \ALU.operand2_5\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__21683\,
            I => \ALU.operand2_5\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__21674\,
            I => \ALU.a3_b_5_cascade_\
        );

    \I__3431\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21665\
        );

    \I__3430\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21665\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__3428\ : Odrv12
    port map (
            O => \N__21662\,
            I => \ALU.madd_94\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__21659\,
            I => \ALU.g_RNIT0COZ0Z_1_cascade_\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__21656\,
            I => \ALU.operand2_7_ns_1_1_cascade_\
        );

    \I__3425\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__21647\,
            I => \ALU.e_RNIPKVJZ0Z_1\
        );

    \I__3422\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__21638\,
            I => \ALU.madd_4\
        );

    \I__3419\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__21629\,
            I => \ALU.madd_12_0_tz\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \ALU.dout_6_ns_1_15_cascade_\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__21623\,
            I => \ALU.N_747_cascade_\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__21620\,
            I => \ALU.aluOut_0_cascade_\
        );

    \I__3413\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__3411\ : Span4Mux_s2_h
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__3409\ : Span4Mux_h
    port map (
            O => \N__21605\,
            I => \N__21602\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__21602\,
            I => \ALU.g0_0_0_N_2L1\
        );

    \I__3407\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21596\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__21596\,
            I => \ALU.dout_3_ns_1_7\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__3404\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__3402\ : Odrv12
    port map (
            O => \N__21584\,
            I => \ALU.a_15_m5_0\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__21581\,
            I => \ALU.d_RNI9BO713Z0Z_0_cascade_\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__21578\,
            I => \ALU.operand2_7_ns_1_0_cascade_\
        );

    \I__3399\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21569\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__21569\,
            I => \N__21565\
        );

    \I__3396\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21560\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__21565\,
            I => \N__21557\
        );

    \I__3394\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21554\
        );

    \I__3393\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21551\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21546\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__21557\,
            I => \N__21546\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__21554\,
            I => \ctrlOut_0\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__21551\,
            I => \ctrlOut_0\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__21546\,
            I => \ctrlOut_0\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__21539\,
            I => \ALU.operand2_0_cascade_\
        );

    \I__3386\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21532\
        );

    \I__3385\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21529\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__21532\,
            I => \ALU.hZ0Z_0\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__21529\,
            I => \ALU.hZ0Z_0\
        );

    \I__3382\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21521\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__21521\,
            I => \ALU.d_RNIE4R7Z0Z_0\
        );

    \I__3380\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21515\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__21515\,
            I => \ALU.g0_7_a3_0Z0Z_0\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__21512\,
            I => \ALU.N_8_1_cascade_\
        );

    \I__3377\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__21506\,
            I => \ALU.g0_2Z0Z_1\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__21503\,
            I => \ALU.g0_7_m4_0_1_cascade_\
        );

    \I__3374\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__21497\,
            I => \ALU.N_9_2\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__21494\,
            I => \ALU.dout_3_ns_1_0_cascade_\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__21491\,
            I => \ALU.dout_6_ns_1_0_cascade_\
        );

    \I__3370\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21481\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__21487\,
            I => \N__21478\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__21486\,
            I => \N__21475\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__21485\,
            I => \N__21472\
        );

    \I__3366\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21466\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21463\
        );

    \I__3364\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21460\
        );

    \I__3363\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21457\
        );

    \I__3362\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21454\
        );

    \I__3361\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21451\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21448\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__21469\,
            I => \N__21445\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__21466\,
            I => \N__21441\
        );

    \I__3357\ : Span4Mux_v
    port map (
            O => \N__21463\,
            I => \N__21438\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__21460\,
            I => \N__21431\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21431\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__21454\,
            I => \N__21431\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__21451\,
            I => \N__21428\
        );

    \I__3352\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21421\
        );

    \I__3351\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21421\
        );

    \I__3350\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21421\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__21441\,
            I => \N__21416\
        );

    \I__3348\ : Span4Mux_h
    port map (
            O => \N__21438\,
            I => \N__21416\
        );

    \I__3347\ : Span4Mux_v
    port map (
            O => \N__21431\,
            I => \N__21413\
        );

    \I__3346\ : Odrv12
    port map (
            O => \N__21428\,
            I => \ALU.N_201_0\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__21421\,
            I => \ALU.N_201_0\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__21416\,
            I => \ALU.N_201_0\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__21413\,
            I => \ALU.N_201_0\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__3341\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__21398\,
            I => \N__21395\
        );

    \I__3339\ : Span4Mux_h
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__3338\ : Span4Mux_v
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__21389\,
            I => \ALU.d_RNIQ74VBZ0Z_8\
        );

    \I__3336\ : InMux
    port map (
            O => \N__21386\,
            I => \bfn_6_10_0_\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__3334\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21377\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__21377\,
            I => \N__21374\
        );

    \I__3332\ : Span12Mux_h
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__3331\ : Odrv12
    port map (
            O => \N__21371\,
            I => \ALU.d_RNI6B7KDZ0Z_9\
        );

    \I__3330\ : InMux
    port map (
            O => \N__21368\,
            I => \ALU.un2_addsub_cry_8\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__3328\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__21350\,
            I => \ALU.N_192_0_i\
        );

    \I__3323\ : InMux
    port map (
            O => \N__21347\,
            I => \ALU.un2_addsub_cry_9\
        );

    \I__3322\ : InMux
    port map (
            O => \N__21344\,
            I => \ALU.un2_addsub_cry_10\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__3320\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__3318\ : Span4Mux_h
    port map (
            O => \N__21332\,
            I => \N__21329\
        );

    \I__3317\ : Span4Mux_h
    port map (
            O => \N__21329\,
            I => \N__21326\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__21323\,
            I => \ALU.N_180_0_i\
        );

    \I__3314\ : InMux
    port map (
            O => \N__21320\,
            I => \ALU.un2_addsub_cry_11\
        );

    \I__3313\ : InMux
    port map (
            O => \N__21317\,
            I => \ALU.un2_addsub_cry_12\
        );

    \I__3312\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21308\
        );

    \I__3311\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21305\
        );

    \I__3310\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21301\
        );

    \I__3309\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21298\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21291\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21291\
        );

    \I__3306\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21288\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__21301\,
            I => \N__21285\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21282\
        );

    \I__3303\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21277\
        );

    \I__3302\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21277\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__21291\,
            I => \N__21274\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__21288\,
            I => \ALU.N_171_0\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__21285\,
            I => \ALU.N_171_0\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__21282\,
            I => \ALU.N_171_0\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__21277\,
            I => \ALU.N_171_0\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__21274\,
            I => \ALU.N_171_0\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__3294\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__3291\ : Span4Mux_v
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__21248\,
            I => \ALU.d_RNI1M3JEZ0Z_14\
        );

    \I__3289\ : InMux
    port map (
            O => \N__21245\,
            I => \ALU.un2_addsub_cry_13\
        );

    \I__3288\ : InMux
    port map (
            O => \N__21242\,
            I => \ALU.un2_addsub_cry_14\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__3286\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21227\
        );

    \I__3285\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21227\
        );

    \I__3284\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21227\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__3282\ : Span4Mux_v
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__21218\,
            I => \ALU.a0_b_11\
        );

    \I__3279\ : InMux
    port map (
            O => \N__21215\,
            I => \ALU.un2_addsub_cry_0\
        );

    \I__3278\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__21209\,
            I => \N__21206\
        );

    \I__3276\ : Sp12to4
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__3275\ : Span12Mux_s4_h
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__3274\ : Odrv12
    port map (
            O => \N__21200\,
            I => \ALU.d_RNIEDJEAZ0Z_2\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__3272\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__21188\,
            I => \N__21185\
        );

    \I__3269\ : Span4Mux_h
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__21182\,
            I => \ALU.N_240_0_i\
        );

    \I__3267\ : InMux
    port map (
            O => \N__21179\,
            I => \ALU.un2_addsub_cry_1\
        );

    \I__3266\ : InMux
    port map (
            O => \N__21176\,
            I => \ALU.un2_addsub_cry_2\
        );

    \I__3265\ : InMux
    port map (
            O => \N__21173\,
            I => \ALU.un2_addsub_cry_3\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__21170\,
            I => \N__21167\
        );

    \I__3263\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__3261\ : Span4Mux_h
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__3260\ : Span4Mux_v
    port map (
            O => \N__21158\,
            I => \N__21155\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__21155\,
            I => \ALU.d_RNIVR3QAZ0Z_5\
        );

    \I__3258\ : InMux
    port map (
            O => \N__21152\,
            I => \ALU.un2_addsub_cry_4\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__3256\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__3254\ : Span4Mux_v
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__3253\ : Span4Mux_v
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__3252\ : Span4Mux_h
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__21131\,
            I => \ALU.d_RNIGLK5BZ0Z_6\
        );

    \I__3250\ : InMux
    port map (
            O => \N__21128\,
            I => \ALU.un2_addsub_cry_5\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__3248\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__3245\ : Span4Mux_h
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__3244\ : Span4Mux_s1_h
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__21104\,
            I => \ALU.d_RNITAM9DZ0Z_7\
        );

    \I__3241\ : InMux
    port map (
            O => \N__21101\,
            I => \ALU.un2_addsub_cry_6\
        );

    \I__3240\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21090\
        );

    \I__3239\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21086\
        );

    \I__3238\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21083\
        );

    \I__3237\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21076\
        );

    \I__3236\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21076\
        );

    \I__3235\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21076\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__21090\,
            I => \N__21073\
        );

    \I__3233\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21070\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__21086\,
            I => \N__21067\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21064\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__21076\,
            I => \N__21061\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__21073\,
            I => \N__21058\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__21070\,
            I => \N__21054\
        );

    \I__3227\ : Span4Mux_v
    port map (
            O => \N__21067\,
            I => \N__21049\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__21064\,
            I => \N__21049\
        );

    \I__3225\ : Span4Mux_h
    port map (
            O => \N__21061\,
            I => \N__21044\
        );

    \I__3224\ : Span4Mux_h
    port map (
            O => \N__21058\,
            I => \N__21044\
        );

    \I__3223\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21041\
        );

    \I__3222\ : Odrv12
    port map (
            O => \N__21054\,
            I => \ALU.N_205_0\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__21049\,
            I => \ALU.N_205_0\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__21044\,
            I => \ALU.N_205_0\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__21041\,
            I => \ALU.N_205_0\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__21032\,
            I => \ALU.operand2_9_cascade_\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__21029\,
            I => \ALU.a_15_m2_ns_1Z0Z_9_cascade_\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__21026\,
            I => \ALU.d_RNIO7LUZ0Z_13_cascade_\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__21023\,
            I => \ALU.operand2_13_cascade_\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__21020\,
            I => \ALU.N_177_0_cascade_\
        );

    \I__3213\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21014\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__3211\ : Odrv12
    port map (
            O => \N__21011\,
            I => \ALU.madd_484_3\
        );

    \I__3210\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__3208\ : Span4Mux_v
    port map (
            O => \N__21002\,
            I => \N__20999\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__20999\,
            I => \ALU.madd_484_1\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__20996\,
            I => \ALU.madd_484_2_cascade_\
        );

    \I__3205\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__20987\,
            I => \ALU.madd_484_0\
        );

    \I__3202\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20978\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__20978\,
            I => \ALU.madd_484_12\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \ALU.m270_nsZ0Z_1_cascade_\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__20972\,
            I => \N__20967\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__20971\,
            I => \N__20963\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__20970\,
            I => \N__20960\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20957\
        );

    \I__3194\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20950\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20950\
        );

    \I__3192\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20950\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__20957\,
            I => \ctrlOut_12\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__20950\,
            I => \ctrlOut_12\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__20945\,
            I => \N__20941\
        );

    \I__3188\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20937\
        );

    \I__3187\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20934\
        );

    \I__3186\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20931\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20926\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20926\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__20931\,
            I => \ctrlOut_15\
        );

    \I__3182\ : Odrv12
    port map (
            O => \N__20926\,
            I => \ctrlOut_15\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__20921\,
            I => \ALU.N_7_0_cascade_\
        );

    \I__3180\ : InMux
    port map (
            O => \N__20918\,
            I => \N__20908\
        );

    \I__3179\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20908\
        );

    \I__3178\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20908\
        );

    \I__3177\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20905\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__20908\,
            I => \N__20902\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__20905\,
            I => \N__20899\
        );

    \I__3174\ : Sp12to4
    port map (
            O => \N__20902\,
            I => \N__20896\
        );

    \I__3173\ : Span4Mux_v
    port map (
            O => \N__20899\,
            I => \N__20891\
        );

    \I__3172\ : Span12Mux_s5_h
    port map (
            O => \N__20896\,
            I => \N__20888\
        );

    \I__3171\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20885\
        );

    \I__3170\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20882\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__20891\,
            I => \ALU.N_179_0\
        );

    \I__3168\ : Odrv12
    port map (
            O => \N__20888\,
            I => \ALU.N_179_0\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__20885\,
            I => \ALU.N_179_0\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__20882\,
            I => \ALU.N_179_0\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__20873\,
            I => \ALU.a_15_m2_ns_1Z0Z_13_cascade_\
        );

    \I__3164\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20861\
        );

    \I__3163\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20861\
        );

    \I__3162\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20858\
        );

    \I__3161\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20855\
        );

    \I__3160\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20852\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__20861\,
            I => \N__20849\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__20858\,
            I => \N__20846\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__20855\,
            I => \N__20843\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__20852\,
            I => \N__20840\
        );

    \I__3155\ : Span4Mux_v
    port map (
            O => \N__20849\,
            I => \N__20833\
        );

    \I__3154\ : Span4Mux_s2_h
    port map (
            O => \N__20846\,
            I => \N__20833\
        );

    \I__3153\ : Span4Mux_v
    port map (
            O => \N__20843\,
            I => \N__20833\
        );

    \I__3152\ : Span4Mux_h
    port map (
            O => \N__20840\,
            I => \N__20830\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__20833\,
            I => \ALU.operand2_9\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__20830\,
            I => \ALU.operand2_9\
        );

    \I__3149\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__20822\,
            I => \ALU.N_220\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__3146\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__20813\,
            I => \ALU.N_250\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__20810\,
            I => \ALU.N_250_cascade_\
        );

    \I__3143\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__20804\,
            I => \ALU.N_254\
        );

    \I__3141\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__20798\,
            I => \ALU.N_218\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__20795\,
            I => \ALU.N_218_cascade_\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__20792\,
            I => \ALU.N_361_cascade_\
        );

    \I__3137\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20785\
        );

    \I__3136\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20782\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__20785\,
            I => \ALU.N_252\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__20782\,
            I => \ALU.N_252\
        );

    \I__3133\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__20774\,
            I => \ALU.N_257\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__20771\,
            I => \ALU.N_249_cascade_\
        );

    \I__3130\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20762\
        );

    \I__3129\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20762\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__20762\,
            I => \ALU.N_253\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__20759\,
            I => \ALU.c_RNIUGCLVZ0Z_11_cascade_\
        );

    \I__3126\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20752\
        );

    \I__3125\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20749\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__20752\,
            I => \ALU.N_415\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__20749\,
            I => \ALU.N_415\
        );

    \I__3122\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20741\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__20741\,
            I => \ALU.N_310\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__20738\,
            I => \ALU.lshift_3_ns_1_4_cascade_\
        );

    \I__3119\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__3117\ : Span4Mux_h
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__20723\,
            I => \ALU.N_273_0\
        );

    \I__3114\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__20717\,
            I => \ALU.N_461\
        );

    \I__3112\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20708\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__20708\,
            I => \ALU.N_474\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__20705\,
            I => \ALU.N_530_cascade_\
        );

    \I__3108\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20696\
        );

    \I__3107\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20696\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__20696\,
            I => \ALU.N_635\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__20693\,
            I => \ALU.d_RNIP8ITN1Z0Z_5_cascade_\
        );

    \I__3104\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__20687\,
            I => \N__20684\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__20684\,
            I => \ALU.d_RNILBFG4Z0Z_2\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__20681\,
            I => \ALU.a_15_m3_2_cascade_\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__20678\,
            I => \ALU.d_RNIE937BZ0Z_0_cascade_\
        );

    \I__3099\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__20672\,
            I => \ALU.a_15_m4_2\
        );

    \I__3097\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20663\
        );

    \I__3096\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20663\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__20663\,
            I => \FTDI.N_28\
        );

    \I__3094\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__20657\,
            I => \ALU.a_15_m1_0\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \ALU.a_15_m4_ns_1_0_cascade_\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__20651\,
            I => \ALU.a_15_m4_0_cascade_\
        );

    \I__3090\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__20645\,
            I => \ALU.a_15_m3_0\
        );

    \I__3088\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20639\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__20636\,
            I => \N__20633\
        );

    \I__3085\ : Span4Mux_v
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__3084\ : Span4Mux_s1_v
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__20627\,
            I => \ALU.a_15_m4_bm_1Z0Z_8\
        );

    \I__3082\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__20621\,
            I => \ALU.a_15_m0_0\
        );

    \I__3080\ : InMux
    port map (
            O => \N__20618\,
            I => \N__20615\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__20609\,
            I => i53_mux_0
        );

    \I__3076\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__20603\,
            I => \ALU.madd_33\
        );

    \I__3074\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__20597\,
            I => \ALU.madd_68_0_tz\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__20591\,
            I => \ALU.madd_68\
        );

    \I__3070\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20582\
        );

    \I__3069\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20582\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20579\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__20579\,
            I => \ALU.madd_89_0\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__20576\,
            I => \ALU.madd_68_cascade_\
        );

    \I__3065\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20567\
        );

    \I__3064\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20567\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__20567\,
            I => \N__20563\
        );

    \I__3062\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20560\
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__20563\,
            I => \ALU.a7_b_1\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__20560\,
            I => \ALU.a7_b_1\
        );

    \I__3059\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20549\
        );

    \I__3058\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20549\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__20549\,
            I => \ALU.madd_108\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__20546\,
            I => \ALU.madd_108_cascade_\
        );

    \I__3055\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20534\
        );

    \I__3054\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20534\
        );

    \I__3053\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20534\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__3051\ : Span4Mux_h
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__20528\,
            I => \ALU.madd_134\
        );

    \I__3049\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20519\
        );

    \I__3048\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20519\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20516\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__20513\,
            I => \ALU.madd_153\
        );

    \I__3044\ : CEMux
    port map (
            O => \N__20510\,
            I => \N__20506\
        );

    \I__3043\ : CEMux
    port map (
            O => \N__20509\,
            I => \N__20503\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20500\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__20503\,
            I => \N__20497\
        );

    \I__3040\ : Span4Mux_s1_h
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__3039\ : Span12Mux_v
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__3038\ : Span4Mux_h
    port map (
            O => \N__20494\,
            I => \N__20488\
        );

    \I__3037\ : Odrv12
    port map (
            O => \N__20491\,
            I => \FTDI.N_201_2\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__20488\,
            I => \FTDI.N_201_2\
        );

    \I__3035\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__20480\,
            I => \N__20475\
        );

    \I__3033\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20472\
        );

    \I__3032\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20469\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__20475\,
            I => \aluOperation_3\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__20472\,
            I => \aluOperation_3\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__20469\,
            I => \aluOperation_3\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__20462\,
            I => \ALU.m681Z0Z_1_cascade_\
        );

    \I__3027\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20450\
        );

    \I__3026\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20445\
        );

    \I__3025\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20445\
        );

    \I__3024\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20436\
        );

    \I__3023\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20436\
        );

    \I__3022\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20436\
        );

    \I__3021\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20436\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20428\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20428\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20428\
        );

    \I__3017\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20425\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__20428\,
            I => \N__20420\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__20425\,
            I => \N__20420\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__20420\,
            I => \ALU.N_730_mux\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__20417\,
            I => \ALU.a7_b_0_cascade_\
        );

    \I__3012\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__20408\,
            I => \N__20404\
        );

    \I__3009\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__20404\,
            I => \ALU.madd_59\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__20401\,
            I => \ALU.madd_59\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__3005\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__3001\ : Span4Mux_h
    port map (
            O => \N__20381\,
            I => \N__20378\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__20378\,
            I => \ALU.madd_484_5\
        );

    \I__2999\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20372\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__2997\ : Odrv12
    port map (
            O => \N__20369\,
            I => \ALU.madd_128_0_tz_0\
        );

    \I__2996\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20360\
        );

    \I__2995\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20360\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__2993\ : Odrv12
    port map (
            O => \N__20357\,
            I => \ALU.madd_104\
        );

    \I__2992\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__2990\ : Span12Mux_s4_h
    port map (
            O => \N__20348\,
            I => \N__20344\
        );

    \I__2989\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20341\
        );

    \I__2988\ : Odrv12
    port map (
            O => \N__20344\,
            I => \ALU.madd_149\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__20341\,
            I => \ALU.madd_149\
        );

    \I__2986\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__20333\,
            I => \ALU.madd_128_0_tz\
        );

    \I__2984\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20324\
        );

    \I__2983\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20324\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__20321\,
            I => \ALU.madd_128_0\
        );

    \I__2980\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__2978\ : Span4Mux_h
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__20309\,
            I => \ALU.madd_N_1_i\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__20306\,
            I => \ALU.madd_20_0_cascade_\
        );

    \I__2975\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20294\
        );

    \I__2974\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20294\
        );

    \I__2973\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20294\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__20294\,
            I => \ALU.madd_20\
        );

    \I__2971\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20286\
        );

    \I__2970\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20281\
        );

    \I__2969\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20281\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__20286\,
            I => \N__20278\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20273\
        );

    \I__2966\ : Span12Mux_s9_h
    port map (
            O => \N__20278\,
            I => \N__20270\
        );

    \I__2965\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20265\
        );

    \I__2964\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20265\
        );

    \I__2963\ : Span4Mux_v
    port map (
            O => \N__20273\,
            I => \N__20262\
        );

    \I__2962\ : Span12Mux_v
    port map (
            O => \N__20270\,
            I => \N__20259\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__20265\,
            I => \ctrlOut_2\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__20262\,
            I => \ctrlOut_2\
        );

    \I__2959\ : Odrv12
    port map (
            O => \N__20259\,
            I => \ctrlOut_2\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__20252\,
            I => \ALU.N_5_0_cascade_\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__20249\,
            I => \ALU.N_240_0_cascade_\
        );

    \I__2956\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__20243\,
            I => \ALU.madd_24_0_tz\
        );

    \I__2954\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__2952\ : Span4Mux_h
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__20231\,
            I => \ALU.madd_8_0\
        );

    \I__2950\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__2948\ : Span4Mux_h
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__20219\,
            I => \ALU.madd_5\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__20216\,
            I => \ALU.madd_8_0_cascade_\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__20213\,
            I => \ALU.N_706_cascade_\
        );

    \I__2944\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__20207\,
            I => \ALU.N_754\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__20204\,
            I => \ALU.aluOut_7_cascade_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20198\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__2939\ : Span4Mux_h
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__2938\ : Span4Mux_v
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__20189\,
            I => \ALU.a7_b_0_6\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2935\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__20174\,
            I => \ALU.m271_nsZ0Z_1\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__20171\,
            I => \ALU.N_708_cascade_\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__20168\,
            I => \ALU.dout_6_ns_1_9_cascade_\
        );

    \I__2929\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20162\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__20162\,
            I => \ALU.N_756\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__20159\,
            I => \ALU.N_751_cascade_\
        );

    \I__2926\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__20153\,
            I => \ALU.N_703\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__20150\,
            I => \ALU.rshift_3_ns_1_4_cascade_\
        );

    \I__2923\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__2921\ : Span12Mux_s11_v
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__2920\ : Odrv12
    port map (
            O => \N__20138\,
            I => \ALU.N_472\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__20135\,
            I => \ALU.N_472_cascade_\
        );

    \I__2918\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__2916\ : Span4Mux_v
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__2915\ : Span4Mux_v
    port map (
            O => \N__20123\,
            I => \N__20119\
        );

    \I__2914\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20116\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__20119\,
            I => \ALU.N_476\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__20116\,
            I => \ALU.N_476\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__20111\,
            I => \ALU.m272_nsZ0Z_1_cascade_\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__2909\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__2907\ : Span4Mux_v
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__20093\,
            I => \ALU.N_191_0_0\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \N__20084\
        );

    \I__2903\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20069\
        );

    \I__2902\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20069\
        );

    \I__2901\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20069\
        );

    \I__2900\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20069\
        );

    \I__2899\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20069\
        );

    \I__2898\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20069\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__20069\,
            I => \ctrlOut_10\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__20066\,
            I => \N__20062\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__20065\,
            I => \N__20059\
        );

    \I__2894\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20054\
        );

    \I__2893\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20054\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__2890\ : IoSpan4Mux
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__2889\ : Span4Mux_s2_h
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__20042\,
            I => \N__20037\
        );

    \I__2887\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20032\
        );

    \I__2886\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20032\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__20037\,
            I => \ALU.N_191_0\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__20032\,
            I => \ALU.N_191_0\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \ALU.N_191_0_cascade_\
        );

    \I__2882\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20015\
        );

    \I__2881\ : InMux
    port map (
            O => \N__20023\,
            I => \N__20015\
        );

    \I__2880\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20015\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__20010\
        );

    \I__2878\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20007\
        );

    \I__2877\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20004\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__20010\,
            I => \ALU.operand2_10\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__20007\,
            I => \ALU.operand2_10\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__20004\,
            I => \ALU.operand2_10\
        );

    \I__2873\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__2871\ : Span4Mux_s3_h
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__19988\,
            I => \ALU.a1_b_10\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__19985\,
            I => \ALU.a1_b_10_cascade_\
        );

    \I__2868\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19975\
        );

    \I__2867\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19975\
        );

    \I__2866\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19972\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__19975\,
            I => \N__19969\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19964\
        );

    \I__2863\ : Span12Mux_v
    port map (
            O => \N__19969\,
            I => \N__19964\
        );

    \I__2862\ : Odrv12
    port map (
            O => \N__19964\,
            I => \ALU.madd_203\
        );

    \I__2861\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__19955\,
            I => \N__19951\
        );

    \I__2858\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__19951\,
            I => \ALU.a9_b_2\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__19948\,
            I => \ALU.a9_b_2\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__19943\,
            I => \ALU.dout_3_ns_1_9_cascade_\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \ALU.N_186_0_cascade_\
        );

    \I__2853\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__19934\,
            I => \ALU.a1_b_11\
        );

    \I__2851\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19925\
        );

    \I__2850\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19925\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__19925\,
            I => \ALU.a0_b_12\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__19922\,
            I => \ALU.a1_b_11_cascade_\
        );

    \I__2847\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19912\
        );

    \I__2845\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19909\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__19912\,
            I => \N__19904\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19904\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__19901\,
            I => \ALU.madd_255\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__19898\,
            I => \ALU.dout_6_ns_1_8_cascade_\
        );

    \I__2839\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__19892\,
            I => \ALU.dout_3_ns_1_8\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__19889\,
            I => \ALU.N_707_cascade_\
        );

    \I__2836\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__19883\,
            I => \ALU.N_755\
        );

    \I__2834\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__2832\ : Odrv12
    port map (
            O => \N__19874\,
            I => \ALU.N_283_0\
        );

    \I__2831\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__19868\,
            I => \N__19864\
        );

    \I__2829\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19861\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__19864\,
            I => \N__19858\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__19861\,
            I => \ctrlOut_7\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__19858\,
            I => \ctrlOut_7\
        );

    \I__2825\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__19850\,
            I => \N__19846\
        );

    \I__2823\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19843\
        );

    \I__2822\ : Span4Mux_v
    port map (
            O => \N__19846\,
            I => \N__19839\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19834\
        );

    \I__2820\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19831\
        );

    \I__2819\ : IoSpan4Mux
    port map (
            O => \N__19839\,
            I => \N__19828\
        );

    \I__2818\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19823\
        );

    \I__2817\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19823\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__19834\,
            I => \N__19816\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__19831\,
            I => \N__19813\
        );

    \I__2814\ : Span4Mux_s1_h
    port map (
            O => \N__19828\,
            I => \N__19808\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19808\
        );

    \I__2812\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19805\
        );

    \I__2811\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19802\
        );

    \I__2810\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19799\
        );

    \I__2809\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19796\
        );

    \I__2808\ : Span4Mux_s1_h
    port map (
            O => \N__19816\,
            I => \N__19789\
        );

    \I__2807\ : Span4Mux_h
    port map (
            O => \N__19813\,
            I => \N__19789\
        );

    \I__2806\ : Span4Mux_v
    port map (
            O => \N__19808\,
            I => \N__19789\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19785\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__19802\,
            I => \N__19778\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19778\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19778\
        );

    \I__2801\ : Span4Mux_v
    port map (
            O => \N__19789\,
            I => \N__19775\
        );

    \I__2800\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19772\
        );

    \I__2799\ : Span12Mux_s6_v
    port map (
            O => \N__19785\,
            I => \N__19767\
        );

    \I__2798\ : Span12Mux_v
    port map (
            O => \N__19778\,
            I => \N__19767\
        );

    \I__2797\ : Span4Mux_s1_h
    port map (
            O => \N__19775\,
            I => \N__19764\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__19772\,
            I => \ALU.N_211_0\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__19767\,
            I => \ALU.N_211_0\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__19764\,
            I => \ALU.N_211_0\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__2792\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__19748\,
            I => \N__19744\
        );

    \I__2789\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19741\
        );

    \I__2788\ : Span4Mux_h
    port map (
            O => \N__19744\,
            I => \N__19738\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__19741\,
            I => \ctrlOut_9\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__19738\,
            I => \ctrlOut_9\
        );

    \I__2785\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19727\
        );

    \I__2784\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19727\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__19721\,
            I => \ALU.madd_367\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__2779\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__19712\,
            I => \ALU.d_RNIRV558Z0Z_13\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__19709\,
            I => \ALU.d_RNIRV558Z0Z_13_cascade_\
        );

    \I__2776\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__19700\,
            I => \ALU.madd_371\
        );

    \I__2773\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19691\
        );

    \I__2772\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19691\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__19691\,
            I => \ALU.a2_b_12\
        );

    \I__2770\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__19685\,
            I => \N__19681\
        );

    \I__2768\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19678\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__19681\,
            I => \N__19672\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19672\
        );

    \I__2765\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19669\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__19672\,
            I => \ALU.madd_259\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__19669\,
            I => \ALU.madd_259\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \ALU.N_240_0_i_cascade_\
        );

    \I__2761\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19655\
        );

    \I__2760\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19655\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__19652\,
            I => \N__19648\
        );

    \I__2757\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__19648\,
            I => \ALU.N_9_0\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__19645\,
            I => \ALU.N_9_0\
        );

    \I__2754\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19634\
        );

    \I__2753\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19634\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__2751\ : Span4Mux_v
    port map (
            O => \N__19631\,
            I => \N__19627\
        );

    \I__2750\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19624\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__19627\,
            I => \N__19621\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__19624\,
            I => \N__19618\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__19621\,
            I => \ALU.N_10_0\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__19618\,
            I => \ALU.N_10_0\
        );

    \I__2745\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__19604\,
            I => \ALU.N_253_0\
        );

    \I__2741\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__2739\ : Span4Mux_s2_v
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__19592\,
            I => \ALU.d_RNIUV3H4Z0Z_0\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__19589\,
            I => \N__19585\
        );

    \I__2736\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19580\
        );

    \I__2735\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19580\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__19577\,
            I => \N__19572\
        );

    \I__2732\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19567\
        );

    \I__2731\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19567\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__19572\,
            I => \ALU.N_635_0\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__19567\,
            I => \ALU.N_635_0\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__2727\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19550\
        );

    \I__2726\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19550\
        );

    \I__2725\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19550\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__19541\,
            I => \N__19536\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__19540\,
            I => \N__19533\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__19539\,
            I => \N__19530\
        );

    \I__2718\ : Sp12to4
    port map (
            O => \N__19536\,
            I => \N__19527\
        );

    \I__2717\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19522\
        );

    \I__2716\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19522\
        );

    \I__2715\ : Span12Mux_s3_v
    port map (
            O => \N__19527\,
            I => \N__19519\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__19522\,
            I => \ALU.N_724\
        );

    \I__2713\ : Odrv12
    port map (
            O => \N__19519\,
            I => \ALU.N_724\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \ALU.N_220_cascade_\
        );

    \I__2711\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19507\
        );

    \I__2710\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__19507\,
            I => \ALU.N_222\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__19504\,
            I => \ALU.N_222\
        );

    \I__2707\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__19490\,
            I => \ALU.madd_484_4\
        );

    \I__2703\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__19484\,
            I => \ALU.N_241_0\
        );

    \I__2701\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__19478\,
            I => \ALU.lshift_3_ns_1_15\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__2698\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__19469\,
            I => \ALU.dout_3_ns_1_14\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__19466\,
            I => \ALU.lshift_3_ns_1_14_cascade_\
        );

    \I__2695\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__19460\,
            I => \ALU.N_256\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__19457\,
            I => \ALU.N_224_cascade_\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__19454\,
            I => \ALU.d_RNI8DL9U1Z0Z_3_cascade_\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__19451\,
            I => \ALU.N_221_cascade_\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__19448\,
            I => \ALU.N_588_cascade_\
        );

    \I__2689\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__19442\,
            I => \ALU.N_575\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__19439\,
            I => \ALU.N_575_cascade_\
        );

    \I__2686\ : InMux
    port map (
            O => \N__19436\,
            I => \N__19433\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__19433\,
            I => \ALU.rshift_3_ns_1_8\
        );

    \I__2684\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__2682\ : Span4Mux_s1_v
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__19421\,
            I => \ALU.m55_bmZ0\
        );

    \I__2680\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__2678\ : Odrv12
    port map (
            O => \N__19412\,
            I => \ALU.m55_amZ0\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \ALU.m650_nsZ0Z_1_cascade_\
        );

    \I__2676\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19400\
        );

    \I__2675\ : InMux
    port map (
            O => \N__19405\,
            I => \N__19400\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__19400\,
            I => \ALU.N_15_0\
        );

    \I__2673\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__19394\,
            I => \N_727\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__19391\,
            I => \ALU.N_577_cascade_\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \ALU.N_528_cascade_\
        );

    \I__2669\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__19379\,
            I => \N__19375\
        );

    \I__2666\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__19375\,
            I => \ALU.N_633\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__19372\,
            I => \ALU.N_633\
        );

    \I__2663\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__2661\ : Span4Mux_h
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__19358\,
            I => \ALU.madd_144\
        );

    \I__2659\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__2657\ : Span4Mux_s3_h
    port map (
            O => \N__19349\,
            I => \N__19345\
        );

    \I__2656\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19342\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__19345\,
            I => \ALU.madd_113\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__19342\,
            I => \ALU.madd_113\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__19337\,
            I => \ALU.madd_154_cascade_\
        );

    \I__2652\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19330\
        );

    \I__2651\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19327\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19322\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__19327\,
            I => \N__19322\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__19316\,
            I => \ALU.madd_99\
        );

    \I__2645\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__19310\,
            I => \ALU.madd_73\
        );

    \I__2643\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19303\
        );

    \I__2642\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19300\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__19303\,
            I => \ALU.madd_109\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__19300\,
            I => \ALU.madd_109\
        );

    \I__2639\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__19289\,
            I => \N__19285\
        );

    \I__2636\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19282\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__19285\,
            I => \ALU.madd_154\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__19282\,
            I => \ALU.madd_154\
        );

    \I__2633\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__19271\,
            I => \N__19266\
        );

    \I__2630\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19261\
        );

    \I__2629\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19261\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__19266\,
            I => \ALU.madd_118\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__19261\,
            I => \ALU.madd_118\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__2625\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__19247\,
            I => \ALU.m641_nsZ0Z_1\
        );

    \I__2622\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__2620\ : Span4Mux_s0_v
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__19235\,
            I => \ALU.m645_nsZ0Z_1\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \ALU.N_283_0_cascade_\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__19229\,
            I => \ALU.madd_74_0_cascade_\
        );

    \I__2616\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19220\
        );

    \I__2615\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19220\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__19220\,
            I => \ALU.madd_83\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__19217\,
            I => \N__19212\
        );

    \I__2612\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19207\
        );

    \I__2611\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19207\
        );

    \I__2610\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19204\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__19207\,
            I => \ALU.madd_46\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__19204\,
            I => \ALU.madd_46\
        );

    \I__2607\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19193\
        );

    \I__2606\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19193\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__19193\,
            I => \ALU.madd_69\
        );

    \I__2604\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__19187\,
            I => \ALU.madd_74_0\
        );

    \I__2602\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19180\
        );

    \I__2601\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19177\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__19180\,
            I => \ALU.madd_79_0\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__19177\,
            I => \ALU.madd_79_0\
        );

    \I__2598\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19164\
        );

    \I__2597\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19164\
        );

    \I__2596\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19159\
        );

    \I__2595\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19159\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__19164\,
            I => \N__19156\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__19159\,
            I => \ALU.madd_51\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__19156\,
            I => \ALU.madd_51\
        );

    \I__2591\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19144\
        );

    \I__2590\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19144\
        );

    \I__2589\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19141\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__19144\,
            I => \N__19136\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19136\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__19136\,
            I => \ALU.madd_58\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \ALU.madd_79_0_cascade_\
        );

    \I__2584\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__19127\,
            I => \ALU.madd_56\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__19124\,
            I => \ALU.madd_88_cascade_\
        );

    \I__2581\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__19118\,
            I => \ALU.madd_114\
        );

    \I__2579\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__19112\,
            I => \ALU.madd_41\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__19109\,
            I => \ALU.madd_73_cascade_\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__2575\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19099\
        );

    \I__2574\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19095\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__19092\
        );

    \I__2572\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19086\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__19095\,
            I => \N__19082\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__19092\,
            I => \N__19077\
        );

    \I__2569\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19074\
        );

    \I__2568\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19069\
        );

    \I__2567\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19069\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__19086\,
            I => \N__19066\
        );

    \I__2565\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19063\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19060\
        );

    \I__2563\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19055\
        );

    \I__2562\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19055\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__19077\,
            I => \ALU.operand2_7\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__19074\,
            I => \ALU.operand2_7\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__19069\,
            I => \ALU.operand2_7\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__19066\,
            I => \ALU.operand2_7\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__19063\,
            I => \ALU.operand2_7\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__19060\,
            I => \ALU.operand2_7\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__19055\,
            I => \ALU.operand2_7\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__2553\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19033\
        );

    \I__2552\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__19033\,
            I => \ALU.a0_b_7\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__19030\,
            I => \ALU.a0_b_7\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__19025\,
            I => \ALU.madd_12_cascade_\
        );

    \I__2548\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__19019\,
            I => \ALU.madd_34\
        );

    \I__2546\ : InMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__19010\,
            I => \ALU.madd_42\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__19007\,
            I => \ALU.madd_34_cascade_\
        );

    \I__2542\ : InMux
    port map (
            O => \N__19004\,
            I => \N__18997\
        );

    \I__2541\ : InMux
    port map (
            O => \N__19003\,
            I => \N__18997\
        );

    \I__2540\ : InMux
    port map (
            O => \N__19002\,
            I => \N__18994\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__18997\,
            I => \ALU.madd_37\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__18994\,
            I => \ALU.madd_37\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__18989\,
            I => \ALU.madd_56_cascade_\
        );

    \I__2536\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__18980\,
            I => \ALU.madd_52_0\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__18977\,
            I => \N__18973\
        );

    \I__2532\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18965\
        );

    \I__2531\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18965\
        );

    \I__2530\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18965\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__18959\,
            I => \ALU.madd_25\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__2525\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18947\
        );

    \I__2524\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18947\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__18947\,
            I => \ALU.madd_12\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__18944\,
            I => \ALU.un2_addsub_axb_6_cascade_\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18936\
        );

    \I__2520\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18931\
        );

    \I__2519\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18931\
        );

    \I__2518\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18928\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__2514\ : Span4Mux_h
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__18919\,
            I => \ALU.madd_64_0\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__18916\,
            I => \ALU.madd_64_0\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__18911\,
            I => \ALU.a8_b_0_cascade_\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__18908\,
            I => \ALU.madd_10_cascade_\
        );

    \I__2509\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__18899\,
            I => \ALU.madd_24\
        );

    \I__2506\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__18887\,
            I => \ALU.madd_29\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__18884\,
            I => \ALU.madd_24_cascade_\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__2500\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__18875\,
            I => \ALU.madd_i1_mux_1\
        );

    \I__2498\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__18866\,
            I => \ALU.madd_i3_mux_0\
        );

    \I__2495\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18859\
        );

    \I__2494\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18856\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__18859\,
            I => \N__18853\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__18856\,
            I => \ALU.a4_b_2\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__18853\,
            I => \ALU.a4_b_2\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__2489\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__18842\,
            I => \ALU.a6_b_0\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__18839\,
            I => \ALU.operand2_10_cascade_\
        );

    \I__2486\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18830\
        );

    \I__2485\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18830\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__2483\ : Span4Mux_s3_h
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__18821\,
            I => \ALU.a4_b_10\
        );

    \I__2480\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__18815\,
            I => \ALU.a3_b_10\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \ALU.a3_b_10_cascade_\
        );

    \I__2477\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__18806\,
            I => \N__18802\
        );

    \I__2475\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18799\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__18802\,
            I => \ALU.madd_305\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__18799\,
            I => \ALU.madd_305\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__18794\,
            I => \ALU.madd_5_cascade_\
        );

    \I__2471\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18785\
        );

    \I__2470\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18785\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__18785\,
            I => \ALU.madd_19\
        );

    \I__2468\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18775\
        );

    \I__2467\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18775\
        );

    \I__2466\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18772\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__18775\,
            I => \ALU.madd_17\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__18772\,
            I => \ALU.madd_17\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__18767\,
            I => \ALU.madd_19_cascade_\
        );

    \I__2462\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__18761\,
            I => \ALU.madd_47\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__2459\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__2456\ : Span4Mux_s1_h
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__18743\,
            I => \ALU.g0_0_a3_0\
        );

    \I__2454\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18735\
        );

    \I__2453\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18732\
        );

    \I__2452\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18724\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__18735\,
            I => \N__18721\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__18732\,
            I => \N__18718\
        );

    \I__2449\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18713\
        );

    \I__2448\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18710\
        );

    \I__2447\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18703\
        );

    \I__2446\ : InMux
    port map (
            O => \N__18728\,
            I => \N__18703\
        );

    \I__2445\ : InMux
    port map (
            O => \N__18727\,
            I => \N__18703\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__18724\,
            I => \N__18698\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__18721\,
            I => \N__18698\
        );

    \I__2442\ : Span4Mux_h
    port map (
            O => \N__18718\,
            I => \N__18695\
        );

    \I__2441\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18690\
        );

    \I__2440\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18690\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18685\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__18710\,
            I => \N__18685\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__18703\,
            I => \ALU.operand2_8\
        );

    \I__2436\ : Odrv4
    port map (
            O => \N__18698\,
            I => \ALU.operand2_8\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__18695\,
            I => \ALU.operand2_8\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__18690\,
            I => \ALU.operand2_8\
        );

    \I__2433\ : Odrv12
    port map (
            O => \N__18685\,
            I => \ALU.operand2_8\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__18674\,
            I => \N__18670\
        );

    \I__2431\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18665\
        );

    \I__2430\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18662\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__18669\,
            I => \N__18659\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__18668\,
            I => \N__18656\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__18665\,
            I => \N__18652\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__18662\,
            I => \N__18649\
        );

    \I__2425\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18644\
        );

    \I__2424\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18641\
        );

    \I__2423\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18637\
        );

    \I__2422\ : Span4Mux_h
    port map (
            O => \N__18652\,
            I => \N__18632\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__18649\,
            I => \N__18632\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__18648\,
            I => \N__18629\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__18647\,
            I => \N__18624\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18619\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18619\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__18640\,
            I => \N__18615\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18609\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__18632\,
            I => \N__18609\
        );

    \I__2413\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18600\
        );

    \I__2412\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18600\
        );

    \I__2411\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18600\
        );

    \I__2410\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18600\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__18619\,
            I => \N__18597\
        );

    \I__2408\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18592\
        );

    \I__2407\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18592\
        );

    \I__2406\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18589\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__18609\,
            I => \N__18586\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__18600\,
            I => \ALU.N_199_0\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__18597\,
            I => \ALU.N_199_0\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__18592\,
            I => \ALU.N_199_0\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__18589\,
            I => \ALU.N_199_0\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__18586\,
            I => \ALU.N_199_0\
        );

    \I__2399\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__18572\,
            I => \ALU.a3_b_8\
        );

    \I__2397\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__18560\,
            I => \ALU.madd_275\
        );

    \I__2393\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__2391\ : Span4Mux_s3_h
    port map (
            O => \N__18551\,
            I => \N__18546\
        );

    \I__2390\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18541\
        );

    \I__2389\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18541\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__18546\,
            I => \N__18538\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__18541\,
            I => \N__18535\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__18538\,
            I => \ALU.madd_217\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__18535\,
            I => \ALU.madd_217\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__2383\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18522\
        );

    \I__2382\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18519\
        );

    \I__2381\ : InMux
    port map (
            O => \N__18525\,
            I => \N__18516\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__18522\,
            I => \N__18512\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__18519\,
            I => \N__18509\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18506\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__18515\,
            I => \N__18503\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__18512\,
            I => \N__18497\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__18509\,
            I => \N__18497\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__18506\,
            I => \N__18494\
        );

    \I__2373\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18489\
        );

    \I__2372\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18489\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__18497\,
            I => \ALU.madd_222\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__18494\,
            I => \ALU.madd_222\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__18489\,
            I => \ALU.madd_222\
        );

    \I__2368\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18476\
        );

    \I__2367\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18476\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__18476\,
            I => \N__18471\
        );

    \I__2365\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18466\
        );

    \I__2364\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18466\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__18471\,
            I => \N__18463\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__18466\,
            I => \ALU.madd_212\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__18463\,
            I => \ALU.madd_212\
        );

    \I__2360\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18454\
        );

    \I__2359\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__18454\,
            I => \N__18448\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__18451\,
            I => \ALU.madd_284\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__18448\,
            I => \ALU.madd_284\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__18443\,
            I => \ALU.madd_279_cascade_\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__2353\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__2351\ : Span4Mux_s3_h
    port map (
            O => \N__18431\,
            I => \N__18427\
        );

    \I__2350\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__18427\,
            I => \ALU.madd_349\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__18424\,
            I => \ALU.madd_349\
        );

    \I__2347\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18415\
        );

    \I__2346\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18412\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__18415\,
            I => \ALU.d_RNIV96U8Z0Z_13\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__18412\,
            I => \ALU.d_RNIV96U8Z0Z_13\
        );

    \I__2343\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__18398\,
            I => \N__18394\
        );

    \I__2339\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18391\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__18394\,
            I => \ALU.madd_310_0\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__18391\,
            I => \ALU.madd_310_0\
        );

    \I__2336\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__18383\,
            I => \ALU.madd_330_0\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__18380\,
            I => \ALU.c_RNIF549Z0Z_10_cascade_\
        );

    \I__2333\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__18374\,
            I => \ALU.a_RNIBLBOZ0Z_10\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \ALU.operand2_7_ns_1_10_cascade_\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__18368\,
            I => \ALU.un9_addsub_axb_12_cascade_\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \ALU.d_RNIV96U8Z0Z_13_cascade_\
        );

    \I__2328\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__18359\,
            I => \N__18355\
        );

    \I__2326\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18352\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__18355\,
            I => \ALU.madd_314\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__18352\,
            I => \ALU.madd_314\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__18347\,
            I => \ALU.madd_310_0_cascade_\
        );

    \I__2322\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18338\
        );

    \I__2321\ : InMux
    port map (
            O => \N__18343\,
            I => \N__18338\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__18338\,
            I => \ALU.madd_334\
        );

    \I__2319\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__18332\,
            I => \ALU.a1_b_12\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \ALU.a2_b_9_cascade_\
        );

    \I__2316\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__18323\,
            I => \ALU.a9_b_4\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__18320\,
            I => \ALU.a10_b_3_cascade_\
        );

    \I__2313\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18311\
        );

    \I__2312\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18311\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__18311\,
            I => \ALU.madd_319\
        );

    \I__2310\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__18302\,
            I => \ALU.madd_366\
        );

    \I__2307\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__18296\,
            I => \ALU.madd_484_11\
        );

    \I__2305\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__18287\,
            I => \ALU.madd_376\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__18284\,
            I => \ALU.madd_484_17_cascade_\
        );

    \I__2301\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__18278\,
            I => \ALU.madd_484_15\
        );

    \I__2299\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__18272\,
            I => \ALU.madd_484_20\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__2296\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18262\
        );

    \I__2295\ : InMux
    port map (
            O => \N__18265\,
            I => \N__18259\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__18262\,
            I => \N__18256\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__18259\,
            I => \N__18253\
        );

    \I__2292\ : Span4Mux_h
    port map (
            O => \N__18256\,
            I => \N__18250\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__18253\,
            I => \ALU.madd_309\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__18250\,
            I => \ALU.madd_309\
        );

    \I__2289\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18238\
        );

    \I__2287\ : InMux
    port map (
            O => \N__18241\,
            I => \N__18235\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__18238\,
            I => \N__18232\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__18235\,
            I => \N__18229\
        );

    \I__2284\ : Span4Mux_s3_h
    port map (
            O => \N__18232\,
            I => \N__18226\
        );

    \I__2283\ : Odrv12
    port map (
            O => \N__18229\,
            I => \ALU.madd_362\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__18226\,
            I => \ALU.madd_362\
        );

    \I__2281\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__18218\,
            I => \ALU.madd_391\
        );

    \I__2279\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__18206\,
            I => \ALU.a5_b_9\
        );

    \I__2275\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__2273\ : Span4Mux_h
    port map (
            O => \N__18197\,
            I => \N__18193\
        );

    \I__2272\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18190\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__18193\,
            I => \ALU.a6_b_8\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__18190\,
            I => \ALU.a6_b_8\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__18185\,
            I => \ALU.a7_b_7_cascade_\
        );

    \I__2268\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__18179\,
            I => \ALU.madd_381\
        );

    \I__2266\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__18173\,
            I => \ALU.madd_484_16\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__18170\,
            I => \ALU.dout_6_ns_1_12_cascade_\
        );

    \I__2263\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__18164\,
            I => \ALU.N_711\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__18161\,
            I => \ALU.N_759_cascade_\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__18158\,
            I => \ALU.aluOut_12_cascade_\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__2258\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18146\
        );

    \I__2257\ : InMux
    port map (
            O => \N__18151\,
            I => \N__18146\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__18146\,
            I => \ALU.a12_b_2\
        );

    \I__2255\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18127\
        );

    \I__2254\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18127\
        );

    \I__2253\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18127\
        );

    \I__2252\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18127\
        );

    \I__2251\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18127\
        );

    \I__2250\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18124\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__18127\,
            I => \N__18117\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__18124\,
            I => \N__18114\
        );

    \I__2247\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18105\
        );

    \I__2246\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18105\
        );

    \I__2245\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18105\
        );

    \I__2244\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18105\
        );

    \I__2243\ : Span4Mux_h
    port map (
            O => \N__18117\,
            I => \N__18101\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__18114\,
            I => \N__18098\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__18105\,
            I => \N__18095\
        );

    \I__2240\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18092\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__18101\,
            I => \N__18087\
        );

    \I__2238\ : Sp12to4
    port map (
            O => \N__18098\,
            I => \N__18084\
        );

    \I__2237\ : Span12Mux_h
    port map (
            O => \N__18095\,
            I => \N__18079\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18079\
        );

    \I__2235\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18074\
        );

    \I__2234\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18074\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__18087\,
            I => \ALU.N_90_0\
        );

    \I__2232\ : Odrv12
    port map (
            O => \N__18084\,
            I => \ALU.N_90_0\
        );

    \I__2231\ : Odrv12
    port map (
            O => \N__18079\,
            I => \ALU.N_90_0\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__18074\,
            I => \ALU.N_90_0\
        );

    \I__2229\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__18062\,
            I => \N__18058\
        );

    \I__2227\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18055\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__18058\,
            I => \N__18049\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__18055\,
            I => \N__18046\
        );

    \I__2224\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18039\
        );

    \I__2223\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18039\
        );

    \I__2222\ : InMux
    port map (
            O => \N__18052\,
            I => \N__18039\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__18049\,
            I => \N__18034\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__18046\,
            I => \N__18034\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__18039\,
            I => \ctrlOut_3\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__18034\,
            I => \ctrlOut_3\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__18029\,
            I => \ALU.N_235_0_cascade_\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__18026\,
            I => \ALU.a12_b_3_cascade_\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__18023\,
            I => \N__18019\
        );

    \I__2214\ : InMux
    port map (
            O => \N__18022\,
            I => \N__18014\
        );

    \I__2213\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18014\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__18014\,
            I => \ctrlOut_4\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__18011\,
            I => \ALU.a_15_m2_ns_1Z0Z_14_cascade_\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__18008\,
            I => \ALU.lshift_15_ns_1_14_cascade_\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__18005\,
            I => \ALU.lshift_14_cascade_\
        );

    \I__2208\ : InMux
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__17999\,
            I => \ALU.a_15_m2_14\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__17996\,
            I => \ALU.a_15_m4_14_cascade_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__17987\,
            I => \ALU.a_15_m3_14\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__17984\,
            I => \ALU.dout_3_ns_1_12_cascade_\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__17981\,
            I => \ALU.rshift_3_ns_1_6_cascade_\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__17978\,
            I => \ALU.N_474_cascade_\
        );

    \I__2199\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17972\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__17972\,
            I => \ALU.rshift_15_ns_1_6\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__17969\,
            I => \ALU.rshift_6_cascade_\
        );

    \I__2196\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17963\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__17960\,
            I => \ALU.N_291_0\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__17957\,
            I => \ALU.dout_6_ns_1_14_cascade_\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__17954\,
            I => \ALU.aluOut_15_cascade_\
        );

    \I__2191\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17948\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__17948\,
            I => \ALU.N_761\
        );

    \I__2189\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__17942\,
            I => \ALU.N_713\
        );

    \I__2187\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17930\
        );

    \I__2186\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17930\
        );

    \I__2185\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17930\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__17930\,
            I => \ALU.a_cnv_0Z0Z_0\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__17927\,
            I => \N__17918\
        );

    \I__2182\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17914\
        );

    \I__2181\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17911\
        );

    \I__2180\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17908\
        );

    \I__2179\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17897\
        );

    \I__2178\ : InMux
    port map (
            O => \N__17922\,
            I => \N__17897\
        );

    \I__2177\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17897\
        );

    \I__2176\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17897\
        );

    \I__2175\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17897\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__17914\,
            I => \aluResults_1\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__17911\,
            I => \aluResults_1\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__17908\,
            I => \aluResults_1\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__17897\,
            I => \aluResults_1\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__2169\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17879\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__17884\,
            I => \N__17876\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__17883\,
            I => \N__17873\
        );

    \I__2166\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17870\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__17879\,
            I => \N__17867\
        );

    \I__2164\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17862\
        );

    \I__2163\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17862\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__17870\,
            I => \ALU.b_cnv_0Z0Z_0\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__17867\,
            I => \ALU.b_cnv_0Z0Z_0\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__17862\,
            I => \ALU.b_cnv_0Z0Z_0\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__17855\,
            I => \N__17849\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__17854\,
            I => \N__17844\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__17853\,
            I => \N__17841\
        );

    \I__2156\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17836\
        );

    \I__2155\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17823\
        );

    \I__2154\ : InMux
    port map (
            O => \N__17848\,
            I => \N__17823\
        );

    \I__2153\ : InMux
    port map (
            O => \N__17847\,
            I => \N__17823\
        );

    \I__2152\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17823\
        );

    \I__2151\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17823\
        );

    \I__2150\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17823\
        );

    \I__2149\ : InMux
    port map (
            O => \N__17839\,
            I => \N__17820\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__17836\,
            I => \aluResults_2\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__17823\,
            I => \aluResults_2\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__17820\,
            I => \aluResults_2\
        );

    \I__2145\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17808\
        );

    \I__2144\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17803\
        );

    \I__2143\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17803\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17799\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__17803\,
            I => \N__17796\
        );

    \I__2140\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17793\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__17799\,
            I => \ALU.N_169_0\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__17796\,
            I => \ALU.N_169_0\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__17793\,
            I => \ALU.N_169_0\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__17786\,
            I => \ALU.c_RNIEP354Z0Z_14_cascade_\
        );

    \I__2135\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17780\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__17780\,
            I => \ALU.c_RNIJENJ8_0Z0Z_15\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__17777\,
            I => \testClock_0_cascade_\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__17774\,
            I => \ALU.a_cnv_0Z0Z_0_cascade_\
        );

    \I__2131\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__17768\,
            I => \ALU.N_53_0\
        );

    \I__2129\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17759\
        );

    \I__2128\ : InMux
    port map (
            O => \N__17764\,
            I => \N__17759\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__17756\,
            I => \aluResults_0\
        );

    \I__2125\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__17750\,
            I => \testClock_0\
        );

    \I__2123\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17740\
        );

    \I__2122\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17731\
        );

    \I__2121\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17731\
        );

    \I__2120\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17731\
        );

    \I__2119\ : InMux
    port map (
            O => \N__17743\,
            I => \N__17731\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__17740\,
            I => \testClockZ0\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__17731\,
            I => \testClockZ0\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__17726\,
            I => \ALU.madd_41_cascade_\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__17723\,
            I => \ALU.madd_46_cascade_\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__17720\,
            I => \ALU.madd_39_cascade_\
        );

    \I__2113\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17711\
        );

    \I__2112\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17711\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__17708\,
            I => \ALU.a6_b_3\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__17705\,
            I => \ALU.madd_78_0_tz_cascade_\
        );

    \I__2108\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__17699\,
            I => \ALU.madd_78_0\
        );

    \I__2106\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__17693\,
            I => \ALU.madd_39\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__17690\,
            I => \ALU.madd_78_0_cascade_\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__17687\,
            I => \ALU.madd_114_cascade_\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__17684\,
            I => \ALU.g1_2_cascade_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__17678\,
            I => \ALU.a4_b_0_7\
        );

    \I__2099\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17672\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__17669\,
            I => \ALU.g2_0_0_0\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__17666\,
            I => \ALU.un2_addsub_axb_5_cascade_\
        );

    \I__2095\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__17654\,
            I => \ALU.a6_b_0_7\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__17651\,
            I => \ALU.a6_b_0_cascade_\
        );

    \I__2090\ : InMux
    port map (
            O => \N__17648\,
            I => \N__17642\
        );

    \I__2089\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17642\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__17642\,
            I => \ALU.madd_275_0\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__17639\,
            I => \ALU.madd_42_cascade_\
        );

    \I__2086\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__17633\,
            I => \ALU.madd_42_0\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__17630\,
            I => \ALU.e_RNIM09HZ0Z_7_cascade_\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__17627\,
            I => \ALU.operand2_7_ns_1_7_cascade_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__17618\,
            I => \N__17615\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__17615\,
            I => \ALU.a2_b_6\
        );

    \I__2078\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__17609\,
            I => \N__17606\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__17603\,
            I => \ALU.a0_b_8\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__17600\,
            I => \ALU.a2_b_6_cascade_\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__17597\,
            I => \ALU.a5_b_6_cascade_\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__17594\,
            I => \ALU.operand2_5_cascade_\
        );

    \I__2071\ : InMux
    port map (
            O => \N__17591\,
            I => \N__17585\
        );

    \I__2070\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17585\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__17585\,
            I => \N__17582\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__17579\,
            I => \ALU.madd_176_0\
        );

    \I__2066\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17570\
        );

    \I__2065\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17570\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__17567\,
            I => \N__17563\
        );

    \I__2062\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17560\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__17563\,
            I => \ALU.madd_218_0\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__17560\,
            I => \ALU.madd_218_0\
        );

    \I__2059\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17551\
        );

    \I__2058\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17548\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__17551\,
            I => \ALU.a7_b_4\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__17548\,
            I => \ALU.a7_b_4\
        );

    \I__2055\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__2053\ : Span4Mux_s1_h
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__17534\,
            I => \N__17529\
        );

    \I__2051\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17526\
        );

    \I__2050\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17523\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__17529\,
            I => \ALU.a6_b_5\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__17526\,
            I => \ALU.a6_b_5\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__17523\,
            I => \ALU.a6_b_5\
        );

    \I__2046\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__2044\ : Span4Mux_s2_h
    port map (
            O => \N__17510\,
            I => \N__17506\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__17509\,
            I => \N__17503\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__17506\,
            I => \N__17500\
        );

    \I__2041\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17497\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__17500\,
            I => \ALU.a5_b_6\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__17497\,
            I => \ALU.a5_b_6\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__17492\,
            I => \N__17487\
        );

    \I__2037\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17484\
        );

    \I__2036\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17481\
        );

    \I__2035\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17478\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__17484\,
            I => \N__17475\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__17481\,
            I => \N__17472\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__17478\,
            I => \N__17469\
        );

    \I__2031\ : Span12Mux_s2_h
    port map (
            O => \N__17475\,
            I => \N__17466\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__17472\,
            I => \N__17461\
        );

    \I__2029\ : Span4Mux_s2_h
    port map (
            O => \N__17469\,
            I => \N__17461\
        );

    \I__2028\ : Odrv12
    port map (
            O => \N__17466\,
            I => \ALU.madd_320\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__17461\,
            I => \ALU.madd_320\
        );

    \I__2026\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17451\
        );

    \I__2025\ : InMux
    port map (
            O => \N__17455\,
            I => \N__17448\
        );

    \I__2024\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17445\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__17451\,
            I => \ALU.madd_325_0\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__17448\,
            I => \ALU.madd_325_0\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__17445\,
            I => \ALU.madd_325_0\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \ALU.madd_274_cascade_\
        );

    \I__2019\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17428\
        );

    \I__2017\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17425\
        );

    \I__2016\ : Span4Mux_v
    port map (
            O => \N__17428\,
            I => \N__17422\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__17425\,
            I => \N__17419\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__17422\,
            I => \ALU.madd_254\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__17419\,
            I => \ALU.madd_254\
        );

    \I__2012\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__2010\ : Span4Mux_s2_h
    port map (
            O => \N__17408\,
            I => \N__17404\
        );

    \I__2009\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17401\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__17404\,
            I => \ALU.madd_344\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__17401\,
            I => \ALU.madd_344\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__17396\,
            I => \ALU.madd_29_cascade_\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__17393\,
            I => \ALU.madd_47_cascade_\
        );

    \I__2004\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__17384\,
            I => \ALU.madd_265_0\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__17381\,
            I => \N__17377\
        );

    \I__2000\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17374\
        );

    \I__1999\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17371\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__17374\,
            I => \N__17368\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__1996\ : Span12Mux_h
    port map (
            O => \N__17368\,
            I => \N__17362\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__17362\,
            I => \ALU.madd_260\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__17359\,
            I => \ALU.madd_260\
        );

    \I__1992\ : InMux
    port map (
            O => \N__17354\,
            I => \N__17348\
        );

    \I__1991\ : InMux
    port map (
            O => \N__17353\,
            I => \N__17348\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__17348\,
            I => \ALU.madd_329\
        );

    \I__1989\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17339\
        );

    \I__1988\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17339\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__17339\,
            I => \ALU.madd_407\
        );

    \I__1986\ : InMux
    port map (
            O => \N__17336\,
            I => \N__17333\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__17333\,
            I => \ALU.madd_412\
        );

    \I__1984\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__17327\,
            I => \ALU.madd_i3_mux_1\
        );

    \I__1982\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__17321\,
            I => \ALU.madd_330\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__1979\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17312\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__17312\,
            I => \N__17309\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__17309\,
            I => \N__17306\
        );

    \I__1976\ : Span4Mux_s0_h
    port map (
            O => \N__17306\,
            I => \N__17303\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__17303\,
            I => \ALU.madd_141_1\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__17300\,
            I => \N__17296\
        );

    \I__1973\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17291\
        );

    \I__1972\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17284\
        );

    \I__1971\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17284\
        );

    \I__1970\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17284\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__17291\,
            I => \ALU.madd_270_0\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__17284\,
            I => \ALU.madd_270_0\
        );

    \I__1967\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__17276\,
            I => \ALU.madd_250_0\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__17273\,
            I => \ALU.madd_250_0_cascade_\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__1963\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__1960\ : Span4Mux_s0_h
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__17255\,
            I => \ALU.madd_250\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__17252\,
            I => \N__17247\
        );

    \I__1957\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17244\
        );

    \I__1956\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17239\
        );

    \I__1955\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17239\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__17244\,
            I => \N__17236\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__17239\,
            I => \N__17233\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__17236\,
            I => \ALU.a3_b_9\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__17233\,
            I => \ALU.a3_b_9\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \ALU.madd_250_cascade_\
        );

    \I__1949\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17221\
        );

    \I__1948\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17218\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__17221\,
            I => \N__17215\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__17218\,
            I => \N__17208\
        );

    \I__1945\ : Span4Mux_s2_h
    port map (
            O => \N__17215\,
            I => \N__17205\
        );

    \I__1944\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17198\
        );

    \I__1943\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17198\
        );

    \I__1942\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17198\
        );

    \I__1941\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17195\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__17208\,
            I => \ALU.madd_207\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__17205\,
            I => \ALU.madd_207\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__17198\,
            I => \ALU.madd_207\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__17195\,
            I => \ALU.madd_207\
        );

    \I__1936\ : InMux
    port map (
            O => \N__17186\,
            I => \N__17180\
        );

    \I__1935\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17180\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__17180\,
            I => \ALU.madd_274\
        );

    \I__1933\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__17174\,
            I => \ALU.madd_372_0\
        );

    \I__1931\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17165\
        );

    \I__1930\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17165\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__17165\,
            I => \ALU.madd_382\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__17162\,
            I => \ALU.madd_377_cascade_\
        );

    \I__1927\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17156\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__17156\,
            I => \N__17152\
        );

    \I__1925\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__17152\,
            I => \ALU.a13_b_1\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__17149\,
            I => \ALU.a13_b_1\
        );

    \I__1922\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__17141\,
            I => \ALU.madd_397\
        );

    \I__1920\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17132\
        );

    \I__1919\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17132\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__17132\,
            I => \ALU.madd_392\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__17129\,
            I => \ALU.madd_397_cascade_\
        );

    \I__1916\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17120\
        );

    \I__1915\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17120\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__17117\,
            I => \ALU.madd_339\
        );

    \I__1912\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__17111\,
            I => \ALU.madd_406\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__17108\,
            I => \ALU.a5_b_8_cascade_\
        );

    \I__1909\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17102\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__17102\,
            I => \ALU.madd_387\
        );

    \I__1907\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17093\
        );

    \I__1906\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17093\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__17093\,
            I => \ALU.madd_329_0\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__17090\,
            I => \ALU.madd_387_cascade_\
        );

    \I__1903\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17084\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__17084\,
            I => \ALU.madd_402\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__17081\,
            I => \ALU.madd_402_cascade_\
        );

    \I__1900\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__17075\,
            I => \ALU.madd_354\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__17072\,
            I => \ALU.madd_412_cascade_\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__17069\,
            I => \ALU.madd_324_0_cascade_\
        );

    \I__1896\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__17063\,
            I => \N__17060\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__17060\,
            I => \ALU.madd_372\
        );

    \I__1893\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__17054\,
            I => \ALU.madd_396\
        );

    \I__1891\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__17048\,
            I => \ALU.madd_484_21\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__17045\,
            I => \ALU.madd_411_cascade_\
        );

    \I__1888\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__17039\,
            I => \ALU.madd_484_24\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__1885\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17027\
        );

    \I__1884\ : InMux
    port map (
            O => \N__17032\,
            I => \N__17027\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__17027\,
            I => \ALU.a8_b_6\
        );

    \I__1882\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17018\
        );

    \I__1881\ : InMux
    port map (
            O => \N__17023\,
            I => \N__17018\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__17018\,
            I => \ALU.a9_b_5\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__1878\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__17009\,
            I => \ALU.madd_377\
        );

    \I__1876\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__17003\,
            I => \ALU.a11_b_3\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \ALU.a11_b_3_cascade_\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__16997\,
            I => \N__16993\
        );

    \I__1872\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16988\
        );

    \I__1871\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16988\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__16988\,
            I => \ctrlOut_14\
        );

    \I__1869\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__16982\,
            I => \N__16977\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16972\
        );

    \I__1866\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16972\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__16977\,
            I => \N__16967\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__16972\,
            I => \N__16967\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__16967\,
            I => \N__16963\
        );

    \I__1862\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16960\
        );

    \I__1861\ : Span4Mux_s0_h
    port map (
            O => \N__16963\,
            I => \N__16957\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__16960\,
            I => \RXbuffer_6\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__16957\,
            I => \RXbuffer_6\
        );

    \I__1858\ : InMux
    port map (
            O => \N__16952\,
            I => \N__16949\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__16949\,
            I => \N__16945\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__16948\,
            I => \N__16942\
        );

    \I__1855\ : Span4Mux_s2_v
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__1854\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__16939\,
            I => \testWordZ0Z_14\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__16936\,
            I => \testWordZ0Z_14\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__16931\,
            I => \ALU.a7_b_6_cascade_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16922\
        );

    \I__1849\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16922\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__16922\,
            I => \ALU.a6_b_7\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__1846\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__16913\,
            I => \ALU.a7_b_6\
        );

    \I__1844\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__16907\,
            I => \ALU.madd_324_0\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__16904\,
            I => \ALU.a13_b_1_cascade_\
        );

    \I__1841\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__16898\,
            I => \ALU.un2_addsub_axb_14\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__16895\,
            I => \ALU.un2_addsub_axb_9_cascade_\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__16892\,
            I => \N_662_0_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__16886\,
            I => \N_665_0\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__16883\,
            I => \N_301_0_cascade_\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \N_668_0_cascade_\
        );

    \I__1833\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__16874\,
            I => \ALU.m300_nsZ0Z_1\
        );

    \I__1831\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16868\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__16865\,
            I => \N__16860\
        );

    \I__1828\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16855\
        );

    \I__1827\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16855\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__16860\,
            I => \N_662_0\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__16855\,
            I => \N_662_0\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \N_670_0_cascade_\
        );

    \I__1823\ : CEMux
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__16844\,
            I => \N__16840\
        );

    \I__1821\ : CEMux
    port map (
            O => \N__16843\,
            I => \N__16837\
        );

    \I__1820\ : Span4Mux_s2_v
    port map (
            O => \N__16840\,
            I => \N__16834\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__16837\,
            I => \N__16831\
        );

    \I__1818\ : Sp12to4
    port map (
            O => \N__16834\,
            I => \N__16828\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__16831\,
            I => \N__16825\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__16828\,
            I => \CONTROL.results_cnvZ0Z_0\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__16825\,
            I => \CONTROL.results_cnvZ0Z_0\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__16820\,
            I => \N_51_0_cascade_\
        );

    \I__1813\ : InMux
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__1811\ : IoSpan4Mux
    port map (
            O => \N__16811\,
            I => \N__16807\
        );

    \I__1810\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16804\
        );

    \I__1809\ : IoSpan4Mux
    port map (
            O => \N__16807\,
            I => \N__16799\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__16804\,
            I => \N__16799\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__16799\,
            I => \testWordZ0Z_15\
        );

    \I__1806\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__16793\,
            I => \N__16789\
        );

    \I__1804\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16786\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__16789\,
            I => \ALU.madd_129\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__16786\,
            I => \ALU.madd_129\
        );

    \I__1801\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__16778\,
            I => \ALU.a5_b_4\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__16775\,
            I => \ALU.a5_b_4_cascade_\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \ALU.madd_133_cascade_\
        );

    \I__1797\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16763\
        );

    \I__1796\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16763\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__16760\,
            I => \N__16756\
        );

    \I__1793\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16753\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__16756\,
            I => \N__16750\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__16753\,
            I => \N__16747\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__16750\,
            I => \ALU.madd_237_0_tz_0\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__16747\,
            I => \ALU.madd_237_0_tz_0\
        );

    \I__1788\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16736\
        );

    \I__1787\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16736\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__16736\,
            I => \ALU.madd_133\
        );

    \I__1785\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16729\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16722\
        );

    \I__1782\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16717\
        );

    \I__1781\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16717\
        );

    \I__1780\ : Sp12to4
    port map (
            O => \N__16722\,
            I => \N__16712\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16712\
        );

    \I__1778\ : Span12Mux_v
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__16709\,
            I => \ALU.madd_138\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__16706\,
            I => \ALU.madd_128_0_0_0_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16694\
        );

    \I__1774\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16694\
        );

    \I__1773\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16694\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__16694\,
            I => \ALU.madd_70\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__16691\,
            I => \ALU.madd_237_0_tz_0_1_cascade_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16682\
        );

    \I__1769\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16679\
        );

    \I__1768\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16674\
        );

    \I__1767\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16674\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__16682\,
            I => \N__16669\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__16679\,
            I => \N__16669\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__16674\,
            I => \N__16666\
        );

    \I__1763\ : Span12Mux_v
    port map (
            O => \N__16669\,
            I => \N__16663\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__16666\,
            I => \ALU.g0_0_0\
        );

    \I__1761\ : Odrv12
    port map (
            O => \N__16663\,
            I => \ALU.g0_0_0\
        );

    \I__1760\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__1758\ : Sp12to4
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__1757\ : Odrv12
    port map (
            O => \N__16649\,
            I => \ALU.N_1537_0_0_1\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__16646\,
            I => \ALU.i6_mux_cascade_\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \ALU.un2_addsub_axb_7_cascade_\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__16640\,
            I => \ALU.a0_b_8_cascade_\
        );

    \I__1753\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16633\
        );

    \I__1752\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16630\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__16633\,
            I => \ALU.madd_103\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__16630\,
            I => \ALU.madd_103\
        );

    \I__1749\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__16622\,
            I => \ALU.madd_124\
        );

    \I__1747\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16610\
        );

    \I__1746\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16610\
        );

    \I__1745\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16610\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__16610\,
            I => \ALU.madd_148\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__16607\,
            I => \ALU.madd_148_cascade_\
        );

    \I__1742\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16598\
        );

    \I__1741\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16598\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__16598\,
            I => \ALU.madd_247_0_tz_0\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__1738\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16587\
        );

    \I__1737\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16584\
        );

    \I__1736\ : InMux
    port map (
            O => \N__16590\,
            I => \N__16581\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__16587\,
            I => \ALU.madd_143\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__16584\,
            I => \ALU.madd_143\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__16581\,
            I => \ALU.madd_143\
        );

    \I__1732\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16567\
        );

    \I__1731\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16567\
        );

    \I__1730\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16564\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__16567\,
            I => \ALU.madd_181\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__16564\,
            I => \ALU.madd_181\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__16559\,
            I => \ALU.madd_280_cascade_\
        );

    \I__1726\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16550\
        );

    \I__1725\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16550\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__16547\,
            I => \ALU.madd_285\
        );

    \I__1722\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16541\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__16541\,
            I => \ALU.madd_326\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__16538\,
            I => \N__16534\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__16537\,
            I => \N__16531\
        );

    \I__1718\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16526\
        );

    \I__1717\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16526\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__16520\,
            I => \ALU.a4_b_7\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__16517\,
            I => \ALU.a4_b_7_cascade_\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__16514\,
            I => \ALU.madd_233_cascade_\
        );

    \I__1711\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16507\
        );

    \I__1710\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16504\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__16507\,
            I => \N__16499\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__16504\,
            I => \N__16499\
        );

    \I__1707\ : Odrv12
    port map (
            O => \N__16499\,
            I => \ALU.madd_237\
        );

    \I__1706\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16492\
        );

    \I__1705\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16489\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__16492\,
            I => \ALU.madd_242\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__16489\,
            I => \ALU.madd_242\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__16484\,
            I => \ALU.madd_247_cascade_\
        );

    \I__1701\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__16478\,
            I => \ALU.madd_295_0\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__1698\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__16469\,
            I => \ALU.madd_N_10\
        );

    \I__1696\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__16463\,
            I => \ALU.madd_247\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__16460\,
            I => \ALU.madd_N_10_cascade_\
        );

    \I__1693\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__16454\,
            I => \ALU.madd_N_5_0\
        );

    \I__1691\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16444\
        );

    \I__1690\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16444\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__16449\,
            I => \N__16441\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__16444\,
            I => \N__16438\
        );

    \I__1687\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16435\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__16438\,
            I => \ALU.madd_190\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__16435\,
            I => \ALU.madd_190\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__16430\,
            I => \N__16427\
        );

    \I__1683\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16421\
        );

    \I__1682\ : InMux
    port map (
            O => \N__16426\,
            I => \N__16421\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__16421\,
            I => \N__16418\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__16418\,
            I => \ALU.madd_238_0\
        );

    \I__1679\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__16412\,
            I => \ALU.madd_233\
        );

    \I__1677\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16404\
        );

    \I__1676\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16399\
        );

    \I__1675\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16399\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__16404\,
            I => \ALU.madd_327\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__16399\,
            I => \ALU.madd_327\
        );

    \I__1672\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16388\
        );

    \I__1671\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16388\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__16388\,
            I => \ALU.madd_208\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__16385\,
            I => \ALU.N_225_0_cascade_\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__16382\,
            I => \ALU.madd_290_0_cascade_\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__16379\,
            I => \ALU.madd_299_cascade_\
        );

    \I__1666\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16373\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__16370\,
            I => \N__16365\
        );

    \I__1663\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16360\
        );

    \I__1662\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16360\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__16365\,
            I => \N__16357\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__16360\,
            I => \N__16354\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__16357\,
            I => \ALU.g0_11\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__16354\,
            I => \ALU.g0_11\
        );

    \I__1657\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16346\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__16346\,
            I => \N__16342\
        );

    \I__1655\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16339\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__16342\,
            I => \ALU.madd_299\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__16339\,
            I => \ALU.madd_299\
        );

    \I__1652\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__16328\,
            I => \ALU.madd_223_0\
        );

    \I__1649\ : InMux
    port map (
            O => \N__16325\,
            I => \N__16321\
        );

    \I__1648\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16318\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__16321\,
            I => \ALU.madd_228\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__16318\,
            I => \ALU.madd_228\
        );

    \I__1645\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16309\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__16312\,
            I => \N__16304\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__16309\,
            I => \N__16301\
        );

    \I__1642\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16296\
        );

    \I__1641\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16296\
        );

    \I__1640\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16293\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__16301\,
            I => \ALU.madd_170\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__16296\,
            I => \ALU.madd_170\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__16293\,
            I => \ALU.madd_170\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__16286\,
            I => \ALU.madd_265_0_cascade_\
        );

    \I__1635\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16280\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16275\
        );

    \I__1633\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16272\
        );

    \I__1632\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16269\
        );

    \I__1631\ : Odrv12
    port map (
            O => \N__16275\,
            I => \ALU.madd_280\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__16272\,
            I => \ALU.madd_280\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__16269\,
            I => \ALU.madd_280\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__16262\,
            I => \ALU.madd_223_0_cascade_\
        );

    \I__1627\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16256\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__16256\,
            I => \ALU.N_1533_0\
        );

    \I__1625\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__16250\,
            I => \N__16247\
        );

    \I__1623\ : Span4Mux_s2_h
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__16244\,
            I => \ALU.N_1559_0\
        );

    \I__1621\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16235\
        );

    \I__1620\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16235\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__16235\,
            I => \ALU.madd_165_0_tz\
        );

    \I__1618\ : InMux
    port map (
            O => \N__16232\,
            I => \N__16228\
        );

    \I__1617\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16225\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__16228\,
            I => \ALU.madd_165_0\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__16225\,
            I => \ALU.madd_165_0\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__1613\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16214\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__16214\,
            I => \ALU.a5_b_5\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__16211\,
            I => \ALU.a5_b_5_cascade_\
        );

    \I__1610\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16204\
        );

    \I__1609\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16201\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__16204\,
            I => \N__16196\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__16201\,
            I => \N__16196\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__16196\,
            I => \ALU.a4_b_6\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__16193\,
            I => \ALU.madd_175_cascade_\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__16190\,
            I => \N__16186\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__16189\,
            I => \N__16182\
        );

    \I__1602\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16178\
        );

    \I__1601\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16171\
        );

    \I__1600\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16171\
        );

    \I__1599\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16171\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__16178\,
            I => \N__16166\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__16171\,
            I => \N__16166\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__16166\,
            I => \ALU.madd_232\
        );

    \I__1595\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16160\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__16160\,
            I => \ALU.madd_175\
        );

    \I__1593\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16151\
        );

    \I__1592\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16151\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__16151\,
            I => \ALU.madd_213_0\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \ALU.a7_b_4_cascade_\
        );

    \I__1589\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16142\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__16142\,
            I => \ALU.madd_i1_mux_2\
        );

    \I__1587\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16135\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__16138\,
            I => \N__16132\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__16135\,
            I => \N__16129\
        );

    \I__1584\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16126\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__16129\,
            I => \ALU.madd_289\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__16126\,
            I => \ALU.madd_289\
        );

    \I__1581\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16115\
        );

    \I__1580\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16115\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__16115\,
            I => \ALU.madd_227\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__16112\,
            I => \ALU.madd_227_cascade_\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__16109\,
            I => \ALU.madd_165_0_0_cascade_\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__16106\,
            I => \ALU.madd_170_0_tz_cascade_\
        );

    \I__1575\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16098\
        );

    \I__1574\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16093\
        );

    \I__1573\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16093\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16090\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__16093\,
            I => \ALU.madd_90\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__16090\,
            I => \ALU.madd_90\
        );

    \I__1569\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__16082\,
            I => \ALU.madd_340_0\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__16079\,
            I => \ALU.g0_1_cascade_\
        );

    \I__1566\ : InMux
    port map (
            O => \N__16076\,
            I => \N__16073\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__16073\,
            I => \ALU.g2\
        );

    \I__1564\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16067\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__16067\,
            I => \ALU.N_1545_1\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__16064\,
            I => \ALU.g0_3_cascade_\
        );

    \I__1561\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__16058\,
            I => \ALU.madd_350_0\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__16055\,
            I => \ALU.madd_350_0_cascade_\
        );

    \I__1558\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16044\
        );

    \I__1557\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16044\
        );

    \I__1556\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16041\
        );

    \I__1555\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16038\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__16044\,
            I => \ALU.madd_335\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__16041\,
            I => \ALU.madd_335\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__16038\,
            I => \ALU.madd_335\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__16031\,
            I => \ALU.a4_b_8_cascade_\
        );

    \I__1550\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16022\
        );

    \I__1549\ : InMux
    port map (
            O => \N__16027\,
            I => \N__16022\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__16022\,
            I => \ALU.madd_269\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__16019\,
            I => \ALU.madd_i1_mux_cascade_\
        );

    \I__1546\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__16013\,
            I => \N__16009\
        );

    \I__1544\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16006\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__16009\,
            I => \N__16003\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__16006\,
            I => \N__16000\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__16003\,
            I => \ALU.g0_14\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__16000\,
            I => \ALU.g0_14\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__15995\,
            I => \ALU.madd_i3_mux_cascade_\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__15992\,
            I => \ALU.madd_331_cascade_\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__15989\,
            I => \N__15985\
        );

    \I__1536\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15980\
        );

    \I__1535\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15980\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__15980\,
            I => \ALU.madd_328\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__15977\,
            I => \ALU.N_275_0_cascade_\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__15971\,
            I => \ALU.g0_0_0_N_3L3\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__15968\,
            I => \ALU.g0_0_0_N_4L5_cascade_\
        );

    \I__1529\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__15962\,
            I => \ALU.g0_0_0_N_3L3_0\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__15959\,
            I => \ALU.a5_b_9_cascade_\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__15956\,
            I => \ALU.operand2_8_cascade_\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__15953\,
            I => \N__15950\
        );

    \I__1524\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__15941\,
            I => \N__15938\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__15938\,
            I => \ALU.a1_b_8\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__15935\,
            I => \ALU.a1_b_8_cascade_\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__15932\,
            I => \N_661_0_cascade_\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \ALU.un2_addsub_axb_8_cascade_\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__15926\,
            I => \N__15922\
        );

    \I__1515\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15916\
        );

    \I__1514\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15916\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__15921\,
            I => \N__15913\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__15916\,
            I => \N__15910\
        );

    \I__1511\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__15910\,
            I => \RXbuffer_0\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__15907\,
            I => \RXbuffer_0\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__15902\,
            I => \N__15898\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__15901\,
            I => \N__15893\
        );

    \I__1506\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15887\
        );

    \I__1505\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15887\
        );

    \I__1504\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15884\
        );

    \I__1503\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15881\
        );

    \I__1502\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15878\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__15887\,
            I => \N__15875\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15870\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__15881\,
            I => \N__15870\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__15878\,
            I => \RXbuffer_7\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__15875\,
            I => \RXbuffer_7\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__15870\,
            I => \RXbuffer_7\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__15863\,
            I => \N__15858\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__15862\,
            I => \N__15854\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__15861\,
            I => \N__15851\
        );

    \I__1492\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15847\
        );

    \I__1491\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15842\
        );

    \I__1490\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15842\
        );

    \I__1489\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15839\
        );

    \I__1488\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15836\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__15847\,
            I => \N__15833\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__15842\,
            I => \N__15830\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__15839\,
            I => \N__15827\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__15836\,
            I => \RXbuffer_1\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__15833\,
            I => \RXbuffer_1\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__15830\,
            I => \RXbuffer_1\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__15827\,
            I => \RXbuffer_1\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__15818\,
            I => \N__15815\
        );

    \I__1479\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15806\
        );

    \I__1478\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15806\
        );

    \I__1477\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15803\
        );

    \I__1476\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15798\
        );

    \I__1475\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15798\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__15806\,
            I => \N__15795\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__15803\,
            I => \N__15788\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__15798\,
            I => \N__15788\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__15795\,
            I => \N__15788\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__15788\,
            I => \N__15785\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__15785\,
            I => \RXbuffer_3\
        );

    \I__1468\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__1466\ : Span4Mux_s0_v
    port map (
            O => \N__15776\,
            I => \N__15772\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__15775\,
            I => \N__15769\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__15772\,
            I => \N__15766\
        );

    \I__1463\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15763\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__15766\,
            I => \testWordZ0Z_13\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__15763\,
            I => \testWordZ0Z_13\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__15758\,
            I => \ALU.m304_nsZ0Z_1_cascade_\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__15755\,
            I => \ALU.i73_mux_1_cascade_\
        );

    \I__1458\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15749\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__15749\,
            I => \clkdivZ0Z_16\
        );

    \I__1456\ : InMux
    port map (
            O => \N__15746\,
            I => \bfn_1_18_0_\
        );

    \I__1455\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__15740\,
            I => \clkdivZ0Z_17\
        );

    \I__1453\ : InMux
    port map (
            O => \N__15737\,
            I => clkdiv_cry_16
        );

    \I__1452\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15731\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__15731\,
            I => \clkdivZ0Z_18\
        );

    \I__1450\ : InMux
    port map (
            O => \N__15728\,
            I => clkdiv_cry_17
        );

    \I__1449\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15722\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__15722\,
            I => \clkdivZ0Z_19\
        );

    \I__1447\ : InMux
    port map (
            O => \N__15719\,
            I => clkdiv_cry_18
        );

    \I__1446\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15713\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__15713\,
            I => \clkdivZ0Z_20\
        );

    \I__1444\ : InMux
    port map (
            O => \N__15710\,
            I => clkdiv_cry_19
        );

    \I__1443\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__15704\,
            I => \clkdivZ0Z_21\
        );

    \I__1441\ : InMux
    port map (
            O => \N__15701\,
            I => clkdiv_cry_20
        );

    \I__1440\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__15695\,
            I => \clkdivZ0Z_22\
        );

    \I__1438\ : InMux
    port map (
            O => \N__15692\,
            I => clkdiv_cry_21
        );

    \I__1437\ : InMux
    port map (
            O => \N__15689\,
            I => clkdiv_cry_22
        );

    \I__1436\ : IoInMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__1434\ : Span12Mux_s7_v
    port map (
            O => \N__15680\,
            I => \N__15676\
        );

    \I__1433\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__1432\ : Odrv12
    port map (
            O => \N__15676\,
            I => \GPIO3_c\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__15673\,
            I => \GPIO3_c\
        );

    \I__1430\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__15665\,
            I => \clkdivZ0Z_7\
        );

    \I__1428\ : InMux
    port map (
            O => \N__15662\,
            I => clkdiv_cry_6
        );

    \I__1427\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__15656\,
            I => \clkdivZ0Z_8\
        );

    \I__1425\ : InMux
    port map (
            O => \N__15653\,
            I => \bfn_1_17_0_\
        );

    \I__1424\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15647\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__15647\,
            I => \clkdivZ0Z_9\
        );

    \I__1422\ : InMux
    port map (
            O => \N__15644\,
            I => clkdiv_cry_8
        );

    \I__1421\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__15638\,
            I => \clkdivZ0Z_10\
        );

    \I__1419\ : InMux
    port map (
            O => \N__15635\,
            I => clkdiv_cry_9
        );

    \I__1418\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__15629\,
            I => \clkdivZ0Z_11\
        );

    \I__1416\ : InMux
    port map (
            O => \N__15626\,
            I => clkdiv_cry_10
        );

    \I__1415\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__15620\,
            I => \clkdivZ0Z_12\
        );

    \I__1413\ : InMux
    port map (
            O => \N__15617\,
            I => clkdiv_cry_11
        );

    \I__1412\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15611\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__15611\,
            I => \clkdivZ0Z_13\
        );

    \I__1410\ : InMux
    port map (
            O => \N__15608\,
            I => clkdiv_cry_12
        );

    \I__1409\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15602\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__15602\,
            I => \clkdivZ0Z_14\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15599\,
            I => clkdiv_cry_13
        );

    \I__1406\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15593\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__15593\,
            I => \clkdivZ0Z_15\
        );

    \I__1404\ : InMux
    port map (
            O => \N__15590\,
            I => clkdiv_cry_14
        );

    \I__1403\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15583\
        );

    \I__1402\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15580\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__15583\,
            I => \ALU.madd_324\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__15580\,
            I => \ALU.madd_324\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__15575\,
            I => \ALU.madd_326_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15567\
        );

    \I__1397\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15562\
        );

    \I__1396\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15562\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__15567\,
            I => \ALU.madd_325\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__15562\,
            I => \ALU.madd_325\
        );

    \I__1393\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__15554\,
            I => \clkdivZ0Z_0\
        );

    \I__1391\ : InMux
    port map (
            O => \N__15551\,
            I => \bfn_1_16_0_\
        );

    \I__1390\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__15545\,
            I => \clkdivZ0Z_1\
        );

    \I__1388\ : InMux
    port map (
            O => \N__15542\,
            I => clkdiv_cry_0
        );

    \I__1387\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15536\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__15536\,
            I => \clkdivZ0Z_2\
        );

    \I__1385\ : InMux
    port map (
            O => \N__15533\,
            I => clkdiv_cry_1
        );

    \I__1384\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15527\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__15527\,
            I => \clkdivZ0Z_3\
        );

    \I__1382\ : InMux
    port map (
            O => \N__15524\,
            I => clkdiv_cry_2
        );

    \I__1381\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__15518\,
            I => \clkdivZ0Z_4\
        );

    \I__1379\ : InMux
    port map (
            O => \N__15515\,
            I => clkdiv_cry_3
        );

    \I__1378\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15509\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__15509\,
            I => \clkdivZ0Z_5\
        );

    \I__1376\ : InMux
    port map (
            O => \N__15506\,
            I => clkdiv_cry_4
        );

    \I__1375\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__15500\,
            I => \clkdivZ0Z_6\
        );

    \I__1373\ : InMux
    port map (
            O => \N__15497\,
            I => clkdiv_cry_5
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__15494\,
            I => \ALU.madd_144_cascade_\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__15491\,
            I => \ALU.madd_324_cascade_\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__15488\,
            I => \ALU.madd_N_9_cascade_\
        );

    \I__1369\ : InMux
    port map (
            O => \N__15485\,
            I => \N__15482\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__15482\,
            I => \ALU.madd_191_0\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__15479\,
            I => \N__15473\
        );

    \I__1366\ : InMux
    port map (
            O => \N__15478\,
            I => \N__15468\
        );

    \I__1365\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15468\
        );

    \I__1364\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15463\
        );

    \I__1363\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15463\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__15468\,
            I => \N__15460\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__15463\,
            I => \N__15455\
        );

    \I__1360\ : Span4Mux_s1_h
    port map (
            O => \N__15460\,
            I => \N__15455\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__15455\,
            I => \ALU.madd_186\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__15452\,
            I => \ALU.madd_191_0_cascade_\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__15449\,
            I => \ALU.a8_b_3_cascade_\
        );

    \I__1356\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15441\
        );

    \I__1355\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15438\
        );

    \I__1354\ : InMux
    port map (
            O => \N__15444\,
            I => \N__15435\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__15441\,
            I => \ALU.a8_b_3\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__15438\,
            I => \ALU.a8_b_3\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__15435\,
            I => \ALU.a8_b_3\
        );

    \I__1350\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__15422\,
            I => \ALU.g0_0_2\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__15419\,
            I => \ALU.g0_0_cascade_\
        );

    \I__1346\ : InMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__15413\,
            I => \ALU.N_1527_1_0\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__15410\,
            I => \N__15407\
        );

    \I__1343\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15404\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__15404\,
            I => \N__15401\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__15401\,
            I => \N__15398\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__15398\,
            I => \ALU.g2_0_1\
        );

    \I__1339\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__15392\,
            I => \ALU.g1\
        );

    \I__1337\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15386\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__15383\,
            I => \ALU.g0_1_0\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__15380\,
            I => \ALU.madd_124_0_cascade_\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__15377\,
            I => \ALU.madd_124_cascade_\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \ALU.madd_171_cascade_\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__15371\,
            I => \ALU.madd_161_0_cascade_\
        );

    \I__1330\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__15365\,
            I => \ALU.madd_161\
        );

    \I__1328\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15356\
        );

    \I__1327\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15356\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__15353\,
            I => \ALU.madd_166\
        );

    \I__1324\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15347\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__15347\,
            I => \ALU.madd_171\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__15344\,
            I => \ALU.madd_161_cascade_\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \ALU.N_217_0_cascade_\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \ALU.un9_addsub_axb_10_cascade_\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__15335\,
            I => \ALU.a3_b_0_10_cascade_\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__15332\,
            I => \ALU.g0_2_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__15326\,
            I => \ALU.N_1555_0\
        );

    \I__1315\ : InMux
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__15320\,
            I => \ALU.N_1527_0\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__15317\,
            I => \ALU.madd_254_0_tz_cascade_\
        );

    \I__1312\ : InMux
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__15311\,
            I => \ALU.madd_141\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__15308\,
            I => \ALU.madd_254_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15301\
        );

    \I__1308\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15298\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__15301\,
            I => \ALU.madd_254_0_tz\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__15298\,
            I => \ALU.madd_254_0_tz\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__15293\,
            I => \N__15290\
        );

    \I__1304\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__15287\,
            I => \ALU.m292_nsZ0Z_1\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__15284\,
            I => \ALU.N_90_0_cascade_\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__15281\,
            I => \N__15277\
        );

    \I__1300\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15272\
        );

    \I__1299\ : InMux
    port map (
            O => \N__15277\,
            I => \N__15272\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__15272\,
            I => \ctrlOut_6\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__15269\,
            I => \ALU.madd_315_0_cascade_\
        );

    \I__1296\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15263\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__15263\,
            I => \ALU.a12_b_1\
        );

    \I__1294\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15257\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__15257\,
            I => \ALU.madd_315_0\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__15254\,
            I => \ALU.a12_b_1_cascade_\
        );

    \I__1291\ : InMux
    port map (
            O => \N__15251\,
            I => \N__15245\
        );

    \I__1290\ : InMux
    port map (
            O => \N__15250\,
            I => \N__15245\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__15245\,
            I => \ALU.madd_264\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__15242\,
            I => \ALU.madd_141_0_cascade_\
        );

    \I__1287\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__15236\,
            I => \ALU.N_1545_0\
        );

    \I__1285\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__15230\,
            I => \ALU.madd_166_0\
        );

    \I__1283\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15215\
        );

    \I__1282\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15215\
        );

    \I__1281\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15215\
        );

    \I__1280\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15215\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__15215\,
            I => \ctrlOut_5\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__15212\,
            I => \ALU.N_223_0_cascade_\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \ALU.a9_b_3_cascade_\
        );

    \I__1276\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15200\
        );

    \I__1275\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15200\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__15200\,
            I => \ALU.a7_b_5\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__15197\,
            I => \N__15194\
        );

    \I__1272\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15191\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__15191\,
            I => \ALU.a9_b_3\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__15188\,
            I => \ALU.g0_0_a3_2_0_cascade_\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__15185\,
            I => \N__15181\
        );

    \I__1268\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15176\
        );

    \I__1267\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15176\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__15176\,
            I => \ctrlOut_8\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \ALU.m289_nsZ0Z_1_cascade_\
        );

    \INVFTDI.TXshift_1C\ : INV
    port map (
            O => \INVFTDI.TXshift_1C_net\,
            I => \N__47602\
        );

    \INVFTDI.TXshift_0C\ : INV
    port map (
            O => \INVFTDI.TXshift_0C_net\,
            I => \N__47607\
        );

    \INVFTDI.baudAcc_1C\ : INV
    port map (
            O => \INVFTDI.baudAcc_1C_net\,
            I => \N__47604\
        );

    \INVFTDI.TXstate_0C\ : INV
    port map (
            O => \INVFTDI.TXstate_0C_net\,
            I => \N__47601\
        );

    \INVFTDI.gap_2C\ : INV
    port map (
            O => \INVFTDI.gap_2C_net\,
            I => \N__47599\
        );

    \INVFTDI.baudAcc_0C\ : INV
    port map (
            O => \INVFTDI.baudAcc_0C_net\,
            I => \N__47603\
        );

    \INVFTDI.gap_0C\ : INV
    port map (
            O => \INVFTDI.gap_0C_net\,
            I => \N__47609\
        );

    \INVFTDI.RXreadyC\ : INV
    port map (
            O => \INVFTDI.RXreadyC_net\,
            I => \N__47617\
        );

    \INVFTDI.RXbuffer_0C\ : INV
    port map (
            O => \INVFTDI.RXbuffer_0C_net\,
            I => \N__47667\
        );

    \INVFTDI.RXbuffer_3C\ : INV
    port map (
            O => \INVFTDI.RXbuffer_3C_net\,
            I => \N__47654\
        );

    \IN_MUX_bfv_13_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_2_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.madd_cry_7\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_7,
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_15,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.un9_addsub_cry_7\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.un2_addsub_cry_7\,
            carryinitout => \bfn_6_10_0_\
        );

    \testState_RNIB7C_0_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__30743\,
            GLOBALBUFFEROUTPUT => \testState_i_g_2\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \FTDI.RXbuffer_3_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32266\,
            lcout => \RXbuffer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_3C_net\,
            ce => \N__20510\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_4_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25538\,
            lcout => \RXbuffer_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_3C_net\,
            ce => \N__20510\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_0_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15850\,
            lcout => \RXbuffer_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_0C_net\,
            ce => \N__20509\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41534\,
            lcout => \RXbuffer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_0C_net\,
            ce => \N__20509\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_2_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15813\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RXbuffer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_0C_net\,
            ce => \N__20509\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_5_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16966\,
            lcout => \RXbuffer_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_0C_net\,
            ce => \N__20509\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_6_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15892\,
            lcout => \RXbuffer_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_0C_net\,
            ce => \N__20509\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_7_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RXbuffer_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_0C_net\,
            ce => \N__20509\,
            sr => \_gnd_net_\
        );

    \ALU.f_8_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48261\,
            in1 => \N__47893\,
            in2 => \_gnd_net_\,
            in3 => \N__47808\,
            lcout => \ALU.fZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47674\,
            ce => \N__36363\,
            sr => \_gnd_net_\
        );

    \ALU.m198_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110111011"
        )
    port map (
            in0 => \N__30200\,
            in1 => \N__29739\,
            in2 => \N__15185\,
            in3 => \N__25206\,
            lcout => \ALU.N_199_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_24_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__41486\,
            in1 => \N__41201\,
            in2 => \N__15926\,
            in3 => \N__15184\,
            lcout => \ctrlOut_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_8_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__41204\,
            in1 => \N__26844\,
            in2 => \N__41508\,
            in3 => \N__15925\,
            lcout => \testWordZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_25_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__41487\,
            in1 => \N__41202\,
            in2 => \N__15862\,
            in3 => \N__19747\,
            lcout => \ctrlOut_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_9_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__41205\,
            in1 => \N__27155\,
            in2 => \N__41509\,
            in3 => \N__15857\,
            lcout => \testWordZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_13_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__25534\,
            in1 => \N__41490\,
            in2 => \N__15775\,
            in3 => \N__41199\,
            lcout => \testWordZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_15_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__41200\,
            in1 => \N__16810\,
            in2 => \N__41507\,
            in3 => \N__15897\,
            lcout => \testWordZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_31_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__41488\,
            in1 => \N__41203\,
            in2 => \N__15902\,
            in3 => \N__20940\,
            lcout => \ctrlOut_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47677\,
            ce => \N__41054\,
            sr => \_gnd_net_\
        );

    \testWord_21_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15227\,
            in1 => \N__41489\,
            in2 => \N__25545\,
            in3 => \N__18104\,
            lcout => \ctrlOut_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47683\,
            ce => \N__41053\,
            sr => \_gnd_net_\
        );

    \ALU.m289_ns_1_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000010000"
        )
    port map (
            in0 => \N__30206\,
            in1 => \N__26568\,
            in2 => \N__29756\,
            in3 => \N__15225\,
            lcout => OPEN,
            ltout => \ALU.m289_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1K464_5_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__15226\,
            in1 => \N__29436\,
            in2 => \N__15173\,
            in3 => \N__40390\,
            lcout => \ALU.N_290_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m222_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011111101111"
        )
    port map (
            in0 => \N__30205\,
            in1 => \N__25216\,
            in2 => \N__29755\,
            in3 => \N__15224\,
            lcout => \ALU.N_223_0\,
            ltout => \ALU.N_223_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVULB7_5_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__24311\,
            in1 => \N__46942\,
            in2 => \N__15212\,
            in3 => \N__21728\,
            lcout => \ALU.a7_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINF4M7_3_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23916\,
            in1 => \N__39849\,
            in2 => \N__24242\,
            in3 => \N__24044\,
            lcout => \ALU.a9_b_3\,
            ltout => \ALU.a9_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_260_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__42687\,
            in1 => \N__40102\,
            in2 => \N__15209\,
            in3 => \N__15206\,
            lcout => \ALU.madd_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_264_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__15205\,
            in1 => \N__40103\,
            in2 => \N__15197\,
            in3 => \N__42688\,
            lcout => \ALU.madd_264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_166_0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010011010"
        )
    port map (
            in0 => \N__46715\,
            in1 => \N__41737\,
            in2 => \N__46973\,
            in3 => \N__42690\,
            lcout => \ALU.madd_166_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_a3_2_0_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__42692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46956\,
            lcout => OPEN,
            ltout => \ALU.g0_0_a3_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g2_0_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001101010"
        )
    port map (
            in0 => \N__18526\,
            in1 => \N__17516\,
            in2 => \N__15188\,
            in3 => \N__17543\,
            lcout => \ALU.g2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_2_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17454\,
            in1 => \N__15239\,
            in2 => \N__17492\,
            in3 => \N__16049\,
            lcout => \ALU.g0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_315_0_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011010010"
        )
    port map (
            in0 => \N__27598\,
            in1 => \N__41738\,
            in2 => \N__39854\,
            in3 => \N__42691\,
            lcout => \ALU.madd_315_0\,
            ltout => \ALU.madd_315_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_335_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16027\,
            in1 => \N__15250\,
            in2 => \N__15269\,
            in3 => \N__15266\,
            lcout => \ALU.madd_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI8LNC7_12_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25355\,
            in2 => \_gnd_net_\,
            in3 => \N__37773\,
            lcout => \ALU.a12_b_1\,
            ltout => \ALU.a12_b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_339_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__16028\,
            in1 => \N__15260\,
            in2 => \N__15254\,
            in3 => \N__15251\,
            lcout => \ALU.madd_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_5_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38315\,
            in1 => \N__25353\,
            in2 => \N__39608\,
            in3 => \N__36984\,
            lcout => OPEN,
            ltout => \ALU.madd_141_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_4_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__37235\,
            in1 => \N__27600\,
            in2 => \N__15242\,
            in3 => \N__15304\,
            lcout => \ALU.N_1545_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_166_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__15233\,
            in1 => \N__39850\,
            in2 => \_gnd_net_\,
            in3 => \N__37757\,
            lcout => \ALU.madd_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_252_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36983\,
            in1 => \N__39600\,
            in2 => \N__25371\,
            in3 => \N__38311\,
            lcout => \ALU.madd_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_254_0_tz_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__39601\,
            in1 => \N__25352\,
            in2 => \N__38336\,
            in3 => \N__36982\,
            lcout => \ALU.madd_254_0_tz\,
            ltout => \ALU.madd_254_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_254_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__37234\,
            in1 => \N__27599\,
            in2 => \N__15317\,
            in3 => \N__15314\,
            lcout => \ALU.madd_254\,
            ltout => \ALU.madd_254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_340_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17491\,
            in2 => \N__15308\,
            in3 => \N__17455\,
            lcout => \ALU.madd_340_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__15305\,
            in1 => \N__27601\,
            in2 => \N__17318\,
            in3 => \N__37236\,
            lcout => \ALU.N_1545_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFD4D4_3_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101110111"
        )
    port map (
            in0 => \N__18053\,
            in1 => \N__29404\,
            in2 => \N__15293\,
            in3 => \N__42012\,
            lcout => \ALU.N_293_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_3_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__18091\,
            in1 => \N__22203\,
            in2 => \N__15818\,
            in3 => \N__41506\,
            lcout => \testWordZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47688\,
            ce => \N__41052\,
            sr => \_gnd_net_\
        );

    \testWord_19_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__18054\,
            in1 => \N__15814\,
            in2 => \N__41510\,
            in3 => \N__18090\,
            lcout => \ctrlOut_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47688\,
            ce => \N__41052\,
            sr => \_gnd_net_\
        );

    \ALU.m292_ns_1_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001010"
        )
    port map (
            in0 => \N__29729\,
            in1 => \N__18052\,
            in2 => \N__26588\,
            in3 => \N__30195\,
            lcout => \ALU.m292_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m89_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__21902\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30323\,
            lcout => \ALU.N_90_0\,
            ltout => \ALU.N_90_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_22_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__41502\,
            in2 => \N__15284\,
            in3 => \N__15280\,
            lcout => \ctrlOut_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47688\,
            ce => \N__41052\,
            sr => \_gnd_net_\
        );

    \ALU.m216_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001111111"
        )
    port map (
            in0 => \N__30194\,
            in1 => \N__25225\,
            in2 => \N__15281\,
            in3 => \N__29728\,
            lcout => \ALU.N_217_0\,
            ltout => \ALU.N_217_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIT7NA7_6_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__29980\,
            in1 => \N__42958\,
            in2 => \N__15341\,
            in3 => \N__26727\,
            lcout => \ALU.a4_b_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1DA1A_10_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111100010"
        )
    port map (
            in0 => \N__20023\,
            in1 => \N__26498\,
            in2 => \N__20065\,
            in3 => \N__27602\,
            lcout => OPEN,
            ltout => \ALU.un9_addsub_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIV2S0F_10_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15338\,
            in3 => \N__39571\,
            lcout => \ALU.a_RNIV2S0FZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILMFN5_10_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__20024\,
            in1 => \_gnd_net_\,
            in2 => \N__20066\,
            in3 => \N__26497\,
            lcout => \ALU.N_192_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVRI59_10_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__26499\,
            in1 => \N__41994\,
            in2 => \N__20108\,
            in3 => \N__20022\,
            lcout => OPEN,
            ltout => \ALU.a3_b_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_15_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28274\,
            in1 => \N__15389\,
            in2 => \N__15335\,
            in3 => \N__18407\,
            lcout => OPEN,
            ltout => \ALU.g0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_14_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18458\,
            in1 => \N__15329\,
            in2 => \N__15332\,
            in3 => \N__19688\,
            lcout => \ALU.g0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_16_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__15323\,
            in1 => \_gnd_net_\,
            in2 => \N__18530\,
            in3 => \N__18557\,
            lcout => \ALU.N_1555_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_17_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__39471\,
            in1 => \N__15445\,
            in2 => \N__18758\,
            in3 => \N__37937\,
            lcout => \ALU.N_1527_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_165_0_tz_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__37934\,
            in1 => \N__39595\,
            in2 => \N__27586\,
            in3 => \N__38308\,
            lcout => \ALU.madd_165_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_163_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38309\,
            in1 => \N__27534\,
            in2 => \N__39607\,
            in3 => \N__37935\,
            lcout => \ALU.madd_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_171_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110111010010"
        )
    port map (
            in0 => \N__41955\,
            in1 => \N__47089\,
            in2 => \N__16220\,
            in3 => \N__16208\,
            lcout => \ALU.madd_171\,
            ltout => \ALU.madd_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_190_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__17590\,
            in1 => \N__15368\,
            in2 => \N__15374\,
            in3 => \N__15361\,
            lcout => \ALU.madd_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_161_0_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__37936\,
            in1 => \N__39599\,
            in2 => \N__40112\,
            in3 => \N__37195\,
            lcout => OPEN,
            ltout => \ALU.madd_161_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_161_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__38310\,
            in1 => \_gnd_net_\,
            in2 => \N__15371\,
            in3 => \N__27535\,
            lcout => \ALU.madd_161\,
            ltout => \ALU.madd_161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_186_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15362\,
            in1 => \N__15350\,
            in2 => \N__15344\,
            in3 => \N__17591\,
            lcout => \ALU.madd_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_208_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__27595\,
            in1 => \N__15444\,
            in2 => \N__37758\,
            in3 => \N__21234\,
            lcout => \ALU.madd_208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIF74M7_3_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23944\,
            in1 => \N__40093\,
            in2 => \N__24312\,
            in3 => \N__24022\,
            lcout => \ALU.a8_b_3\,
            ltout => \ALU.a8_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_212_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__27596\,
            in1 => \N__21235\,
            in2 => \N__15449\,
            in3 => \N__37731\,
            lcout => \ALU.madd_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_24_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__37732\,
            in1 => \N__27597\,
            in2 => \N__21239\,
            in3 => \N__15446\,
            lcout => \ALU.N_1527_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_22_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001101100"
        )
    port map (
            in0 => \N__17251\,
            in1 => \N__15428\,
            in2 => \N__17270\,
            in3 => \N__17225\,
            lcout => OPEN,
            ltout => \ALU.g0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_11_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16253\,
            in1 => \N__16012\,
            in2 => \N__15419\,
            in3 => \N__15395\,
            lcout => \ALU.g0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__15416\,
            in1 => \N__16279\,
            in2 => \N__15410\,
            in3 => \N__16658\,
            lcout => \ALU.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_13_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__39397\,
            in1 => \N__37199\,
            in2 => \N__40772\,
            in3 => \N__38317\,
            lcout => \ALU.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_10_ma_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15586\,
            lcout => \ALU.madd_cry_10_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_124_0_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__39814\,
            in1 => \N__46918\,
            in2 => \N__37233\,
            in3 => \N__38316\,
            lcout => OPEN,
            ltout => \ALU.madd_124_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_124_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__37742\,
            in1 => \N__40094\,
            in2 => \N__15380\,
            in3 => \_gnd_net_\,
            lcout => \ALU.madd_124\,
            ltout => \ALU.madd_124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_144_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16637\,
            in2 => \N__15377\,
            in3 => \N__16796\,
            lcout => \ALU.madd_144\,
            ltout => \ALU.madd_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_158_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20354\,
            in2 => \N__15494\,
            in3 => \N__19355\,
            lcout => \ALU.madd_324\,
            ltout => \ALU.madd_324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_9_l_ofx_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__19295\,
            in1 => \N__15570\,
            in2 => \N__15491\,
            in3 => \N__19277\,
            lcout => \ALU.madd_axb_9_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_134_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__23749\,
            in1 => \N__36994\,
            in2 => \N__15953\,
            in3 => \N__47051\,
            lcout => \ALU.madd_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_196_0_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15477\,
            in1 => \N__16574\,
            in2 => \N__16595\,
            in3 => \N__16617\,
            lcout => OPEN,
            ltout => \ALU.madd_N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m4_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__15476\,
            in1 => \N__20318\,
            in2 => \N__15488\,
            in3 => \N__16407\,
            lcout => \ALU.madd_N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_127_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46911\,
            in1 => \N__37194\,
            in2 => \N__40120\,
            in3 => \N__37741\,
            lcout => \ALU.madd_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_196_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16618\,
            in1 => \N__20524\,
            in2 => \N__15479\,
            in3 => \N__15485\,
            lcout => \ALU.madd_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_191_0_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16573\,
            in2 => \_gnd_net_\,
            in3 => \N__16591\,
            lcout => \ALU.madd_191_0\,
            ltout => \ALU.madd_191_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_200_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__16619\,
            in1 => \N__15478\,
            in2 => \N__15452\,
            in3 => \N__20525\,
            lcout => \ALU.madd_326\,
            ltout => \ALU.madd_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_10_l_ofx_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__16408\,
            in1 => \N__15587\,
            in2 => \N__15575\,
            in3 => \N__15572\,
            lcout => \ALU.madd_axb_10_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_0_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15557\,
            in2 => \_gnd_net_\,
            in3 => \N__15551\,
            lcout => \clkdivZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => clkdiv_cry_0,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_1_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15548\,
            in2 => \_gnd_net_\,
            in3 => \N__15542\,
            lcout => \clkdivZ0Z_1\,
            ltout => OPEN,
            carryin => clkdiv_cry_0,
            carryout => clkdiv_cry_1,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_2_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15539\,
            in2 => \_gnd_net_\,
            in3 => \N__15533\,
            lcout => \clkdivZ0Z_2\,
            ltout => OPEN,
            carryin => clkdiv_cry_1,
            carryout => clkdiv_cry_2,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_3_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15530\,
            in2 => \_gnd_net_\,
            in3 => \N__15524\,
            lcout => \clkdivZ0Z_3\,
            ltout => OPEN,
            carryin => clkdiv_cry_2,
            carryout => clkdiv_cry_3,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_4_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15521\,
            in2 => \_gnd_net_\,
            in3 => \N__15515\,
            lcout => \clkdivZ0Z_4\,
            ltout => OPEN,
            carryin => clkdiv_cry_3,
            carryout => clkdiv_cry_4,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_5_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15512\,
            in2 => \_gnd_net_\,
            in3 => \N__15506\,
            lcout => \clkdivZ0Z_5\,
            ltout => OPEN,
            carryin => clkdiv_cry_4,
            carryout => clkdiv_cry_5,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_6_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15503\,
            in2 => \_gnd_net_\,
            in3 => \N__15497\,
            lcout => \clkdivZ0Z_6\,
            ltout => OPEN,
            carryin => clkdiv_cry_5,
            carryout => clkdiv_cry_6,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_7_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15668\,
            in2 => \_gnd_net_\,
            in3 => \N__15662\,
            lcout => \clkdivZ0Z_7\,
            ltout => OPEN,
            carryin => clkdiv_cry_6,
            carryout => clkdiv_cry_7,
            clk => \N__47691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_8_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15659\,
            in2 => \_gnd_net_\,
            in3 => \N__15653\,
            lcout => \clkdivZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => clkdiv_cry_8,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_9_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15650\,
            in2 => \_gnd_net_\,
            in3 => \N__15644\,
            lcout => \clkdivZ0Z_9\,
            ltout => OPEN,
            carryin => clkdiv_cry_8,
            carryout => clkdiv_cry_9,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_10_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15641\,
            in2 => \_gnd_net_\,
            in3 => \N__15635\,
            lcout => \clkdivZ0Z_10\,
            ltout => OPEN,
            carryin => clkdiv_cry_9,
            carryout => clkdiv_cry_10,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_11_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15632\,
            in2 => \_gnd_net_\,
            in3 => \N__15626\,
            lcout => \clkdivZ0Z_11\,
            ltout => OPEN,
            carryin => clkdiv_cry_10,
            carryout => clkdiv_cry_11,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_12_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15623\,
            in2 => \_gnd_net_\,
            in3 => \N__15617\,
            lcout => \clkdivZ0Z_12\,
            ltout => OPEN,
            carryin => clkdiv_cry_11,
            carryout => clkdiv_cry_12,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_13_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15614\,
            in2 => \_gnd_net_\,
            in3 => \N__15608\,
            lcout => \clkdivZ0Z_13\,
            ltout => OPEN,
            carryin => clkdiv_cry_12,
            carryout => clkdiv_cry_13,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_14_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15605\,
            in2 => \_gnd_net_\,
            in3 => \N__15599\,
            lcout => \clkdivZ0Z_14\,
            ltout => OPEN,
            carryin => clkdiv_cry_13,
            carryout => clkdiv_cry_14,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_15_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15596\,
            in2 => \_gnd_net_\,
            in3 => \N__15590\,
            lcout => \clkdivZ0Z_15\,
            ltout => OPEN,
            carryin => clkdiv_cry_14,
            carryout => clkdiv_cry_15,
            clk => \N__47692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_16_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15752\,
            in2 => \_gnd_net_\,
            in3 => \N__15746\,
            lcout => \clkdivZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => clkdiv_cry_16,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_17_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15743\,
            in2 => \_gnd_net_\,
            in3 => \N__15737\,
            lcout => \clkdivZ0Z_17\,
            ltout => OPEN,
            carryin => clkdiv_cry_16,
            carryout => clkdiv_cry_17,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_18_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15734\,
            in2 => \_gnd_net_\,
            in3 => \N__15728\,
            lcout => \clkdivZ0Z_18\,
            ltout => OPEN,
            carryin => clkdiv_cry_17,
            carryout => clkdiv_cry_18,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_19_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15725\,
            in2 => \_gnd_net_\,
            in3 => \N__15719\,
            lcout => \clkdivZ0Z_19\,
            ltout => OPEN,
            carryin => clkdiv_cry_18,
            carryout => clkdiv_cry_19,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_20_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15716\,
            in2 => \_gnd_net_\,
            in3 => \N__15710\,
            lcout => \clkdivZ0Z_20\,
            ltout => OPEN,
            carryin => clkdiv_cry_19,
            carryout => clkdiv_cry_20,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_21_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15707\,
            in2 => \_gnd_net_\,
            in3 => \N__15701\,
            lcout => \clkdivZ0Z_21\,
            ltout => OPEN,
            carryin => clkdiv_cry_20,
            carryout => clkdiv_cry_21,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_22_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15698\,
            in2 => \_gnd_net_\,
            in3 => \N__15692\,
            lcout => \clkdivZ0Z_22\,
            ltout => OPEN,
            carryin => clkdiv_cry_21,
            carryout => clkdiv_cry_22,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_23_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15679\,
            in2 => \_gnd_net_\,
            in3 => \N__15689\,
            lcout => \GPIO3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.results_e_0_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15782\,
            lcout => \aluResults_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47642\,
            ce => \N__16847\,
            sr => \_gnd_net_\
        );

    \testWord_18_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__20277\,
            in1 => \N__41431\,
            in2 => \N__41544\,
            in3 => \N__18120\,
            lcout => \ctrlOut_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47648\,
            ce => \N__41059\,
            sr => \_gnd_net_\
        );

    \ALU.m304_ns_1_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111110101"
        )
    port map (
            in0 => \N__22402\,
            in1 => \N__22687\,
            in2 => \N__33300\,
            in3 => \N__20276\,
            lcout => OPEN,
            ltout => \ALU.m304_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m304_ns_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011011110111"
        )
    port map (
            in0 => \N__33261\,
            in1 => \N__22280\,
            in2 => \N__15758\,
            in3 => \N__38733\,
            lcout => \N_305_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_2_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__18122\,
            in1 => \N__41538\,
            in2 => \N__41475\,
            in3 => \N__22409\,
            lcout => \testWordZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47648\,
            ce => \N__41059\,
            sr => \_gnd_net_\
        );

    \testWord_1_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__22692\,
            in1 => \N__41430\,
            in2 => \N__15863\,
            in3 => \N__18121\,
            lcout => \testWordZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47648\,
            ce => \N__41059\,
            sr => \_gnd_net_\
        );

    \testWord_5_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__18123\,
            in1 => \N__25546\,
            in2 => \N__41476\,
            in3 => \N__33263\,
            lcout => \testWordZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47648\,
            ce => \N__41059\,
            sr => \_gnd_net_\
        );

    \ALU.m656_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101111100"
        )
    port map (
            in0 => \N__21568\,
            in1 => \N__33259\,
            in2 => \N__22719\,
            in3 => \N__22403\,
            lcout => OPEN,
            ltout => \ALU.i73_mux_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m657_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__22281\,
            in1 => \N__33262\,
            in2 => \N__15755\,
            in3 => \N__22691\,
            lcout => i53_mux_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_8_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48109\,
            in1 => \N__47894\,
            in2 => \_gnd_net_\,
            in3 => \N__47809\,
            lcout => \ALU.gZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47655\,
            ce => \N__36069\,
            sr => \_gnd_net_\
        );

    \testWord_16_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__41423\,
            in1 => \N__18139\,
            in2 => \N__15921\,
            in3 => \N__21564\,
            lcout => \ctrlOut_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \testWord_23_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__18141\,
            in1 => \N__41425\,
            in2 => \N__15901\,
            in3 => \N__19867\,
            lcout => \ctrlOut_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \testWord_7_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__15896\,
            in1 => \N__41429\,
            in2 => \N__27745\,
            in3 => \N__18143\,
            lcout => \testWordZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \testWord_17_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__18140\,
            in1 => \N__41424\,
            in2 => \N__15861\,
            in3 => \N__21846\,
            lcout => \ctrlOut_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \testWord_4_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__22504\,
            in1 => \N__41428\,
            in2 => \N__32291\,
            in3 => \N__18142\,
            lcout => \testWordZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \testWord_11_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__15811\,
            in1 => \N__41427\,
            in2 => \N__34545\,
            in3 => \N__41206\,
            lcout => \testWordZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \testWord_27_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__41207\,
            in1 => \N__41426\,
            in2 => \N__24892\,
            in3 => \N__15812\,
            lcout => \ctrlOut_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47661\,
            ce => \N__41058\,
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_rep2_e_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__33296\,
            in1 => \N__19576\,
            in2 => \N__19540\,
            in3 => \N__22257\,
            lcout => \aluReadBus_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47668\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_N_3L3_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__21097\,
            in1 => \N__32738\,
            in2 => \N__29898\,
            in3 => \N__37484\,
            lcout => \ALU.g0_0_0_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_e_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__33295\,
            in1 => \N__19575\,
            in2 => \N__19539\,
            in3 => \N__22256\,
            lcout => \aluReadBus\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47668\,
            ce => \N__34710\,
            sr => \_gnd_net_\
        );

    \ALU.m8_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__29837\,
            in1 => \_gnd_net_\,
            in2 => \N__30217\,
            in3 => \N__29746\,
            lcout => \ALU.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m660_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__22430\,
            in2 => \_gnd_net_\,
            in3 => \N__22255\,
            lcout => OPEN,
            ltout => \N_661_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_cnv_0_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101100000000"
        )
    port map (
            in0 => \N__16871\,
            in1 => \N__33294\,
            in2 => \N__15932\,
            in3 => \N__34668\,
            lcout => \CONTROL.aluOperation_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m9_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111011101"
        )
    port map (
            in0 => \N__29745\,
            in1 => \N__30207\,
            in2 => \_gnd_net_\,
            in3 => \N__29836\,
            lcout => \ALU.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m634_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__22431\,
            in1 => \N__22493\,
            in2 => \_gnd_net_\,
            in3 => \N__22720\,
            lcout => \ALU.N_635_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIR21R7_8_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011000101"
        )
    port map (
            in0 => \N__18728\,
            in1 => \N__18627\,
            in2 => \N__26535\,
            in3 => \N__40079\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQ74VB_8_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15929\,
            in3 => \N__21484\,
            lcout => \ALU.d_RNIQ74VBZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN2L24_8_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__18729\,
            in1 => \_gnd_net_\,
            in2 => \N__26536\,
            in3 => \N__18628\,
            lcout => \ALU.N_201_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI60794_8_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__40080\,
            in1 => \_gnd_net_\,
            in2 => \N__18648\,
            in3 => \N__29435\,
            lcout => OPEN,
            ltout => \ALU.N_275_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUSVB61_8_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000011"
        )
    port map (
            in0 => \N__44448\,
            in1 => \N__43165\,
            in2 => \N__15977\,
            in3 => \N__19385\,
            lcout => \ALU.a_15_m3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_N_4L5_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__27593\,
            in1 => \N__37244\,
            in2 => \N__40107\,
            in3 => \N__38332\,
            lcout => OPEN,
            ltout => \ALU.g0_0_0_N_4L5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010001110"
        )
    port map (
            in0 => \N__15974\,
            in1 => \N__15965\,
            in2 => \N__15968\,
            in3 => \N__21617\,
            lcout => \ALU.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_N_3L3_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000000000"
        )
    port map (
            in0 => \N__24325\,
            in1 => \N__18727\,
            in2 => \N__18647\,
            in3 => \N__36995\,
            lcout => \ALU.g0_0_0_N_3L3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRAM58_9_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__21089\,
            in1 => \N__20868\,
            in2 => \N__30023\,
            in3 => \N__40388\,
            lcout => \ALU.a5_b_9\,
            ltout => \ALU.a5_b_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_382_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100111100"
        )
    port map (
            in0 => \N__47099\,
            in1 => \N__18196\,
            in2 => \N__15959\,
            in3 => \N__46944\,
            lcout => \ALU.madd_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVPQD3_8_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32996\,
            in1 => \N__25604\,
            in2 => \_gnd_net_\,
            in3 => \N__30875\,
            lcout => \ALU.operand2_8\,
            ltout => \ALU.operand2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC54P6_8_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__24232\,
            in1 => \N__18614\,
            in2 => \N__15956\,
            in3 => \N__37447\,
            lcout => \ALU.a1_b_8\,
            ltout => \ALU.a1_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_138_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__23750\,
            in1 => \N__36996\,
            in2 => \N__15935\,
            in3 => \N__47097\,
            lcout => \ALU.madd_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGG5I7_8_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000000000"
        )
    port map (
            in0 => \N__24233\,
            in1 => \N__18716\,
            in2 => \N__18640\,
            in3 => \N__42959\,
            lcout => OPEN,
            ltout => \ALU.a4_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_269_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__23783\,
            in1 => \N__40389\,
            in2 => \N__16031\,
            in3 => \N__47098\,
            lcout => \ALU.madd_269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2AVH7_8_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__18618\,
            in1 => \N__18717\,
            in2 => \N__30024\,
            in3 => \N__46736\,
            lcout => \ALU.a6_b_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m3_1_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000110110111"
        )
    port map (
            in0 => \N__17575\,
            in1 => \N__16686\,
            in2 => \N__16537\,
            in3 => \N__16768\,
            lcout => OPEN,
            ltout => \ALU.madd_i1_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m6_0_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18569\,
            in2 => \N__16019\,
            in3 => \N__16283\,
            lcout => OPEN,
            ltout => \ALU.madd_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110110001110"
        )
    port map (
            in0 => \N__16061\,
            in1 => \N__16016\,
            in2 => \N__15995\,
            in3 => \N__16139\,
            lcout => \ALU.madd_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001101010"
        )
    port map (
            in0 => \N__17042\,
            in1 => \N__17414\,
            in2 => \N__18440\,
            in3 => \N__17087\,
            lcout => OPEN,
            ltout => \ALU.madd_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_14_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__17354\,
            in1 => \N__15988\,
            in2 => \N__15992\,
            in3 => \N__17324\,
            lcout => \ALU.madd_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_13_l_ofx_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__16349\,
            in1 => \N__16376\,
            in2 => \N__15989\,
            in3 => \N__17353\,
            lcout => \ALU.madd_axb_13_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_237_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__17576\,
            in1 => \N__16685\,
            in2 => \N__16538\,
            in3 => \N__16769\,
            lcout => \ALU.madd_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_325_0_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101010000"
        )
    port map (
            in0 => \N__22048\,
            in1 => \N__21444\,
            in2 => \N__42990\,
            in3 => \N__40432\,
            lcout => \ALU.madd_325_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_354_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011101000"
        )
    port map (
            in0 => \N__16051\,
            in1 => \N__17186\,
            in2 => \N__16138\,
            in3 => \N__16085\,
            lcout => \ALU.madd_354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g2_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__40084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28084\,
            lcout => \ALU.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_10_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011000110"
        )
    port map (
            in0 => \N__40431\,
            in1 => \N__42957\,
            in2 => \N__21469\,
            in3 => \N__22047\,
            lcout => OPEN,
            ltout => \ALU.g0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_3_2_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20201\,
            in1 => \N__17663\,
            in2 => \N__16079\,
            in3 => \N__16076\,
            lcout => OPEN,
            ltout => \ALU.g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16070\,
            in1 => \N__16050\,
            in2 => \N__16064\,
            in3 => \N__17185\,
            lcout => \ALU.madd_350_0\,
            ltout => \ALU.madd_350_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m6_2_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16145\,
            in2 => \N__16055\,
            in3 => \N__16052\,
            lcout => \ALU.madd_i3_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICJE9B_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010100101011"
        )
    port map (
            in0 => \N__40043\,
            in1 => \N__20642\,
            in2 => \N__21470\,
            in3 => \N__47308\,
            lcout => \ALU.d_RNICJE9BZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIV4344_8_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__24318\,
            in1 => \N__18655\,
            in2 => \_gnd_net_\,
            in3 => \N__18731\,
            lcout => \ALU.N_201_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m3_3_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000111010111"
        )
    port map (
            in0 => \N__16121\,
            in1 => \N__17214\,
            in2 => \N__17300\,
            in3 => \N__16185\,
            lcout => \ALU.madd_i1_mux_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_289_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__17213\,
            in1 => \N__17295\,
            in2 => \N__16189\,
            in3 => \N__16120\,
            lcout => \ALU.madd_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIJ8B8_9_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__20867\,
            in1 => \N__21096\,
            in2 => \N__26494\,
            in3 => \N__42011\,
            lcout => \ALU.a3_b_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_227_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101000"
        )
    port map (
            in0 => \N__19980\,
            in1 => \N__16103\,
            in2 => \N__16312\,
            in3 => \N__16231\,
            lcout => \ALU.madd_227\,
            ltout => \ALU.madd_227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_285_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17294\,
            in1 => \N__17212\,
            in2 => \N__16112\,
            in3 => \N__16181\,
            lcout => \ALU.madd_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_21_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__16241\,
            in1 => \_gnd_net_\,
            in2 => \N__37237\,
            in3 => \N__40086\,
            lcout => OPEN,
            ltout => \ALU.madd_165_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_18_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001000"
        )
    port map (
            in0 => \N__16102\,
            in1 => \N__19982\,
            in2 => \N__16109\,
            in3 => \N__16307\,
            lcout => \ALU.N_1533_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_170_0_tz_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__39807\,
            in1 => \N__46686\,
            in2 => \N__37767\,
            in3 => \N__42662\,
            lcout => OPEN,
            ltout => \ALU.madd_170_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_170_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__46963\,
            in1 => \N__41726\,
            in2 => \N__16106\,
            in3 => \N__23390\,
            lcout => \ALU.madd_170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_223_0_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__19981\,
            in1 => \N__16101\,
            in2 => \_gnd_net_\,
            in3 => \N__16232\,
            lcout => \ALU.madd_223_0\,
            ltout => \ALU.madd_223_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_238_0_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16324\,
            in2 => \N__16262\,
            in3 => \N__16308\,
            lcout => \ALU.madd_238_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_12_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__17299\,
            in1 => \N__17224\,
            in2 => \N__16190\,
            in3 => \N__16259\,
            lcout => \ALU.N_1559_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_165_0_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__40085\,
            in1 => \N__37214\,
            in2 => \_gnd_net_\,
            in3 => \N__16240\,
            lcout => \ALU.madd_165_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_213_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010011100"
        )
    port map (
            in0 => \N__46463\,
            in1 => \N__46693\,
            in2 => \N__40409\,
            in3 => \N__28027\,
            lcout => \ALU.madd_213_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIU9R47_5_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__21766\,
            in1 => \N__40362\,
            in2 => \N__29967\,
            in3 => \N__21700\,
            lcout => \ALU.a5_b_5\,
            ltout => \ALU.a5_b_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_175_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100000"
        )
    port map (
            in0 => \N__41943\,
            in1 => \N__47088\,
            in2 => \N__16211\,
            in3 => \N__16207\,
            lcout => \ALU.madd_175\,
            ltout => \ALU.madd_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_232_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__17554\,
            in1 => \N__16156\,
            in2 => \N__16193\,
            in3 => \N__16393\,
            lcout => \ALU.madd_232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI07LK7_4_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23486\,
            in1 => \N__46962\,
            in2 => \N__26576\,
            in3 => \N__23569\,
            lcout => \ALU.a7_b_4\,
            ltout => \ALU.a7_b_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_228_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16163\,
            in1 => \N__16157\,
            in2 => \N__16148\,
            in3 => \N__16394\,
            lcout => \ALU.madd_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAMNM3_5_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__21699\,
            in1 => \N__21765\,
            in2 => \_gnd_net_\,
            in3 => \N__25229\,
            lcout => \ALU.N_225_0\,
            ltout => \ALU.N_225_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_64_0_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011000110"
        )
    port map (
            in0 => \N__36962\,
            in1 => \N__41942\,
            in2 => \N__16385\,
            in3 => \N__42689\,
            lcout => \ALU.madd_64_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_290_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18475\,
            in1 => \N__17648\,
            in2 => \_gnd_net_\,
            in3 => \N__16278\,
            lcout => OPEN,
            ltout => \ALU.madd_290_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_299_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__16496\,
            in1 => \N__16511\,
            in2 => \N__16382\,
            in3 => \N__16556\,
            lcout => \ALU.madd_299\,
            ltout => \ALU.madd_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_360_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16379\,
            in3 => \N__16368\,
            lcout => \ALU.madd_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_13_ma_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16345\,
            lcout => \ALU.madd_cry_13_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_242_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011101000"
        )
    port map (
            in0 => \N__16334\,
            in1 => \N__16325\,
            in2 => \N__16449\,
            in3 => \N__16313\,
            lcout => \ALU.madd_242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_265_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010100110"
        )
    port map (
            in0 => \N__40419\,
            in1 => \N__42933\,
            in2 => \N__21486\,
            in3 => \N__47087\,
            lcout => \ALU.madd_265_0\,
            ltout => \ALU.madd_265_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_280_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17380\,
            in1 => \N__23775\,
            in2 => \N__16286\,
            in3 => \N__19919\,
            lcout => \ALU.madd_280\,
            ltout => \ALU.madd_280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_295_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17647\,
            in1 => \N__18474\,
            in2 => \N__16559\,
            in3 => \N__16555\,
            lcout => \ALU.madd_295_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_11_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__16544\,
            in1 => \N__16409\,
            in2 => \N__16475\,
            in3 => \_gnd_net_\,
            lcout => \ALU.madd_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI698B8_7_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__19849\,
            in1 => \N__42906\,
            in2 => \N__26496\,
            in3 => \N__19091\,
            lcout => \ALU.a4_b_7\,
            ltout => \ALU.a4_b_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_233_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16688\,
            in1 => \N__17566\,
            in2 => \N__16517\,
            in3 => \N__16759\,
            lcout => \ALU.madd_233\,
            ltout => \ALU.madd_233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_247_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011101000"
        )
    port map (
            in0 => \N__16604\,
            in1 => \N__16450\,
            in2 => \N__16514\,
            in3 => \N__16426\,
            lcout => \ALU.madd_247\,
            ltout => \ALU.madd_247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_300_0_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16510\,
            in1 => \N__16495\,
            in2 => \N__16484\,
            in3 => \N__16481\,
            lcout => \ALU.madd_N_10\,
            ltout => \ALU.madd_N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_12_l_fx_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__16466\,
            in1 => \N__25933\,
            in2 => \N__16460\,
            in3 => \N__16457\,
            lcout => \ALU.madd_axb_12_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_243_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16451\,
            in1 => \N__16603\,
            in2 => \N__16430\,
            in3 => \N__16415\,
            lcout => \ALU.madd_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0B2B8_7_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110010100011"
        )
    port map (
            in0 => \N__19838\,
            in1 => \N__19081\,
            in2 => \N__26495\,
            in3 => \N__46912\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITAM9D_7_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16643\,
            in3 => \N__47049\,
            lcout => \ALU.d_RNITAM9DZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGF4I7_8_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000000000"
        )
    port map (
            in0 => \N__24298\,
            in1 => \N__18730\,
            in2 => \N__18674\,
            in3 => \N__37985\,
            lcout => \ALU.a0_b_8\,
            ltout => \ALU.a0_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_103_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__17624\,
            in1 => \N__37503\,
            in2 => \N__16640\,
            in3 => \N__47050\,
            lcout => \ALU.madd_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITVJU4_7_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__19837\,
            in1 => \N__24297\,
            in2 => \_gnd_net_\,
            in3 => \N__19080\,
            lcout => \ALU.N_213_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_148_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__16636\,
            in1 => \N__16792\,
            in2 => \_gnd_net_\,
            in3 => \N__16625\,
            lcout => \ALU.madd_148\,
            ltout => \ALU.madd_148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_195_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011101000"
        )
    port map (
            in0 => \N__16590\,
            in1 => \N__16572\,
            in2 => \N__16607\,
            in3 => \_gnd_net_\,
            lcout => \ALU.madd_247_0_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_143_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000001000"
        )
    port map (
            in0 => \N__37986\,
            in1 => \N__22085\,
            in2 => \N__22073\,
            in3 => \N__21977\,
            lcout => \ALU.madd_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_181_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__16741\,
            in1 => \N__16702\,
            in2 => \N__16732\,
            in3 => \N__20329\,
            lcout => \ALU.madd_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_129_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101100110"
        )
    port map (
            in0 => \N__17717\,
            in1 => \N__16781\,
            in2 => \N__28088\,
            in3 => \N__42973\,
            lcout => \ALU.madd_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6I7F7_4_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__40368\,
            in2 => \N__24283\,
            in3 => \N__23573\,
            lcout => \ALU.a5_b_4\,
            ltout => \ALU.a5_b_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_133_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__17716\,
            in1 => \N__42972\,
            in2 => \N__16775\,
            in3 => \N__28071\,
            lcout => \ALU.madd_133\,
            ltout => \ALU.madd_133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_185_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101000"
        )
    port map (
            in0 => \N__16725\,
            in1 => \N__16701\,
            in2 => \N__16772\,
            in3 => \N__20330\,
            lcout => \ALU.madd_237_0_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_23_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__38318\,
            in1 => \N__39853\,
            in2 => \_gnd_net_\,
            in3 => \N__20375\,
            lcout => OPEN,
            ltout => \ALU.madd_128_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_7_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101000"
        )
    port map (
            in0 => \N__16742\,
            in1 => \N__16733\,
            in2 => \N__16706\,
            in3 => \N__16703\,
            lcout => OPEN,
            ltout => \ALU.madd_237_0_tz_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_6_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17675\,
            in1 => \_gnd_net_\,
            in2 => \N__16691\,
            in3 => \N__16687\,
            lcout => \ALU.N_1537_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m48_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111101101000"
        )
    port map (
            in0 => \N__22698\,
            in1 => \N__22408\,
            in2 => \N__22600\,
            in3 => \N__48029\,
            lcout => OPEN,
            ltout => \ALU.i6_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m50_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__22324\,
            in1 => \N__22594\,
            in2 => \N__16646\,
            in3 => \N__22699\,
            lcout => OPEN,
            ltout => \N_51_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_0_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__33275\,
            in1 => \N__33434\,
            in2 => \N__16820\,
            in3 => \N__48030\,
            lcout => \aluOperation_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m55_am_LC_3_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__22407\,
            in1 => \N__22322\,
            in2 => \N__22601\,
            in3 => \N__17771\,
            lcout => \ALU.m55_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m641_ns_1_LC_3_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111111"
        )
    port map (
            in0 => \N__22697\,
            in1 => \N__22323\,
            in2 => \N__33303\,
            in3 => \N__20483\,
            lcout => \ALU.m641_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m645_ns_1_LC_3_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000001111"
        )
    port map (
            in0 => \N__22321\,
            in1 => \N__22696\,
            in2 => \N__43180\,
            in3 => \N__33271\,
            lcout => \ALU.m645_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_cnv_0_LC_3_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17924\,
            in1 => \N__20459\,
            in2 => \N__17888\,
            in3 => \N__17839\,
            lcout => \ALU.h_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.results_e_0_1_LC_3_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16952\,
            lcout => \aluResults_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47643\,
            ce => \N__16843\,
            sr => \_gnd_net_\
        );

    \CONTROL.results_e_0_2_LC_3_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16817\,
            lcout => \aluResults_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47643\,
            ce => \N__16843\,
            sr => \_gnd_net_\
        );

    \ALU.m16_LC_3_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__22387\,
            in1 => \N__22276\,
            in2 => \N__22584\,
            in3 => \N__22676\,
            lcout => \N_723\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m55_bm_LC_3_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011111"
        )
    port map (
            in0 => \N__22677\,
            in1 => \N__22388\,
            in2 => \N__22298\,
            in3 => \N__22555\,
            lcout => \ALU.m55_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m661_LC_3_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__22386\,
            in1 => \N__22275\,
            in2 => \N__22582\,
            in3 => \N__22675\,
            lcout => \N_662_0\,
            ltout => \N_662_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_cnv_0_LC_3_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100000000"
        )
    port map (
            in0 => \N__16889\,
            in1 => \N__33245\,
            in2 => \N__16892\,
            in3 => \N__34604\,
            lcout => \CONTROL.operand1_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m664_LC_3_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100101011001"
        )
    port map (
            in0 => \N__22385\,
            in1 => \N__22274\,
            in2 => \N__22583\,
            in3 => \N__22674\,
            lcout => \N_665_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m300_ns_LC_3_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010010111111"
        )
    port map (
            in0 => \N__16877\,
            in1 => \N__22320\,
            in2 => \N__33302\,
            in3 => \N__44324\,
            lcout => OPEN,
            ltout => \N_301_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_3_LC_3_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__44325\,
            in1 => \_gnd_net_\,
            in2 => \N__16883\,
            in3 => \N__22124\,
            lcout => \aluParams_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47649\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m667_LC_3_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100101011011"
        )
    port map (
            in0 => \N__22405\,
            in1 => \N__22319\,
            in2 => \N__22525\,
            in3 => \N__22685\,
            lcout => OPEN,
            ltout => \N_668_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_cnv_0_LC_3_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000010"
        )
    port map (
            in0 => \N__34617\,
            in1 => \N__33264\,
            in2 => \N__16880\,
            in3 => \N__16863\,
            lcout => \CONTROL.aluParams_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m300_ns_1_LC_3_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111110101"
        )
    port map (
            in0 => \N__22406\,
            in1 => \N__22686\,
            in2 => \N__33301\,
            in3 => \N__18065\,
            lcout => \ALU.m300_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m669_LC_3_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111000001"
        )
    port map (
            in0 => \N__22684\,
            in1 => \N__22497\,
            in2 => \N__22325\,
            in3 => \N__22404\,
            lcout => OPEN,
            ltout => \N_670_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.results_cnv_0_LC_3_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101100000000"
        )
    port map (
            in0 => \N__16864\,
            in1 => \N__33260\,
            in2 => \N__16850\,
            in3 => \N__34616\,
            lcout => \CONTROL.results_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1M3JE_14_LC_3_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16901\,
            in2 => \_gnd_net_\,
            in3 => \N__21312\,
            lcout => \ALU.d_RNI1M3JEZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKNU29_14_LC_3_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011000011"
        )
    port map (
            in0 => \N__17811\,
            in1 => \N__40615\,
            in2 => \N__30646\,
            in3 => \N__26375\,
            lcout => \ALU.un2_addsub_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m636_LC_3_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001100"
        )
    port map (
            in0 => \N__22715\,
            in1 => \N__22419\,
            in2 => \N__22526\,
            in3 => \N__22285\,
            lcout => \ALU.N_724\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5SME5_14_LC_3_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010001110100"
        )
    port map (
            in0 => \N__17812\,
            in1 => \N__26380\,
            in2 => \N__30647\,
            in3 => \_gnd_net_\,
            lcout => \ALU.N_171_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9G6T4_9_LC_3_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__20870\,
            in1 => \N__26379\,
            in2 => \_gnd_net_\,
            in3 => \N__21094\,
            lcout => \ALU.N_207_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILOIL8_9_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110010100011"
        )
    port map (
            in0 => \N__21093\,
            in1 => \N__20869\,
            in2 => \N__26445\,
            in3 => \N__39847\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6B7KD_9_LC_3_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16895\,
            in3 => \N__22065\,
            lcout => \ALU.d_RNI6B7KDZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIF9794_9_LC_3_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__21095\,
            in1 => \N__29405\,
            in2 => \_gnd_net_\,
            in3 => \N__39848\,
            lcout => \ALU.N_274_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m252_LC_3_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__19630\,
            in1 => \N__19651\,
            in2 => \_gnd_net_\,
            in3 => \N__21563\,
            lcout => \ALU.N_253_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_362_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__40599\,
            in1 => \N__18835\,
            in2 => \N__38337\,
            in3 => \N__18151\,
            lcout => \ALU.madd_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_366_LC_3_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__18836\,
            in1 => \N__38322\,
            in2 => \N__18155\,
            in3 => \N__40600\,
            lcout => \ALU.madd_366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_0_ma_LC_3_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37471\,
            lcout => \ALU.madd_cry_0_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIH1R53_1_LC_3_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__37472\,
            in1 => \_gnd_net_\,
            in2 => \N__29434\,
            in3 => \N__23342\,
            lcout => \ALU.N_292_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI21MU3_6_LC_3_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__26283\,
            in1 => \N__29413\,
            in2 => \_gnd_net_\,
            in3 => \N__46670\,
            lcout => \ALU.N_291_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICCNU3_7_LC_3_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__46966\,
            in1 => \_gnd_net_\,
            in2 => \N__29433\,
            in3 => \N__19822\,
            lcout => \ALU.N_264_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAB477_6_LC_3_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43688\,
            in1 => \N__46965\,
            in2 => \_gnd_net_\,
            in3 => \N__46669\,
            lcout => \ALU.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIGTNC7_13_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40763\,
            in2 => \_gnd_net_\,
            in3 => \N__37759\,
            lcout => \ALU.a13_b_1\,
            ltout => \ALU.a13_b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_376_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010100000"
        )
    port map (
            in0 => \N__17006\,
            in1 => \N__21296\,
            in2 => \N__16904\,
            in3 => \N__38026\,
            lcout => \ALU.madd_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDU4G5_14_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__17802\,
            in1 => \N__24234\,
            in2 => \_gnd_net_\,
            in3 => \N__30634\,
            lcout => \ALU.N_171_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m168_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001111111"
        )
    port map (
            in0 => \N__30201\,
            in1 => \N__25205\,
            in2 => \N__16997\,
            in3 => \N__29740\,
            lcout => \ALU.N_169_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIDMS7_3_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23920\,
            in1 => \N__39375\,
            in2 => \N__29914\,
            in3 => \N__24029\,
            lcout => \ALU.a11_b_3\,
            ltout => \ALU.a11_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_372_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101011010"
        )
    port map (
            in0 => \N__17155\,
            in1 => \N__21297\,
            in2 => \N__17000\,
            in3 => \N__38027\,
            lcout => \ALU.madd_372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_30_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__41219\,
            in1 => \N__16996\,
            in2 => \N__41477\,
            in3 => \N__16981\,
            lcout => \ctrlOut_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__41056\,
            sr => \_gnd_net_\
        );

    \testWord_14_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__16980\,
            in1 => \N__41438\,
            in2 => \N__16948\,
            in3 => \N__41218\,
            lcout => \testWordZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47669\,
            ce => \N__41056\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI05GC8_7_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__19842\,
            in1 => \N__19102\,
            in2 => \N__30012\,
            in3 => \N__46728\,
            lcout => \ALU.a6_b_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN9HA7_6_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__26732\,
            in1 => \N__26276\,
            in2 => \N__29956\,
            in3 => \N__46943\,
            lcout => \ALU.a7_b_6\,
            ltout => \ALU.a7_b_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_320_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__16928\,
            in1 => \N__40082\,
            in2 => \N__16931\,
            in3 => \N__28085\,
            lcout => \ALU.madd_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_392_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16910\,
            in1 => \N__19733\,
            in2 => \_gnd_net_\,
            in3 => \N__18317\,
            lcout => \ALU.madd_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_324_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__16927\,
            in1 => \N__40083\,
            in2 => \N__16919\,
            in3 => \N__28086\,
            lcout => \ALU.madd_324_0\,
            ltout => \ALU.madd_324_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_396_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19732\,
            in2 => \N__17069\,
            in3 => \N__18316\,
            lcout => \ALU.madd_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGS0L7_6_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__26277\,
            in1 => \N__40081\,
            in2 => \N__30013\,
            in3 => \N__26731\,
            lcout => \ALU.a8_b_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_372_0_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010110100"
        )
    port map (
            in0 => \N__21311\,
            in1 => \N__38035\,
            in2 => \N__39396\,
            in3 => \N__41736\,
            lcout => \ALU.madd_372_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_21_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011111101000"
        )
    port map (
            in0 => \N__17066\,
            in1 => \N__17171\,
            in2 => \N__17015\,
            in3 => \N__17057\,
            lcout => \ALU.madd_484_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1S6M7_5_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__21785\,
            in1 => \N__39808\,
            in2 => \N__30022\,
            in3 => \N__21721\,
            lcout => \ALU.a9_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_411_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__17125\,
            in1 => \N__17144\,
            in2 => \_gnd_net_\,
            in3 => \N__17137\,
            lcout => OPEN,
            ltout => \ALU.madd_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_24_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17051\,
            in1 => \N__17114\,
            in2 => \N__17045\,
            in3 => \N__18275\,
            lcout => \ALU.madd_484_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_381_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__17023\,
            in1 => \N__27554\,
            in2 => \N__17036\,
            in3 => \N__42675\,
            lcout => \ALU.madd_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_377_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__42676\,
            in1 => \N__17035\,
            in2 => \N__27594\,
            in3 => \N__17024\,
            lcout => \ALU.madd_377\,
            ltout => \ALU.madd_377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_397_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17177\,
            in1 => \N__17170\,
            in2 => \N__17162\,
            in3 => \N__17159\,
            lcout => \ALU.madd_397\,
            ltout => \ALU.madd_397_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_407_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17138\,
            in1 => \_gnd_net_\,
            in2 => \N__17129\,
            in3 => \N__17126\,
            lcout => \ALU.madd_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_406_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__17105\,
            in1 => \N__18344\,
            in2 => \_gnd_net_\,
            in3 => \N__17098\,
            lcout => \ALU.madd_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0PL97_8_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__18738\,
            in1 => \N__26514\,
            in2 => \N__18669\,
            in3 => \N__40430\,
            lcout => OPEN,
            ltout => \ALU.a5_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_329_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100000"
        )
    port map (
            in0 => \N__42927\,
            in1 => \N__22064\,
            in2 => \N__17108\,
            in3 => \N__17431\,
            lcout => \ALU.madd_329_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_387_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18358\,
            in1 => \N__18241\,
            in2 => \_gnd_net_\,
            in3 => \N__18265\,
            lcout => \ALU.madd_387\,
            ltout => \ALU.madd_387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_402_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17099\,
            in2 => \N__17090\,
            in3 => \N__18343\,
            lcout => \ALU.madd_402\,
            ltout => \ALU.madd_402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_412_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18430\,
            in2 => \N__17081\,
            in3 => \N__17407\,
            lcout => \ALU.madd_412\,
            ltout => \ALU.madd_412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_417_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17078\,
            in2 => \N__17072\,
            in3 => \N__17344\,
            lcout => \ALU.madd_329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_573_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__17345\,
            in1 => \N__17336\,
            in2 => \_gnd_net_\,
            in3 => \N__17330\,
            lcout => \ALU.madd_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_9_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38329\,
            in1 => \N__25372\,
            in2 => \N__37000\,
            in3 => \N__39594\,
            lcout => \ALU.madd_141_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_270_0_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__25373\,
            in1 => \N__17279\,
            in2 => \N__17252\,
            in3 => \N__38330\,
            lcout => \ALU.madd_270_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_0_rep1_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34681\,
            in1 => \N__34798\,
            in2 => \N__31250\,
            in3 => \N__41112\,
            lcout => \aluOperand2_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_207_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__39394\,
            in1 => \N__19997\,
            in2 => \N__38339\,
            in3 => \N__19961\,
            lcout => \ALU.madd_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_250_0_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__27539\,
            in1 => \N__39593\,
            in2 => \N__36999\,
            in3 => \N__37232\,
            lcout => \ALU.madd_250_0\,
            ltout => \ALU.madd_250_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_250_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25354\,
            in2 => \N__17273\,
            in3 => \N__38331\,
            lcout => \ALU.madd_250\,
            ltout => \ALU.madd_250_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_274_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17250\,
            in2 => \N__17228\,
            in3 => \N__17211\,
            lcout => \ALU.madd_274\,
            ltout => \ALU.madd_274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_344_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011101000"
        )
    port map (
            in0 => \N__17490\,
            in1 => \N__17456\,
            in2 => \N__17438\,
            in3 => \N__17435\,
            lcout => \ALU.madd_344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_25_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__23617\,
            in1 => \N__38029\,
            in2 => \N__24065\,
            in3 => \N__28026\,
            lcout => \ALU.madd_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_29_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001000000"
        )
    port map (
            in0 => \N__28025\,
            in1 => \N__24064\,
            in2 => \N__38046\,
            in3 => \N__23618\,
            lcout => \ALU.madd_29\,
            ltout => \ALU.madd_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_47_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__18905\,
            in1 => \N__38033\,
            in2 => \N__17396\,
            in3 => \N__46473\,
            lcout => \ALU.madd_47\,
            ltout => \ALU.madd_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_5_l_fx_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__18782\,
            in1 => \N__26183\,
            in2 => \N__17393\,
            in3 => \N__18791\,
            lcout => \ALU.madd_axb_5_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_4_l_fx_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18790\,
            in1 => \N__25741\,
            in2 => \_gnd_net_\,
            in3 => \N__18781\,
            lcout => \ALU.madd_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_284_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__17390\,
            in1 => \N__23779\,
            in2 => \N__17381\,
            in3 => \N__19915\,
            lcout => \ALU.madd_284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_309_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__37205\,
            in1 => \N__39322\,
            in2 => \N__35069\,
            in3 => \N__18818\,
            lcout => \ALU.madd_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGGQ26_1_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37485\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37204\,
            lcout => \ALU.a1_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIG1A7_6_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__26284\,
            in1 => \N__36958\,
            in2 => \N__30054\,
            in3 => \N__26729\,
            lcout => \ALU.a2_b_6\,
            ltout => \ALU.a2_b_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_99_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__37486\,
            in1 => \N__17612\,
            in2 => \N__17600\,
            in3 => \N__47096\,
            lcout => \ALU.madd_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILIL37_6_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__26285\,
            in1 => \N__40410\,
            in2 => \N__30055\,
            in3 => \N__26730\,
            lcout => \ALU.a5_b_6\,
            ltout => \ALU.a5_b_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_217_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__17532\,
            in1 => \N__46961\,
            in2 => \N__17597\,
            in3 => \N__42666\,
            lcout => \ALU.madd_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_42_0_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011010010"
        )
    port map (
            in0 => \N__37487\,
            in1 => \N__28034\,
            in2 => \N__36998\,
            in3 => \N__42667\,
            lcout => \ALU.madd_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN9H73_5_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__28541\,
            in1 => \N__31655\,
            in2 => \N__33096\,
            in3 => \N__28883\,
            lcout => \ALU.operand2_5\,
            ltout => \ALU.operand2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINMLB7_5_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101000"
        )
    port map (
            in0 => \N__46672\,
            in1 => \N__30032\,
            in2 => \N__17594\,
            in3 => \N__21784\,
            lcout => \ALU.a6_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_176_0_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011000110"
        )
    port map (
            in0 => \N__36964\,
            in1 => \N__37488\,
            in2 => \N__21485\,
            in3 => \N__22066\,
            lcout => \ALU.madd_176_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_218_0_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101000100"
        )
    port map (
            in0 => \N__22067\,
            in1 => \N__36966\,
            in2 => \N__21487\,
            in3 => \N__41927\,
            lcout => \ALU.madd_218_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_275_0_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011111101000"
        )
    port map (
            in0 => \N__17555\,
            in1 => \N__17533\,
            in2 => \N__17509\,
            in3 => \N__18525\,
            lcout => \ALU.madd_275_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_42_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__37489\,
            in1 => \N__23605\,
            in2 => \N__24376\,
            in3 => \N__28035\,
            lcout => \ALU.madd_42\,
            ltout => \ALU.madd_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m3_2_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19003\,
            in2 => \N__17639\,
            in3 => \N__19022\,
            lcout => \ALU.madd_i1_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_52_0_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__19004\,
            in1 => \_gnd_net_\,
            in2 => \N__24377\,
            in3 => \N__17636\,
            lcout => \ALU.madd_52_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_1_ma_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37490\,
            lcout => \ALU.madd_cry_1_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVQ5R6_2_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36965\,
            in2 => \_gnd_net_\,
            in3 => \N__37702\,
            lcout => \ALU.a2_b_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFDNC8_7_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__19819\,
            in1 => \N__42905\,
            in2 => \N__30056\,
            in3 => \N__19085\,
            lcout => \ALU.a4_b_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIM09H_7_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27875\,
            in1 => \N__28805\,
            in2 => \_gnd_net_\,
            in3 => \N__32079\,
            lcout => OPEN,
            ltout => \ALU.e_RNIM09HZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIKJH32_7_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__33085\,
            in1 => \N__34512\,
            in2 => \N__17630\,
            in3 => \N__31670\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIULB84_7_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__32963\,
            in1 => \N__45203\,
            in2 => \N__17627\,
            in3 => \N__26897\,
            lcout => \ALU.operand2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g1_2_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001111111111"
        )
    port map (
            in0 => \N__18673\,
            in1 => \N__18740\,
            in2 => \N__30057\,
            in3 => \N__41919\,
            lcout => OPEN,
            ltout => \ALU.g1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_25_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010001001011"
        )
    port map (
            in0 => \N__22072\,
            in1 => \N__36963\,
            in2 => \N__17684\,
            in3 => \N__17681\,
            lcout => \ALU.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIL5C37_5_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110010100011"
        )
    port map (
            in0 => \N__21786\,
            in1 => \N__21722\,
            in2 => \N__26603\,
            in3 => \N__40367\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVR3QA_5_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17666\,
            in3 => \N__28070\,
            lcout => \ALU.d_RNIVR3QAZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICFBS3_5_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__21787\,
            in1 => \N__21723\,
            in2 => \_gnd_net_\,
            in3 => \N__26575\,
            lcout => \ALU.N_225_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILT5T4_7_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__19089\,
            in1 => \N__26564\,
            in2 => \_gnd_net_\,
            in3 => \N__19821\,
            lcout => \ALU.N_213_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN01B8_7_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000100000"
        )
    port map (
            in0 => \N__46616\,
            in1 => \N__19820\,
            in2 => \N__26604\,
            in3 => \N__19090\,
            lcout => \ALU.a6_b_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNII0KR6_6_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46615\,
            in2 => \_gnd_net_\,
            in3 => \N__38291\,
            lcout => \ALU.a6_b_0\,
            ltout => \ALU.a6_b_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_41_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__18863\,
            in1 => \N__40366\,
            in2 => \N__17651\,
            in3 => \N__37730\,
            lcout => \ALU.madd_41\,
            ltout => \ALU.madd_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_69_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__19036\,
            in1 => \N__37514\,
            in2 => \N__17726\,
            in3 => \N__46448\,
            lcout => \ALU.madd_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_46_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__23606\,
            in1 => \N__37513\,
            in2 => \N__24375\,
            in3 => \N__28087\,
            lcout => \ALU.madd_46\,
            ltout => \ALU.madd_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_76_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000001000000"
        )
    port map (
            in0 => \N__41721\,
            in1 => \N__42995\,
            in2 => \N__17723\,
            in3 => \N__18940\,
            lcout => \ALU.madd_39\,
            ltout => \ALU.madd_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_118_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101000"
        )
    port map (
            in0 => \N__20366\,
            in1 => \N__17702\,
            in2 => \N__17720\,
            in3 => \N__19226\,
            lcout => \ALU.madd_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDAJB7_3_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__23945\,
            in1 => \N__24030\,
            in2 => \N__24317\,
            in3 => \N__46671\,
            lcout => \ALU.a6_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_78_0_tz_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110110"
        )
    port map (
            in0 => \N__18939\,
            in1 => \N__42994\,
            in2 => \N__19217\,
            in3 => \N__41720\,
            lcout => OPEN,
            ltout => \ALU.madd_78_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_78_0_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17705\,
            in3 => \N__20414\,
            lcout => \ALU.madd_78_0\,
            ltout => \ALU.madd_78_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_114_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__20365\,
            in1 => \N__17696\,
            in2 => \N__17690\,
            in3 => \N__19225\,
            lcout => \ALU.madd_114\,
            ltout => \ALU.madd_114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_8_l_fx_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \N__26068\,
            in1 => \N__19307\,
            in2 => \N__17687\,
            in3 => \N__18872\,
            lcout => \ALU.madd_axb_8_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testClock_RNIAQVB_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__41338\,
            in1 => \N__30290\,
            in2 => \N__30780\,
            in3 => \N__17743\,
            lcout => \testClock_0\,
            ltout => \testClock_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_cnv_0_0_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__17744\,
            in1 => \_gnd_net_\,
            in2 => \N__17777\,
            in3 => \N__17764\,
            lcout => \ALU.a_cnv_0Z0Z_0\,
            ltout => \ALU.a_cnv_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_cnv_0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20435\,
            in1 => \N__17852\,
            in2 => \N__17774\,
            in3 => \N__17925\,
            lcout => \ALU.a_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m52_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__22438\,
            in1 => \N__22729\,
            in2 => \N__22599\,
            in3 => \N__44038\,
            lcout => \ALU.N_53_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testClock_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__41340\,
            in1 => \N__30291\,
            in2 => \N__30782\,
            in3 => \N__17746\,
            lcout => \testClockZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_cnv_0_0_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17745\,
            in1 => \N__17765\,
            in2 => \_gnd_net_\,
            in3 => \N__17753\,
            lcout => \ALU.b_cnv_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_2_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100001010000"
        )
    port map (
            in0 => \N__41339\,
            in1 => \N__21895\,
            in2 => \N__30781\,
            in3 => \N__30292\,
            lcout => \testStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_cnv_0_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17938\,
            in1 => \N__17847\,
            in2 => \N__17927\,
            in3 => \N__20455\,
            lcout => \ALU.e_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_cnv_0_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20454\,
            in1 => \N__17921\,
            in2 => \N__17853\,
            in3 => \N__17937\,
            lcout => \ALU.c_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.G_566_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41399\,
            in1 => \N__30314\,
            in2 => \N__30783\,
            in3 => \N__17747\,
            lcout => \G_566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_cnv_0_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17926\,
            in1 => \N__17939\,
            in2 => \N__17855\,
            in3 => \N__20458\,
            lcout => \ALU.g_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_cnv_0_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17917\,
            in1 => \N__20453\,
            in2 => \N__17883\,
            in3 => \N__17840\,
            lcout => \ALU.b_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_cnv_0_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17882\,
            in1 => \N__17922\,
            in2 => \N__17854\,
            in3 => \N__20457\,
            lcout => \ALU.d_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_cnv_0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17923\,
            in1 => \N__20456\,
            in2 => \N__17884\,
            in3 => \N__17848\,
            lcout => \ALU.f_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIEP354_14_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__17813\,
            in1 => \N__40616\,
            in2 => \_gnd_net_\,
            in3 => \N__29377\,
            lcout => OPEN,
            ltout => \ALU.c_RNIEP354Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI25K7D_14_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43109\,
            in2 => \N__17786\,
            in3 => \N__17783\,
            lcout => \ALU.a_15_m3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJENJ8_0_15_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__38432\,
            in1 => \N__38647\,
            in2 => \N__39082\,
            in3 => \N__44334\,
            lcout => \ALU.c_RNIJENJ8_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJENJ8_15_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000101"
        )
    port map (
            in0 => \N__38646\,
            in1 => \N__39053\,
            in2 => \N__44403\,
            in3 => \N__38431\,
            lcout => \ALU.rshift_15_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIR45G7_6_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__43697\,
            in1 => \N__46960\,
            in2 => \N__39081\,
            in3 => \N__46735\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIS6U9F_9_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__39851\,
            in1 => \N__39054\,
            in2 => \N__17981\,
            in3 => \N__40071\,
            lcout => \ALU.N_474\,
            ltout => \ALU.N_474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNII2IF91_9_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__44323\,
            in1 => \N__19445\,
            in2 => \N__17978\,
            in3 => \N__17975\,
            lcout => OPEN,
            ltout => \ALU.rshift_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIL01TD1_6_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43110\,
            in2 => \N__17969\,
            in3 => \N__17966\,
            lcout => \ALU.d_RNIL01TD1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIKJTS7_15_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__40619\,
            in1 => \N__39076\,
            in2 => \N__32665\,
            in3 => \N__43667\,
            lcout => \ALU.lshift_3_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3FQF1_14_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35401\,
            in1 => \N__33692\,
            in2 => \N__19475\,
            in3 => \N__31556\,
            lcout => \ALU.N_713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNITDBD1_14_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__28298\,
            in1 => \N__35761\,
            in2 => \N__28322\,
            in3 => \N__35588\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI81K02_14_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35402\,
            in1 => \N__30620\,
            in2 => \N__17957\,
            in3 => \N__30596\,
            lcout => \ALU.N_761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIN38K3_15_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30556\,
            in1 => \N__30536\,
            in2 => \_gnd_net_\,
            in3 => \N__35243\,
            lcout => \ALU.aluOut_15\,
            ltout => \ALU.aluOut_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3QSJ7_15_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43653\,
            in2 => \N__17954\,
            in3 => \N__40618\,
            lcout => \ALU.N_590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFR7K3_14_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17951\,
            in1 => \N__17945\,
            in2 => \_gnd_net_\,
            in3 => \N__35242\,
            lcout => \ALU.aluOut_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_14_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__47292\,
            in1 => \N__44089\,
            in2 => \N__43919\,
            in3 => \N__43668\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI58CHC_14_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001100111"
        )
    port map (
            in0 => \N__47293\,
            in1 => \N__40617\,
            in2 => \N__18011\,
            in3 => \N__21304\,
            lcout => \ALU.a_15_m2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIB9KD11_11_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__38732\,
            in1 => \N__19463\,
            in2 => \N__44523\,
            in3 => \N__20789\,
            lcout => OPEN,
            ltout => \ALU.lshift_15_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAD5QQ1_0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__44491\,
            in1 => \N__39200\,
            in2 => \N__18008\,
            in3 => \N__39185\,
            lcout => OPEN,
            ltout => \ALU.lshift_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIEGAQ72_14_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44090\,
            in2 => \N__18005\,
            in3 => \N__18002\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFCGVL2_14_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46331\,
            in2 => \N__17996\,
            in3 => \N__17993\,
            lcout => \c_RNIFCGVL2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI63LF1_12_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__35910\,
            in1 => \N__28565\,
            in2 => \N__36005\,
            in3 => \N__28211\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBAHQ1_12_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35394\,
            in1 => \N__33962\,
            in2 => \N__17984\,
            in3 => \N__31286\,
            lcout => \ALU.N_711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIP9BD1_12_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__35762\,
            in1 => \N__28370\,
            in2 => \N__28349\,
            in3 => \N__35577\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0PJ02_12_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35395\,
            in1 => \N__25499\,
            in2 => \N__18170\,
            in3 => \N__28394\,
            lcout => OPEN,
            ltout => \ALU.N_759_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFEUU3_12_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18167\,
            in2 => \N__18161\,
            in3 => \N__35241\,
            lcout => \ALU.aluOut_12\,
            ltout => \ALU.aluOut_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIIUNC7_12_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__37245\,
            in1 => \_gnd_net_\,
            in2 => \N__18158\,
            in3 => \_gnd_net_\,
            lcout => \ALU.a12_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA6K08_4_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23446\,
            in1 => \N__39821\,
            in2 => \N__30014\,
            in3 => \N__23567\,
            lcout => \ALU.a9_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_20_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__18022\,
            in1 => \N__32292\,
            in2 => \N__41478\,
            in3 => \N__18138\,
            lcout => \ctrlOut_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47670\,
            ce => \N__41057\,
            sr => \_gnd_net_\
        );

    \ALU.m234_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111110101"
        )
    port map (
            in0 => \N__29681\,
            in1 => \N__18061\,
            in2 => \N__25164\,
            in3 => \N__30136\,
            lcout => \ALU.N_235_0\,
            ltout => \ALU.N_235_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRNNS7_3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__29955\,
            in1 => \N__25288\,
            in2 => \N__18029\,
            in3 => \N__24043\,
            lcout => OPEN,
            ltout => \ALU.a12_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_11_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__40626\,
            in1 => \N__23366\,
            in2 => \N__18026\,
            in3 => \N__37761\,
            lcout => \ALU.madd_484_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m228_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001111111"
        )
    port map (
            in0 => \N__30135\,
            in1 => \N__25118\,
            in2 => \N__18023\,
            in3 => \N__29682\,
            lcout => \ALU.N_229_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIOVJ78_3_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__24042\,
            in1 => \N__29954\,
            in2 => \N__23921\,
            in3 => \N__27587\,
            lcout => OPEN,
            ltout => \ALU.a10_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_319_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__37760\,
            in1 => \N__18326\,
            in2 => \N__18320\,
            in3 => \N__25289\,
            lcout => \ALU.madd_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_15_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18308\,
            in1 => \N__19499\,
            in2 => \N__20396\,
            in3 => \N__18299\,
            lcout => \ALU.madd_484_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_17_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19706\,
            in1 => \N__18293\,
            in2 => \_gnd_net_\,
            in3 => \N__20984\,
            lcout => OPEN,
            ltout => \ALU.madd_484_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_20_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18176\,
            in1 => \N__18221\,
            in2 => \N__18284\,
            in3 => \N__18281\,
            lcout => \ALU.madd_484_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_391_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__18362\,
            in1 => \_gnd_net_\,
            in2 => \N__18269\,
            in3 => \N__18245\,
            lcout => \ALU.madd_391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0B2B8_0_7_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010100000"
        )
    port map (
            in0 => \N__46907\,
            in1 => \N__19788\,
            in2 => \N__19106\,
            in3 => \N__26523\,
            lcout => OPEN,
            ltout => \ALU.a7_b_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_16_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011111101000"
        )
    port map (
            in0 => \N__18215\,
            in1 => \N__18203\,
            in2 => \N__18185\,
            in3 => \N__18182\,
            lcout => \ALU.madd_484_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIB0KD9_12_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111001010"
        )
    port map (
            in0 => \N__25462\,
            in1 => \N__20917\,
            in2 => \N__26597\,
            in3 => \N__25326\,
            lcout => OPEN,
            ltout => \ALU.un9_addsub_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFKNTE_12_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18368\,
            in3 => \N__40848\,
            lcout => \ALU.d_RNIFKNTEZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISHLE5_12_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110101"
        )
    port map (
            in0 => \N__25463\,
            in1 => \_gnd_net_\,
            in2 => \N__26596\,
            in3 => \N__20918\,
            lcout => \ALU.N_180_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIV96U8_13_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__25061\,
            in1 => \N__25008\,
            in2 => \N__30031\,
            in3 => \N__38002\,
            lcout => \ALU.d_RNIV96U8Z0Z_13\,
            ltout => \ALU.d_RNIV96U8Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_314_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__39448\,
            in1 => \N__36989\,
            in2 => \N__18365\,
            in3 => \N__18335\,
            lcout => \ALU.madd_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_310_0_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__37418\,
            in1 => \N__40847\,
            in2 => \N__37003\,
            in3 => \N__39447\,
            lcout => \ALU.madd_310_0\,
            ltout => \ALU.madd_310_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_334_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__18809\,
            in1 => \N__18419\,
            in2 => \N__18347\,
            in3 => \N__19677\,
            lcout => \ALU.madd_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIM558_12_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__20916\,
            in1 => \N__37417\,
            in2 => \N__30030\,
            in3 => \N__25461\,
            lcout => \ALU.a1_b_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO82C8_9_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__21098\,
            in1 => \N__20866\,
            in2 => \N__30050\,
            in3 => \N__36985\,
            lcout => OPEN,
            ltout => \ALU.a2_b_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_222_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__18575\,
            in1 => \N__42891\,
            in2 => \N__18329\,
            in3 => \N__47100\,
            lcout => \ALU.madd_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI885I7_8_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000000000"
        )
    port map (
            in0 => \N__24231\,
            in1 => \N__18739\,
            in2 => \N__18668\,
            in3 => \N__41941\,
            lcout => \ALU.a3_b_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_275_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__18482\,
            in1 => \_gnd_net_\,
            in2 => \N__18515\,
            in3 => \N__18550\,
            lcout => \ALU.madd_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_279_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__18549\,
            in1 => \N__18502\,
            in2 => \_gnd_net_\,
            in3 => \N__18481\,
            lcout => OPEN,
            ltout => \ALU.madd_279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_349_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011101000"
        )
    port map (
            in0 => \N__19684\,
            in1 => \N__18457\,
            in2 => \N__18443\,
            in3 => \N__18386\,
            lcout => \ALU.madd_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_330_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18418\,
            in1 => \N__18397\,
            in2 => \_gnd_net_\,
            in3 => \N__18805\,
            lcout => \ALU.madd_330_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIBLBO_10_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28601\,
            in1 => \N__23708\,
            in2 => \_gnd_net_\,
            in3 => \N__45136\,
            lcout => \ALU.a_RNIBLBOZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIF549_10_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45137\,
            in1 => \N__34282\,
            in2 => \_gnd_net_\,
            in3 => \N__34934\,
            lcout => OPEN,
            ltout => \ALU.c_RNIF549Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIVSRV1_10_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__32992\,
            in1 => \N__34513\,
            in2 => \N__18380\,
            in3 => \N__18377\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHGJR4_10_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__24404\,
            in1 => \N__32993\,
            in2 => \N__18371\,
            in3 => \N__26801\,
            lcout => \ALU.operand2_10\,
            ltout => \ALU.operand2_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIF6179_10_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__42787\,
            in1 => \N__30045\,
            in2 => \N__18839\,
            in3 => \N__20040\,
            lcout => \ALU.a4_b_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7U079_10_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__20041\,
            in1 => \N__41959\,
            in2 => \N__30058\,
            in3 => \N__20014\,
            lcout => \ALU.a3_b_10\,
            ltout => \ALU.a3_b_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_305_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__37218\,
            in1 => \N__39395\,
            in2 => \N__18812\,
            in3 => \N__35065\,
            lcout => \ALU.madd_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIV0CK1_7_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__45374\,
            in1 => \N__45356\,
            in2 => \N__35365\,
            in3 => \N__26906\,
            lcout => \ALU.N_754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_17_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__23188\,
            in1 => \N__22970\,
            in2 => \N__23209\,
            in3 => \N__23165\,
            lcout => \ALU.madd_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_5_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010001000"
        )
    port map (
            in0 => \N__24481\,
            in1 => \N__24460\,
            in2 => \N__37004\,
            in3 => \N__37651\,
            lcout => \ALU.madd_5\,
            ltout => \ALU.madd_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_19_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000011000000"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__20240\,
            in2 => \N__18794\,
            in3 => \N__41992\,
            lcout => \ALU.madd_19\,
            ltout => \ALU.madd_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_58_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18780\,
            in2 => \N__18767\,
            in3 => \N__18764\,
            lcout => \ALU.madd_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_a3_0_1_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27566\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37659\,
            lcout => \ALU.g0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKRRR6_4_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42789\,
            in2 => \_gnd_net_\,
            in3 => \N__37115\,
            lcout => \ALU.a4_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKT467_8_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40056\,
            in2 => \_gnd_net_\,
            in3 => \N__38225\,
            lcout => OPEN,
            ltout => \ALU.a8_b_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_93_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__46681\,
            in1 => \N__37116\,
            in2 => \N__18911\,
            in3 => \N__20566\,
            lcout => \ALU.madd_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4KLR6_7_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46813\,
            in2 => \_gnd_net_\,
            in3 => \N__37658\,
            lcout => \ALU.a7_b_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_23_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37660\,
            in1 => \N__42788\,
            in2 => \N__41975\,
            in3 => \N__37114\,
            lcout => OPEN,
            ltout => \ALU.madd_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_24_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__40425\,
            in1 => \N__20246\,
            in2 => \N__18908\,
            in3 => \N__38226\,
            lcout => \ALU.madd_24\,
            ltout => \ALU.madd_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_51_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101000"
        )
    port map (
            in0 => \N__18896\,
            in1 => \N__38001\,
            in2 => \N__18884\,
            in3 => \N__46462\,
            lcout => \ALU.madd_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m6_1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010001110001"
        )
    port map (
            in0 => \N__19150\,
            in1 => \N__19183\,
            in2 => \N__18881\,
            in3 => \N__19169\,
            lcout => \ALU.madd_i3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_37_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__40426\,
            in1 => \N__18862\,
            in2 => \N__18848\,
            in3 => \N__37653\,
            lcout => \ALU.madd_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_12_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__21635\,
            in1 => \N__21644\,
            in2 => \N__42971\,
            in3 => \N__38299\,
            lcout => \ALU.madd_12\,
            ltout => \ALU.madd_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_34_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18972\,
            in2 => \N__19025\,
            in3 => \N__20301\,
            lcout => \ALU.madd_34\,
            ltout => \ALU.madd_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_56_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19016\,
            in2 => \N__19007\,
            in3 => \N__19002\,
            lcout => \ALU.madd_56\,
            ltout => \ALU.madd_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_6_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19170\,
            in1 => \N__19151\,
            in2 => \N__18989\,
            in3 => \N__19184\,
            lcout => \ALU.madd_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_30_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__20302\,
            in1 => \_gnd_net_\,
            in2 => \N__18977\,
            in3 => \N__18952\,
            lcout => \ALU.madd_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_52_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001101010"
        )
    port map (
            in0 => \N__18986\,
            in1 => \N__18976\,
            in2 => \N__18956\,
            in3 => \N__20303\,
            lcout => \ALU.madd_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5R097_6_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001100011"
        )
    port map (
            in0 => \N__26282\,
            in1 => \N__46626\,
            in2 => \N__26602\,
            in3 => \N__26716\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGLK5B_6_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18944\,
            in3 => \N__46443\,
            lcout => \ALU.d_RNIGLK5BZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_74_0_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110111010010"
        )
    port map (
            in0 => \N__42926\,
            in1 => \N__41706\,
            in2 => \N__18941\,
            in3 => \N__20407\,
            lcout => \ALU.madd_74_0\,
            ltout => \ALU.madd_74_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_83_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__19216\,
            in1 => \N__19171\,
            in2 => \N__19229\,
            in3 => \N__19199\,
            lcout => \ALU.madd_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBQJS3_6_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__24263\,
            in1 => \N__26281\,
            in2 => \_gnd_net_\,
            in3 => \N__26715\,
            lcout => \ALU.N_219_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_79_0_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19215\,
            in1 => \N__19198\,
            in2 => \_gnd_net_\,
            in3 => \N__19190\,
            lcout => \ALU.madd_79_0\,
            ltout => \ALU.madd_79_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_88_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__19172\,
            in1 => \N__19149\,
            in2 => \N__19133\,
            in3 => \N__19130\,
            lcout => OPEN,
            ltout => \ALU.madd_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_7_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19306\,
            in2 => \N__19124\,
            in3 => \N__19121\,
            lcout => \ALU.madd_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_73_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100000"
        )
    port map (
            in0 => \N__37500\,
            in1 => \N__46449\,
            in2 => \N__19040\,
            in3 => \N__19115\,
            lcout => \ALU.madd_73\,
            ltout => \ALU.madd_73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_113_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19333\,
            in2 => \N__19109\,
            in3 => \N__21670\,
            lcout => \ALU.madd_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFCMC8_7_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__19853\,
            in1 => \N__19098\,
            in2 => \N__30059\,
            in3 => \N__37997\,
            lcout => \ALU.a0_b_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_154_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19367\,
            in1 => \N__20347\,
            in2 => \_gnd_net_\,
            in3 => \N__19348\,
            lcout => \ALU.madd_154\,
            ltout => \ALU.madd_154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_159_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19337\,
            in3 => \N__19269\,
            lcout => \ALU.madd_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_109_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19334\,
            in1 => \N__21671\,
            in2 => \_gnd_net_\,
            in3 => \N__19313\,
            lcout => \ALU.madd_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_9_ma_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19288\,
            in2 => \_gnd_net_\,
            in3 => \N__19270\,
            lcout => \ALU.madd_cry_9_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m271_ns_1_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110000000"
        )
    port map (
            in0 => \N__24922\,
            in1 => \N__30215\,
            in2 => \N__26627\,
            in3 => \N__29753\,
            lcout => \ALU.m271_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_e_0_3_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__33317\,
            in1 => \N__33385\,
            in2 => \N__19256\,
            in3 => \N__19406\,
            lcout => \aluOperation_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47622\,
            ce => \N__33442\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_m5s2_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20478\,
            in2 => \_gnd_net_\,
            in3 => \N__44029\,
            lcout => \ALU.a_15_sm3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m282_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22573\,
            lcout => \ALU.N_283_0\,
            ltout => \ALU.N_283_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_e_0_4_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000000100010"
        )
    port map (
            in0 => \N__33384\,
            in1 => \N__19244\,
            in2 => \N__19232\,
            in3 => \N__33318\,
            lcout => \aluOperation_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47622\,
            ce => \N__33442\,
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_e_0_2_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33316\,
            in1 => \N__19430\,
            in2 => \_gnd_net_\,
            in3 => \N__19418\,
            lcout => \aluOperation_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47622\,
            ce => \N__33442\,
            sr => \_gnd_net_\
        );

    \ALU.m650_ns_1_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110100001010"
        )
    port map (
            in0 => \N__45697\,
            in1 => \N__22441\,
            in2 => \N__22596\,
            in3 => \N__22724\,
            lcout => OPEN,
            ltout => \ALU.m650_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m650_ns_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101000010010"
        )
    port map (
            in0 => \N__22725\,
            in1 => \N__22299\,
            in2 => \N__19409\,
            in3 => \N__19405\,
            lcout => \N_727\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m14_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__22569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22439\,
            lcout => \ALU.N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_1_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33438\,
            in1 => \N__45698\,
            in2 => \N__33335\,
            in3 => \N__19397\,
            lcout => \aluOperation_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINJ76G_13_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38923\,
            in1 => \N__38755\,
            in2 => \_gnd_net_\,
            in3 => \N__38437\,
            lcout => OPEN,
            ltout => \ALU.N_577_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIN1J811_11_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38696\,
            in2 => \N__19391\,
            in3 => \N__20122\,
            lcout => \ALU.N_633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHDLLS_3_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38697\,
            in1 => \N__20147\,
            in2 => \_gnd_net_\,
            in3 => \N__22985\,
            lcout => OPEN,
            ltout => \ALU.N_528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8DL9U1_3_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__44480\,
            in1 => \_gnd_net_\,
            in2 => \N__19388\,
            in3 => \N__19378\,
            lcout => OPEN,
            ltout => \ALU.d_RNI8DL9U1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7AI932_0_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43097\,
            in2 => \N__19454\,
            in3 => \N__19601\,
            lcout => \ALU.a_15_m3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m713_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__44060\,
            in1 => \N__38922\,
            in2 => \_gnd_net_\,
            in3 => \N__43491\,
            lcout => \ALU.log_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID35S7_9_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40070\,
            in1 => \_gnd_net_\,
            in2 => \N__39837\,
            in3 => \N__43511\,
            lcout => \ALU.N_221\,
            ltout => \ALU.N_221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIDIAPG_11_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__39044\,
            in1 => \N__22934\,
            in2 => \N__19451\,
            in3 => \_gnd_net_\,
            lcout => \ALU.N_253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI30A98_13_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43545\,
            in1 => \N__40765\,
            in2 => \_gnd_net_\,
            in3 => \N__25340\,
            lcout => \ALU.N_588\,
            ltout => \ALU.N_588_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3FF6H_11_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39045\,
            in1 => \_gnd_net_\,
            in2 => \N__19448\,
            in3 => \N__20720\,
            lcout => \ALU.N_575\,
            ltout => \ALU.N_575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIMVPEP_15_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__38436\,
            in1 => \N__38652\,
            in2 => \N__19439\,
            in3 => \N__39046\,
            lcout => \ALU.N_635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1HUMG_11_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__19436\,
            in1 => \N__39384\,
            in2 => \N__39080\,
            in3 => \N__27608\,
            lcout => \ALU.N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIURRD4_0_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__39015\,
            in1 => \N__38653\,
            in2 => \N__43638\,
            in3 => \N__38028\,
            lcout => \ALU.N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUS558_9_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__43510\,
            in1 => \N__39795\,
            in2 => \N__39079\,
            in3 => \N__40069\,
            lcout => \ALU.rshift_3_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBIR3G_13_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__25343\,
            in1 => \N__19481\,
            in2 => \N__39077\,
            in3 => \N__40768\,
            lcout => \ALU.N_257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIQ3U41_14_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__35912\,
            in1 => \N__30728\,
            in2 => \N__35587\,
            in3 => \N__31385\,
            lcout => \ALU.dout_3_ns_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIK6K78_14_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__43673\,
            in1 => \N__40614\,
            in2 => \N__39078\,
            in3 => \N__40766\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIQIGEG_11_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__39387\,
            in1 => \N__39036\,
            in2 => \N__19466\,
            in3 => \N__25344\,
            lcout => \ALU.N_256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI30A98_0_13_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25342\,
            in1 => \_gnd_net_\,
            in2 => \N__43719\,
            in3 => \N__40767\,
            lcout => \ALU.N_225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIID898_0_11_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39386\,
            in1 => \N__43669\,
            in2 => \_gnd_net_\,
            in3 => \N__25341\,
            lcout => OPEN,
            ltout => \ALU.N_224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO0TVG_11_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__19511\,
            in1 => \_gnd_net_\,
            in2 => \N__19457\,
            in3 => \N__39013\,
            lcout => \ALU.N_254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIG4C2T_1_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__23008\,
            in1 => \_gnd_net_\,
            in2 => \N__20819\,
            in3 => \N__38728\,
            lcout => \ALU.N_310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_1_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__42945\,
            in1 => \N__39586\,
            in2 => \N__40433\,
            in3 => \N__39463\,
            lcout => \ALU.madd_484_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINSF07_5_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43665\,
            in1 => \N__40423\,
            in2 => \_gnd_net_\,
            in3 => \N__42946\,
            lcout => \ALU.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIF7TU3_4_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__42947\,
            in1 => \N__23468\,
            in2 => \_gnd_net_\,
            in3 => \N__29426\,
            lcout => \ALU.N_289_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC8LH7_7_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46946\,
            in1 => \N__43666\,
            in2 => \_gnd_net_\,
            in3 => \N__40075\,
            lcout => \ALU.N_220\,
            ltout => \ALU.N_220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIR98G_7_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39014\,
            in2 => \N__19514\,
            in3 => \N__19510\,
            lcout => \ALU.N_252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILPJD8_9_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43664\,
            in1 => \N__39836\,
            in2 => \_gnd_net_\,
            in3 => \N__27603\,
            lcout => \ALU.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_4_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010001000100"
        )
    port map (
            in0 => \N__21488\,
            in1 => \N__46945\,
            in2 => \N__32670\,
            in3 => \N__38324\,
            lcout => \ALU.madd_484_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIDBD49_15_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32661\,
            lcout => \ALU.un9_addsub_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILBFG4_2_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__19487\,
            in1 => \N__29380\,
            in2 => \_gnd_net_\,
            in3 => \N__36980\,
            lcout => \ALU.d_RNILBFG4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m240_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__19639\,
            in1 => \N__19660\,
            in2 => \_gnd_net_\,
            in3 => \N__20290\,
            lcout => \ALU.N_241_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI59DJ3_2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111111"
        )
    port map (
            in0 => \N__20289\,
            in1 => \N__29378\,
            in2 => \N__26577\,
            in3 => \N__28730\,
            lcout => \ALU.N_240_0_i\,
            ltout => \ALU.N_240_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEDJEA_2_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__36979\,
            in1 => \_gnd_net_\,
            in2 => \N__19664\,
            in3 => \N__37201\,
            lcout => \ALU.d_RNIEDJEAZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m10_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__19661\,
            in1 => \N__19640\,
            in2 => \_gnd_net_\,
            in3 => \N__20944\,
            lcout => \ALU.N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_6_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000100010"
        )
    port map (
            in0 => \N__38024\,
            in1 => \N__41722\,
            in2 => \N__33148\,
            in3 => \N__37202\,
            lcout => \ALU.madd_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUV3H4_0_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__19613\,
            in1 => \N__29379\,
            in2 => \_gnd_net_\,
            in3 => \N__38025\,
            lcout => \ALU.d_RNIUV3H4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_0_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38023\,
            in1 => \N__37200\,
            in2 => \N__37002\,
            in3 => \N__38274\,
            lcout => \ALU.madd_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILU4U8_12_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__20895\,
            in1 => \N__37981\,
            in2 => \N__24193\,
            in3 => \N__25452\,
            lcout => \ALU.a0_b_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_rep1_e_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__33355\,
            in1 => \N__19588\,
            in2 => \N__19562\,
            in3 => \N__22294\,
            lcout => \aluReadBus_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47662\,
            ce => \N__34691\,
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_fast_e_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000101"
        )
    port map (
            in0 => \N__22292\,
            in1 => \N__19558\,
            in2 => \N__19589\,
            in3 => \N__33357\,
            lcout => \aluReadBus_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47662\,
            ce => \N__34691\,
            sr => \_gnd_net_\
        );

    \ALU.m246_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001111111"
        )
    port map (
            in0 => \N__30130\,
            in1 => \N__25122\,
            in2 => \N__21859\,
            in3 => \N__29679\,
            lcout => \ALU.N_247_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_e_0_2_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__22291\,
            in1 => \N__19557\,
            in2 => \N__22595\,
            in3 => \N__33358\,
            lcout => \busState_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47662\,
            ce => \N__34691\,
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_e_0_0_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33356\,
            in1 => \N__22293\,
            in2 => \N__22736\,
            in3 => \N__19880\,
            lcout => \busState_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47662\,
            ce => \N__34691\,
            sr => \_gnd_net_\
        );

    \ALU.m210_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111110101"
        )
    port map (
            in0 => \N__29678\,
            in1 => \N__19871\,
            in2 => \N__25165\,
            in3 => \N__30129\,
            lcout => \ALU.N_211_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m204_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001111111"
        )
    port map (
            in0 => \N__30131\,
            in1 => \N__25123\,
            in2 => \N__19757\,
            in3 => \N__29680\,
            lcout => \ALU.N_205_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_367_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19697\,
            in1 => \N__42016\,
            in2 => \N__19718\,
            in3 => \N__39452\,
            lcout => \ALU.madd_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRV558_13_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000100000"
        )
    port map (
            in0 => \N__37429\,
            in1 => \N__25060\,
            in2 => \N__29994\,
            in3 => \N__24999\,
            lcout => \ALU.d_RNIRV558Z0Z_13\,
            ltout => \ALU.d_RNIRV558Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_371_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__19696\,
            in1 => \N__42017\,
            in2 => \N__19709\,
            in3 => \N__39453\,
            lcout => \ALU.madd_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBAHT8_12_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__20915\,
            in1 => \N__36981\,
            in2 => \N__29993\,
            in3 => \N__25453\,
            lcout => \ALU.a2_b_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_259_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010000000"
        )
    port map (
            in0 => \N__19930\,
            in1 => \N__37769\,
            in2 => \N__39383\,
            in3 => \N__19937\,
            lcout => \ALU.madd_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMIK85_11_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__24909\,
            in1 => \N__24134\,
            in2 => \N__31180\,
            in3 => \N__29310\,
            lcout => \ALU.N_186_0\,
            ltout => \ALU.N_186_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3JLT7_1_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19940\,
            in3 => \N__37428\,
            lcout => \ALU.a1_b_11\,
            ltout => \ALU.a1_b_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_255_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__37768\,
            in1 => \N__19931\,
            in2 => \N__19922\,
            in3 => \N__39341\,
            lcout => \ALU.madd_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIU5N11_8_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__31067\,
            in1 => \N__27349\,
            in2 => \N__30974\,
            in3 => \N__27134\,
            lcout => \ALU.dout_3_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIIIOA1_8_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__35989\,
            in1 => \N__47719\,
            in2 => \N__25654\,
            in3 => \N__35899\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI35CK1_8_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__25595\,
            in1 => \N__35366\,
            in2 => \N__19898\,
            in3 => \N__25628\,
            lcout => \ALU.N_755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNITF602_8_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__30908\,
            in1 => \N__35737\,
            in2 => \N__30941\,
            in3 => \N__19895\,
            lcout => OPEN,
            ltout => \ALU.N_707_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI40CO3_8_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35231\,
            in2 => \N__19889\,
            in3 => \N__19886\,
            lcout => \ALU.aluOut_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_26_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__20089\,
            in1 => \N__41501\,
            in2 => \N__41563\,
            in3 => \N__41230\,
            lcout => \ctrlOut_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47678\,
            ce => \N__41055\,
            sr => \_gnd_net_\
        );

    \ALU.m272_ns_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110000000"
        )
    port map (
            in0 => \N__30172\,
            in1 => \N__20087\,
            in2 => \N__26651\,
            in3 => \N__29704\,
            lcout => OPEN,
            ltout => \ALU.m272_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIEUU85_10_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101110111"
        )
    port map (
            in0 => \N__20088\,
            in1 => \N__29367\,
            in2 => \N__20111\,
            in3 => \N__27540\,
            lcout => \ALU.N_273_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g0_7_a3_0_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20082\,
            in2 => \_gnd_net_\,
            in3 => \N__29701\,
            lcout => \ALU.g0_7_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g0_6_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29703\,
            in1 => \N__30021\,
            in2 => \N__20090\,
            in3 => \N__30171\,
            lcout => \ALU.N_191_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m190_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30170\,
            in1 => \N__20083\,
            in2 => \N__24235\,
            in3 => \N__29702\,
            lcout => \ALU.N_191_0\,
            ltout => \ALU.N_191_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBRVD8_10_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__30026\,
            in1 => \N__37391\,
            in2 => \N__20027\,
            in3 => \N__20013\,
            lcout => \ALU.a1_b_10\,
            ltout => \ALU.a1_b_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_203_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__39334\,
            in1 => \N__19954\,
            in2 => \N__19985\,
            in3 => \N__38213\,
            lcout => \ALU.madd_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFO567_9_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39752\,
            in2 => \_gnd_net_\,
            in3 => \N__37145\,
            lcout => \ALU.a9_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI08N11_9_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__38405\,
            in1 => \N__38375\,
            in2 => \N__27353\,
            in3 => \N__27133\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNI1K602_9_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35748\,
            in1 => \N__36131\,
            in2 => \N__19943\,
            in3 => \N__32720\,
            lcout => OPEN,
            ltout => \ALU.N_708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC8CO3_9_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35230\,
            in2 => \N__20171\,
            in3 => \N__20165\,
            lcout => \ALU.aluOut_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIKKOA1_9_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__28160\,
            in1 => \N__28133\,
            in2 => \N__36004\,
            in3 => \N__35897\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI79CK1_9_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35367\,
            in1 => \N__32839\,
            in2 => \N__20168\,
            in3 => \N__32797\,
            lcout => \ALU.N_756\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHBIK1_4_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__27287\,
            in1 => \N__36542\,
            in2 => \N__35754\,
            in3 => \N__28997\,
            lcout => OPEN,
            ltout => \ALU.N_751_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHB2E3_4_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35232\,
            in1 => \_gnd_net_\,
            in2 => \N__20159\,
            in3 => \N__20156\,
            lcout => \ALU.aluOut_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNISKML1_4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__26975\,
            in1 => \N__31862\,
            in2 => \N__35753\,
            in3 => \N__29051\,
            lcout => \ALU.N_703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8MG97_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__43762\,
            in1 => \N__40427\,
            in2 => \N__39139\,
            in3 => \N__42821\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI609EE_6_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__46657\,
            in1 => \N__46837\,
            in2 => \N__20150\,
            in3 => \N__39105\,
            lcout => \ALU.N_472\,
            ltout => \ALU.N_472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6EKGV_6_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38743\,
            in2 => \N__20135\,
            in3 => \N__20132\,
            lcout => \ALU.N_532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_N_1700_i_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38178\,
            lcout => \ALU.N_1700_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNI81NL1_7_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__31814\,
            in1 => \N__31694\,
            in2 => \N__35738\,
            in3 => \N__21599\,
            lcout => OPEN,
            ltout => \ALU.N_706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBDSD3_7_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35220\,
            in2 => \N__20213\,
            in3 => \N__20210\,
            lcout => \ALU.aluOut_7\,
            ltout => \ALU.aluOut_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIE5297_6_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000100000"
        )
    port map (
            in0 => \N__26595\,
            in1 => \N__26280\,
            in2 => \N__20204\,
            in3 => \N__26711\,
            lcout => \ALU.a7_b_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIP6PD3_1_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__25169\,
            in1 => \N__23336\,
            in2 => \_gnd_net_\,
            in3 => \N__23290\,
            lcout => \ALU.N_249_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI64QK7_4_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__23485\,
            in1 => \N__23566\,
            in2 => \N__26626\,
            in3 => \N__37894\,
            lcout => \ALU.a0_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIP0RR6_3_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41926\,
            in2 => \_gnd_net_\,
            in3 => \N__38177\,
            lcout => \ALU.a3_b_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIAE1U4_11_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__24926\,
            in1 => \N__39382\,
            in2 => \N__20186\,
            in3 => \N__29309\,
            lcout => \ALU.N_272_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_89_0_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__38176\,
            in1 => \N__40098\,
            in2 => \N__37156\,
            in3 => \N__46658\,
            lcout => \ALU.madd_89_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_20_0_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__41883\,
            in1 => \N__37098\,
            in2 => \N__38273\,
            in3 => \N__40277\,
            lcout => OPEN,
            ltout => \ALU.madd_20_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_20_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__42823\,
            in1 => \_gnd_net_\,
            in2 => \N__20306\,
            in3 => \N__37627\,
            lcout => \ALU.madd_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC6QK6_5_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40276\,
            in2 => \_gnd_net_\,
            in3 => \N__37094\,
            lcout => \ALU.a5_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m4_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30196\,
            in1 => \N__25215\,
            in2 => \_gnd_net_\,
            in3 => \N__29735\,
            lcout => \ALU.N_5_0\,
            ltout => \ALU.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3GPD3_2_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__25170\,
            in1 => \N__20291\,
            in2 => \N__20252\,
            in3 => \N__28726\,
            lcout => \ALU.N_240_0\,
            ltout => \ALU.N_240_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_24_0_tz_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__42822\,
            in1 => \N__41882\,
            in2 => \N__20249\,
            in3 => \N__37626\,
            lcout => \ALU.madd_24_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_66_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36938\,
            in1 => \N__41704\,
            in2 => \N__42969\,
            in3 => \N__28068\,
            lcout => \ALU.madd_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_8_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__38192\,
            in1 => \N__42916\,
            in2 => \N__37158\,
            in3 => \N__36940\,
            lcout => \ALU.madd_8_0\,
            ltout => \ALU.madd_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_18_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__37656\,
            in1 => \N__20228\,
            in2 => \N__20216\,
            in3 => \N__41973\,
            lcout => \ALU.madd_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_128_0_tz_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__40044\,
            in1 => \N__46839\,
            in2 => \N__37157\,
            in3 => \N__37654\,
            lcout => \ALU.madd_128_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_68_0_tz_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__36939\,
            in1 => \N__41705\,
            in2 => \N__42970\,
            in3 => \N__28069\,
            lcout => \ALU.madd_68_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRALR6_7_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46838\,
            lcout => \ALU.a7_b_0\,
            ltout => \ALU.a7_b_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_59_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__37655\,
            in1 => \N__46638\,
            in2 => \N__20417\,
            in3 => \N__24526\,
            lcout => \ALU.madd_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_5_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011010010"
        )
    port map (
            in0 => \N__40045\,
            in1 => \N__47067\,
            in2 => \N__39852\,
            in3 => \N__46444\,
            lcout => \ALU.madd_484_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_26_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__40046\,
            in1 => \N__46876\,
            in2 => \N__37203\,
            in3 => \N__37657\,
            lcout => \ALU.madd_128_0_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_104_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20573\,
            in1 => \N__20588\,
            in2 => \N__24515\,
            in3 => \N__20594\,
            lcout => \ALU.madd_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_149_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20541\,
            in1 => \N__21948\,
            in2 => \_gnd_net_\,
            in3 => \N__20554\,
            lcout => \ALU.madd_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_128_0_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__38272\,
            in1 => \N__39825\,
            in2 => \_gnd_net_\,
            in3 => \N__20336\,
            lcout => \ALU.madd_128_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_m3_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__20543\,
            in1 => \N__21950\,
            in2 => \_gnd_net_\,
            in3 => \N__20555\,
            lcout => \ALU.madd_N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_68_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__41993\,
            in1 => \N__20606\,
            in2 => \N__42698\,
            in3 => \N__20600\,
            lcout => \ALU.madd_68\,
            ltout => \ALU.madd_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_108_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011101000"
        )
    port map (
            in0 => \N__20587\,
            in1 => \N__24511\,
            in2 => \N__20576\,
            in3 => \N__20572\,
            lcout => \ALU.madd_108\,
            ltout => \ALU.madd_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_153_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__21949\,
            in1 => \_gnd_net_\,
            in2 => \N__20546\,
            in3 => \N__20542\,
            lcout => \ALU.madd_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXready_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__24767\,
            in1 => \N__20668\,
            in2 => \N__24661\,
            in3 => \N__24742\,
            lcout => \RXready\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXreadyC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_RNI29TH_2_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29249\,
            in2 => \_gnd_net_\,
            in3 => \N__24652\,
            lcout => \FTDI.N_201_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_2_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010100000"
        )
    port map (
            in0 => \N__24768\,
            in1 => \N__20669\,
            in2 => \N__24662\,
            in3 => \N__24743\,
            lcout => \FTDI.RXstateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXreadyC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m681_1_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43090\,
            in1 => \N__20479\,
            in2 => \N__48054\,
            in3 => \N__44028\,
            lcout => OPEN,
            ltout => \ALU.m681Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m681_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__33173\,
            in1 => \N__45699\,
            in2 => \N__20462\,
            in3 => \N__26649\,
            lcout => \ALU.N_730_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m57_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30285\,
            in2 => \_gnd_net_\,
            in3 => \N__21883\,
            lcout => \ALU.N_58_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNI67DS1_0_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24766\,
            in1 => \N__24741\,
            in2 => \N__24660\,
            in3 => \N__24688\,
            lcout => \FTDI.gap8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNIV5TH_0_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29250\,
            lcout => \FTDI.N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEN0V7_0_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011010"
        )
    port map (
            in0 => \N__38306\,
            in1 => \_gnd_net_\,
            in2 => \N__38045\,
            in3 => \N__43859\,
            lcout => \ALU.a_15_m1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID9RV5_0_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__44037\,
            in1 => \N__47230\,
            in2 => \N__44524\,
            in3 => \N__20755\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINPK3M_0_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__44159\,
            in1 => \N__20660\,
            in2 => \N__20654\,
            in3 => \N__20624\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITQOAQ2_0_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46310\,
            in2 => \N__20651\,
            in3 => \N__20648\,
            lcout => \ALU.a_15_m5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m4_bm_1_8_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__47229\,
            in1 => \_gnd_net_\,
            in2 => \N__43881\,
            in3 => \N__24579\,
            lcout => \ALU.a_15_m4_bm_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITTVL7_0_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__24580\,
            in1 => \N__38022\,
            in2 => \_gnd_net_\,
            in3 => \N__38307\,
            lcout => \ALU.a_15_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_0_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__22137\,
            in1 => \N__20618\,
            in2 => \_gnd_net_\,
            in3 => \N__43583\,
            lcout => \aluParams_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPD997_6_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__43582\,
            in1 => \N__40424\,
            in2 => \N__38968\,
            in3 => \N__46734\,
            lcout => \ALU.rshift_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI5PUHV_10_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000111011"
        )
    port map (
            in0 => \N__20702\,
            in1 => \N__43139\,
            in2 => \N__44449\,
            in3 => \N__20735\,
            lcout => \ALU.a_15_m3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFL4K8_11_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43674\,
            in1 => \N__39385\,
            in2 => \_gnd_net_\,
            in3 => \N__27589\,
            lcout => \ALU.N_461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3BB3U_5_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38559\,
            in1 => \N__24818\,
            in2 => \_gnd_net_\,
            in3 => \N__20714\,
            lcout => OPEN,
            ltout => \ALU.N_530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIP8ITN1_5_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44393\,
            in2 => \N__20705\,
            in3 => \N__20701\,
            lcout => OPEN,
            ltout => \ALU.d_RNIP8ITN1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFHQSS1_2_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43140\,
            in2 => \N__20693\,
            in3 => \N__20690\,
            lcout => OPEN,
            ltout => \ALU.a_15_m3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDVDOJ2_2_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46311\,
            in2 => \N__20681\,
            in3 => \N__20675\,
            lcout => \ALU.a_15_m5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIE937B_0_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__38560\,
            in1 => \N__44422\,
            in2 => \_gnd_net_\,
            in3 => \N__39180\,
            lcout => OPEN,
            ltout => \ALU.d_RNIE937BZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVM1UL_2_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44139\,
            in2 => \N__20678\,
            in3 => \N__24830\,
            lcout => \ALU.a_15_m4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI75NNF_6_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__38966\,
            in1 => \N__22915\,
            in2 => \N__38603\,
            in3 => \N__22894\,
            lcout => \ALU.lshift_7_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINVVJ11_13_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__38593\,
            in1 => \N__20777\,
            in2 => \N__44492\,
            in3 => \N__20767\,
            lcout => \ALU.lshift_15_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNII1LGE_5_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38967\,
            in1 => \N__22810\,
            in2 => \_gnd_net_\,
            in3 => \N__22895\,
            lcout => \ALU.N_249\,
            ltout => \ALU.N_249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIUGCLV_11_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38528\,
            in2 => \N__20771\,
            in3 => \N__20768\,
            lcout => OPEN,
            ltout => \ALU.c_RNIUGCLVZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILTHAE1_1_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44443\,
            in2 => \N__20759\,
            in3 => \N__22823\,
            lcout => \ALU.lshift_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEUKR11_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44442\,
            in1 => \N__20756\,
            in2 => \_gnd_net_\,
            in3 => \N__20744\,
            lcout => \ALU.d_RNIEUKR11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI83IG7_3_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__43620\,
            in1 => \N__41995\,
            in2 => \N__42997\,
            in3 => \N__39141\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICH0SD_1_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__36957\,
            in1 => \N__38965\,
            in2 => \N__20738\,
            in3 => \N__37426\,
            lcout => \ALU.N_246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFL4K8_0_11_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27558\,
            in1 => \N__43586\,
            in2 => \_gnd_net_\,
            in3 => \N__39389\,
            lcout => \ALU.N_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5MUQE_6_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39142\,
            in1 => \N__20825\,
            in2 => \_gnd_net_\,
            in3 => \N__20801\,
            lcout => \ALU.N_250\,
            ltout => \ALU.N_250_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNISJ8601_11_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__38722\,
            in1 => \_gnd_net_\,
            in2 => \N__20810\,
            in3 => \N__20807\,
            lcout => \ALU.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVUE24_0_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__43587\,
            in1 => \N__39144\,
            in2 => \_gnd_net_\,
            in3 => \N__37962\,
            lcout => \ALU.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIK8CGE_5_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39145\,
            in1 => \N__22803\,
            in2 => \_gnd_net_\,
            in3 => \N__23043\,
            lcout => \ALU.N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8K807_6_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43585\,
            in1 => \N__40402\,
            in2 => \_gnd_net_\,
            in3 => \N__46720\,
            lcout => \ALU.N_218\,
            ltout => \ALU.N_218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGNQGE_3_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39143\,
            in2 => \N__20795\,
            in3 => \N__23024\,
            lcout => \ALU.N_361\,
            ltout => \ALU.N_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1GH4V_7_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38723\,
            in2 => \N__20792\,
            in3 => \N__20788\,
            lcout => \ALU.d_RNI1GH4VZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_28_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__32293\,
            in1 => \N__41159\,
            in2 => \N__20972\,
            in3 => \N__41474\,
            lcout => \ctrlOut_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47650\,
            ce => \N__41060\,
            sr => \_gnd_net_\
        );

    \ALU.m270_ns_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110000000"
        )
    port map (
            in0 => \N__30193\,
            in1 => \N__26637\,
            in2 => \N__20971\,
            in3 => \N__29692\,
            lcout => OPEN,
            ltout => \ALU.m270_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNILQ2U4_12_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__25348\,
            in1 => \N__20966\,
            in2 => \N__20975\,
            in3 => \N__29403\,
            lcout => \ALU.N_271_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m178_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30192\,
            in1 => \N__25139\,
            in2 => \N__20970\,
            in3 => \N__29691\,
            lcout => \ALU.N_179_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIM75G5_15_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__24149\,
            in1 => \N__29402\,
            in2 => \N__20945\,
            in3 => \N__31322\,
            lcout => \ALU.N_7_0\,
            ltout => \ALU.N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_0_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__41976\,
            in1 => \N__37961\,
            in2 => \N__20921\,
            in3 => \N__40826\,
            lcout => \ALU.madd_484_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4K3G5_12_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24148\,
            in1 => \N__20894\,
            in2 => \_gnd_net_\,
            in3 => \N__25442\,
            lcout => \ALU.N_180_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_13_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47233\,
            in1 => \N__24588\,
            in2 => \_gnd_net_\,
            in3 => \N__43861\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNID22SC_13_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010100101011"
        )
    port map (
            in0 => \N__40746\,
            in1 => \N__24969\,
            in2 => \N__20873\,
            in3 => \N__47234\,
            lcout => \ALU.a_15_m2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m714_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44133\,
            in2 => \_gnd_net_\,
            in3 => \N__43584\,
            lcout => \ALU.log_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_3_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010001000100"
        )
    port map (
            in0 => \N__22002\,
            in1 => \N__46729\,
            in2 => \N__40764\,
            in3 => \N__37231\,
            lcout => \ALU.madd_484_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIG6C84_9_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__32990\,
            in1 => \N__28109\,
            in2 => \N__24449\,
            in3 => \N__32849\,
            lcout => \ALU.operand2_9\,
            ltout => \ALU.operand2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHIKU4_9_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21057\,
            in2 => \N__21032\,
            in3 => \N__24144\,
            lcout => \ALU.N_207_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_9_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__47231\,
            in1 => \N__24587\,
            in2 => \_gnd_net_\,
            in3 => \N__43860\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6904C_9_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101001101"
        )
    port map (
            in0 => \N__22003\,
            in1 => \N__47232\,
            in2 => \N__21029\,
            in3 => \N__39832\,
            lcout => \ALU.a_15_m2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_13_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48598\,
            in1 => \N__33940\,
            in2 => \N__45873\,
            in3 => \N__33881\,
            lcout => \ALU.hZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47663\,
            ce => \N__45489\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO7LU_13_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45334\,
            in1 => \N__35446\,
            in2 => \_gnd_net_\,
            in3 => \N__35435\,
            lcout => OPEN,
            ltout => \ALU.d_RNIO7LUZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8DRP4_0_13_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__28439\,
            in1 => \N__32994\,
            in2 => \N__21026\,
            in3 => \N__31103\,
            lcout => \ALU.operand2_13\,
            ltout => \ALU.operand2_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDT3G5_13_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__25053\,
            in1 => \_gnd_net_\,
            in2 => \N__21023\,
            in3 => \N__24153\,
            lcout => \ALU.N_177_0\,
            ltout => \ALU.N_177_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_2_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010100110"
        )
    port map (
            in0 => \N__37376\,
            in1 => \N__36878\,
            in2 => \N__21020\,
            in3 => \N__21313\,
            lcout => OPEN,
            ltout => \ALU.madd_484_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_12_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21017\,
            in1 => \N__21008\,
            in2 => \N__20996\,
            in3 => \N__20993\,
            lcout => \ALU.madd_484_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7TLM8_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__39440\,
            in1 => \N__37968\,
            in2 => \N__36325\,
            in3 => \_gnd_net_\,
            lcout => \ALU.a0_b_11\,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \ALU.un2_addsub_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_0_c_RNI5MA0E_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23351\,
            in2 => \N__23279\,
            in3 => \N__21215\,
            lcout => \ALU.un2_addsub_cry_0_c_RNI5MA0EZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_0\,
            carryout => \ALU.un2_addsub_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_1_c_RNI966GE_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21212\,
            in2 => \N__21197\,
            in3 => \N__21179\,
            lcout => \ALU.un2_addsub_cry_1_c_RNI966GEZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_1\,
            carryout => \ALU.un2_addsub_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_2_c_RNI5IV5F_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41719\,
            in2 => \N__23846\,
            in3 => \N__21176\,
            lcout => \ALU.un2_addsub_cry_2_c_RNI5IV5FZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_2\,
            carryout => \ALU.un2_addsub_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_3_c_RNIOGGJG_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42683\,
            in2 => \N__21800\,
            in3 => \N__21173\,
            lcout => \ALU.un2_addsub_cry_3_c_RNIOGGJGZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_3\,
            carryout => \ALU.un2_addsub_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_4_c_RNI284VE_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28090\,
            in2 => \N__21170\,
            in3 => \N__21152\,
            lcout => \ALU.un2_addsub_cry_4_c_RNI284VEZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_4\,
            carryout => \ALU.un2_addsub_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_5_c_RNIL7IGF_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46474\,
            in2 => \N__21149\,
            in3 => \N__21128\,
            lcout => \ALU.un2_addsub_cry_5_c_RNIL7IGFZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_5\,
            carryout => \ALU.un2_addsub_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_6_c_RNIL4LMI_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47101\,
            in2 => \N__21125\,
            in3 => \N__21101\,
            lcout => \ALU.un2_addsub_cry_6_c_RNIL4LMIZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_6\,
            carryout => \ALU.un2_addsub_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_7_c_RNIL8JHG_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21471\,
            in2 => \N__21404\,
            in3 => \N__21386\,
            lcout => \ALU.un2_addsub_cry_7_c_RNIL8JHGZ0\,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \ALU.un2_addsub_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_8_c_RNIKR81J_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22057\,
            in2 => \N__21383\,
            in3 => \N__21368\,
            lcout => \ALU.un2_addsub_cry_8_c_RNIKR81JZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_8\,
            carryout => \ALU.un2_addsub_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_9_c_RNIVCOFA_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27511\,
            in2 => \N__21365\,
            in3 => \N__21347\,
            lcout => \ALU.un2_addsub_cry_9_c_RNIVCOFAZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_9\,
            carryout => \ALU.un2_addsub_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_10_c_RNIUS1OJ_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25571\,
            in2 => \N__24848\,
            in3 => \N__21344\,
            lcout => \ALU.un2_addsub_cry_10_c_RNIUS1OJZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_10\,
            carryout => \ALU.un2_addsub_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_11_c_RNII7OF9_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25379\,
            in2 => \N__21341\,
            in3 => \N__21320\,
            lcout => \ALU.un2_addsub_cry_11_c_RNII7OFZ0Z9\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_11\,
            carryout => \ALU.un2_addsub_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_12_c_RNIUL1GK_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24973\,
            in2 => \N__24947\,
            in3 => \N__21317\,
            lcout => \ALU.un2_addsub_cry_12_c_RNIUL1GKZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_12\,
            carryout => \ALU.un2_addsub_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_13_c_RNINVE5K_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21314\,
            in2 => \N__21263\,
            in3 => \N__21245\,
            lcout => \ALU.un2_addsub_cry_13_c_RNINVE5KZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_13\,
            carryout => \ALU.un2_addsub_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_14_c_RNINOK69_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32608\,
            in1 => \N__32675\,
            in2 => \_gnd_net_\,
            in3 => \N__21242\,
            lcout => \ALU.un2_addsub_cry_14_c_RNINOKZ0Z69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_10_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111010001"
        )
    port map (
            in0 => \N__34326\,
            in1 => \N__45842\,
            in2 => \N__34415\,
            in3 => \N__48251\,
            lcout => \ALU.hZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47679\,
            ce => \N__45586\,
            sr => \_gnd_net_\
        );

    \ALU.g0_2_1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111011101"
        )
    port map (
            in0 => \N__31260\,
            in1 => \N__25213\,
            in2 => \N__30216\,
            in3 => \N__21518\,
            lcout => \ALU.g0_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIPN2P1_10_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111010"
        )
    port map (
            in0 => \N__28600\,
            in1 => \N__23707\,
            in2 => \N__34514\,
            in3 => \N__34814\,
            lcout => OPEN,
            ltout => \ALU.N_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIULHV4_10_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__25214\,
            in1 => \N__21500\,
            in2 => \N__21512\,
            in3 => \N__21509\,
            lcout => \ALU.N_192_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGNUR_10_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001110111"
        )
    port map (
            in0 => \N__28422\,
            in1 => \N__35026\,
            in2 => \N__24427\,
            in3 => \N__34901\,
            lcout => OPEN,
            ltout => \ALU.g0_7_m4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIT7R92_10_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001010"
        )
    port map (
            in0 => \N__26827\,
            in1 => \N__28525\,
            in2 => \N__21503\,
            in3 => \N__34508\,
            lcout => \ALU.N_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNITA7N_0_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__28933\,
            in1 => \N__27124\,
            in2 => \N__27040\,
            in3 => \N__28952\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIC4ML1_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35707\,
            in1 => \N__31943\,
            in2 => \N__21494\,
            in3 => \N__29138\,
            lcout => \ALU.N_699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIGRS31_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__27126\,
            in1 => \N__27325\,
            in2 => \N__36299\,
            in3 => \N__35051\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1RHK1_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35708\,
            in1 => \N__21536\,
            in2 => \N__21491\,
            in3 => \N__42194\,
            lcout => \ALU.N_747\,
            ltout => \ALU.N_747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHA1E3_0_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35206\,
            in1 => \_gnd_net_\,
            in2 => \N__21623\,
            in3 => \N__27256\,
            lcout => \ALU.aluOut_0\,
            ltout => \ALU.aluOut_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_N_2L1_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__39531\,
            in1 => \_gnd_net_\,
            in2 => \N__21620\,
            in3 => \_gnd_net_\,
            lcout => \ALU.g0_0_0_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIBP7N_7_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__28798\,
            in1 => \N__27870\,
            in2 => \N__27041\,
            in3 => \N__27125\,
            lcout => \ALU.dout_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9BO713_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__37933\,
            in1 => \N__46041\,
            in2 => \N__21593\,
            in3 => \N__38190\,
            lcout => \ALU.d_RNI9BO713Z0Z_0\,
            ltout => \ALU.d_RNI9BO713Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48433\,
            in2 => \N__21581\,
            in3 => \N__42326\,
            lcout => \ALU.hZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47687\,
            ce => \N__45587\,
            sr => \_gnd_net_\
        );

    \ALU.e_RNIHCSL1_0_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__31041\,
            in1 => \N__31597\,
            in2 => \N__28904\,
            in3 => \N__28850\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPDJU2_0_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31262\,
            in1 => \N__21524\,
            in2 => \N__21578\,
            in3 => \N__31607\,
            lcout => OPEN,
            ltout => \ALU.operand2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGTOD3_0_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21575\,
            in1 => \N__29292\,
            in2 => \N__21539\,
            in3 => \N__25220\,
            lcout => \ALU.N_252_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIE4R7_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21535\,
            in1 => \N__42193\,
            in2 => \_gnd_net_\,
            in3 => \N__32068\,
            lcout => \ALU.d_RNIE4R7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIT0CO_1_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34884\,
            in2 => \N__31922\,
            in3 => \N__29117\,
            lcout => OPEN,
            ltout => \ALU.g_RNIT0COZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNILGSL1_1_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__31046\,
            in1 => \N__31598\,
            in2 => \N__21659\,
            in3 => \N__21653\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1MJU2_1_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__31265\,
            in1 => \N__28838\,
            in2 => \N__21656\,
            in3 => \N__31709\,
            lcout => \ALU.operand2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIPKVJ_1_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34883\,
            in1 => \N__44596\,
            in2 => \_gnd_net_\,
            in3 => \N__26933\,
            lcout => \ALU.e_RNIPKVJZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_11_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41863\,
            in1 => \N__37118\,
            in2 => \N__36945\,
            in3 => \N__37647\,
            lcout => \ALU.madd_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMH5R6_2_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36861\,
            in2 => \_gnd_net_\,
            in3 => \N__38179\,
            lcout => \ALU.a2_b_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_12_0_tz_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__41862\,
            in1 => \N__37117\,
            in2 => \N__36944\,
            in3 => \N__37646\,
            lcout => \ALU.madd_12_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIVFBD1_15_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__28496\,
            in1 => \N__35699\,
            in2 => \N__25916\,
            in3 => \N__35576\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC5K02_15_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__33476\,
            in1 => \N__35376\,
            in2 => \N__21626\,
            in3 => \N__33500\,
            lcout => \ALU.N_762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_1_rep2_e_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26881\,
            lcout => \aluOperand1_1_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47689\,
            ce => \N__27727\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5IGD1_5_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__31406\,
            in1 => \N__43400\,
            in2 => \N__35384\,
            in3 => \N__23663\,
            lcout => OPEN,
            ltout => \ALU.N_752_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9M073_5_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35183\,
            in2 => \N__21815\,
            in3 => \N__21809\,
            lcout => \ALU.aluOut_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_fast_e_1_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aluOperand1_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47689\,
            ce => \N__27727\,
            sr => \_gnd_net_\
        );

    \ALU.e_RNI7L7N_5_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__27108\,
            in1 => \N__44641\,
            in2 => \N__27039\,
            in3 => \N__28868\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNI0PML1_5_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35698\,
            in1 => \N__31835\,
            in2 => \N__21812\,
            in3 => \N__29030\,
            lcout => \ALU.N_704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI65RK7_4_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101001011001"
        )
    port map (
            in0 => \N__42904\,
            in1 => \N__26605\,
            in2 => \N__23500\,
            in3 => \N__23559\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI312TB_4_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21803\,
            in3 => \N__42696\,
            lcout => \ALU.d_RNI312TBZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITKRB7_5_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__21788\,
            in1 => \N__41864\,
            in2 => \N__24340\,
            in3 => \N__21724\,
            lcout => \ALU.a3_b_5\,
            ltout => \ALU.a3_b_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_94_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__40292\,
            in1 => \N__22100\,
            in2 => \N__21674\,
            in3 => \N__41695\,
            lcout => \ALU.madd_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIE79M7_4_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__23558\,
            in1 => \N__23493\,
            in2 => \N__24341\,
            in3 => \N__42903\,
            lcout => \ALU.a4_b_4\,
            ltout => \ALU.a4_b_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_98_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101000"
        )
    port map (
            in0 => \N__40291\,
            in1 => \N__22094\,
            in2 => \N__22088\,
            in3 => \N__41694\,
            lcout => \ALU.madd_98\,
            ltout => \ALU.madd_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_139_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__22068\,
            in1 => \N__38034\,
            in2 => \N__21980\,
            in3 => \N__21973\,
            lcout => \ALU.madd_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNO_0_3_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001101"
        )
    port map (
            in0 => \N__24740\,
            in1 => \N__24659\,
            in2 => \N__21934\,
            in3 => \N__24772\,
            lcout => \FTDI.m13_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_1_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001111100000"
        )
    port map (
            in0 => \N__21888\,
            in1 => \N__30805\,
            in2 => \N__30302\,
            in3 => \N__41293\,
            lcout => \testStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001101011100"
        )
    port map (
            in0 => \N__41292\,
            in1 => \N__21887\,
            in2 => \N__30809\,
            in3 => \N__30289\,
            lcout => \testStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m40_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010001"
        )
    port map (
            in0 => \N__22581\,
            in1 => \N__22723\,
            in2 => \N__21860\,
            in3 => \N__22436\,
            lcout => OPEN,
            ltout => \ALU.N_41_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_e_0_1_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111000000"
        )
    port map (
            in0 => \N__22437\,
            in1 => \N__33331\,
            in2 => \N__21824\,
            in3 => \N__22742\,
            lcout => \aluParams_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47618\,
            ce => \N__22139\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPKIOE_7_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__21821\,
            in1 => \N__40111\,
            in2 => \N__38972\,
            in3 => \N__46974\,
            lcout => \ALU.N_473\,
            ltout => \ALU.N_473_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4HG101_7_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38540\,
            in2 => \N__22745\,
            in3 => \N__31767\,
            lcout => \ALU.d_RNI4HG101Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m42_ns_1_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101001100"
        )
    port map (
            in0 => \N__22297\,
            in1 => \N__38888\,
            in2 => \N__22598\,
            in3 => \N__33330\,
            lcout => \ALU.m42_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINEO9E_1_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__38887\,
            in1 => \N__23144\,
            in2 => \N__38678\,
            in3 => \N__23054\,
            lcout => \ALU.lshift_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m286_am_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011010000010"
        )
    port map (
            in0 => \N__22295\,
            in1 => \N__22432\,
            in2 => \N__22597\,
            in3 => \N__22721\,
            lcout => \ALU.m286_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m286_bm_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22722\,
            in1 => \N__22574\,
            in2 => \N__22442\,
            in3 => \N__22296\,
            lcout => \ALU.m286_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICH0SD_3_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__22829\,
            in1 => \N__42015\,
            in2 => \N__38971\,
            in3 => \N__42996\,
            lcout => OPEN,
            ltout => \ALU.N_469_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI41DBT_3_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__44420\,
            in1 => \N__38591\,
            in2 => \N__22166\,
            in3 => \N__22163\,
            lcout => OPEN,
            ltout => \ALU.rshift_15_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO3KRQ1_15_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__44421\,
            in1 => \N__31790\,
            in2 => \N__22157\,
            in3 => \N__31771\,
            lcout => \ALU.rshift_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_2_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__22154\,
            in1 => \N__22138\,
            in2 => \_gnd_net_\,
            in3 => \N__38592\,
            lcout => \aluParams_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6JKM8_9_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__43621\,
            in1 => \N__39855\,
            in2 => \N__38969\,
            in3 => \N__27588\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNICVGTG_11_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__39012\,
            in1 => \N__39286\,
            in2 => \N__22832\,
            in3 => \N__25370\,
            lcout => \ALU.N_477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI19RM6_1_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__43622\,
            in1 => \N__36993\,
            in2 => \N__38970\,
            in3 => \N__37427\,
            lcout => \ALU.rshift_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINEO9E_0_1_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__23053\,
            in1 => \N__39029\,
            in2 => \N__38677\,
            in3 => \N__23143\,
            lcout => \ALU.d_RNINEO9E_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJ1PCQ_1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__44149\,
            in1 => \N__23639\,
            in2 => \N__44521\,
            in3 => \N__22841\,
            lcout => \ALU.d_RNIJ1PCQZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9HFAU_5_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__23052\,
            in1 => \N__22814\,
            in2 => \N__38676\,
            in3 => \N__22787\,
            lcout => OPEN,
            ltout => \ALU.N_311_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKBPO51_5_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44438\,
            in2 => \N__22781\,
            in3 => \N__22840\,
            lcout => OPEN,
            ltout => \ALU.lshift_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPFIBI1_9_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44148\,
            in2 => \N__22778\,
            in3 => \N__22775\,
            lcout => \ALU.d_RNIPFIBI1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA28GU1_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43149\,
            in1 => \N__22763\,
            in2 => \_gnd_net_\,
            in3 => \N__22751\,
            lcout => OPEN,
            ltout => \ALU.d_RNIA28GU1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISQIQP2_1_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46326\,
            in1 => \_gnd_net_\,
            in2 => \N__22955\,
            in3 => \N__22952\,
            lcout => \ALU.a_15_m5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI2CSHH_13_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__39150\,
            in1 => \N__22946\,
            in2 => \N__38727\,
            in3 => \N__22933\,
            lcout => OPEN,
            ltout => \ALU.lshift_7_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIONI011_6_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__38689\,
            in1 => \N__22919\,
            in2 => \N__22898\,
            in3 => \N__22893\,
            lcout => OPEN,
            ltout => \ALU.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINQ8VM1_6_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__44487\,
            in1 => \_gnd_net_\,
            in2 => \N__22871\,
            in3 => \N__27958\,
            lcout => OPEN,
            ltout => \ALU.lshift_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3O3A42_13_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__44150\,
            in1 => \_gnd_net_\,
            in2 => \N__22868\,
            in3 => \N__22865\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI88B4N2_13_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__46330\,
            in1 => \_gnd_net_\,
            in2 => \N__22856\,
            in3 => \N__24791\,
            lcout => \c_RNI88B4N2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIV49JL_1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__39037\,
            in1 => \N__23142\,
            in2 => \N__38729\,
            in3 => \N__22853\,
            lcout => \ALU.N_420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1HDEU1_13_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__23089\,
            in2 => \N__44522\,
            in3 => \N__22847\,
            lcout => \ALU.lshift_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBSS27_1_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__38685\,
            in1 => \N__39149\,
            in2 => \_gnd_net_\,
            in3 => \N__23141\,
            lcout => \ALU.N_416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICIR67_3_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43714\,
            in1 => \N__36953\,
            in2 => \_gnd_net_\,
            in3 => \N__41977\,
            lcout => \ALU.N_377\,
            ltout => \ALU.N_377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIOHBUD_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39147\,
            in2 => \N__23027\,
            in3 => \N__23137\,
            lcout => \ALU.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN9H77_3_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43715\,
            in1 => \N__41978\,
            in2 => \_gnd_net_\,
            in3 => \N__42980\,
            lcout => \ALU.N_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIADS9I_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38724\,
            in1 => \N__23018\,
            in2 => \_gnd_net_\,
            in3 => \N__23012\,
            lcout => \ALU.N_419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGFQD6_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43713\,
            in1 => \N__36952\,
            in2 => \_gnd_net_\,
            in3 => \N__37419\,
            lcout => \ALU.N_376\,
            ltout => \ALU.N_376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEBMRA_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__38725\,
            in1 => \N__39148\,
            in2 => \N__22997\,
            in3 => \N__27245\,
            lcout => OPEN,
            ltout => \ALU.d_RNIEBMRAZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFPKBA1_0_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44444\,
            in2 => \N__22994\,
            in3 => \N__22991\,
            lcout => \ALU.lshift_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICGVRD_3_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__41979\,
            in1 => \N__39146\,
            in2 => \N__36997\,
            in3 => \N__23111\,
            lcout => \ALU.N_468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIG5BH6_3_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23917\,
            in1 => \N__37371\,
            in2 => \N__26598\,
            in3 => \N__24014\,
            lcout => \ALU.a1_b_3\,
            ltout => \ALU.a1_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_13_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__23219\,
            in1 => \N__23158\,
            in2 => \N__23192\,
            in3 => \N__23189\,
            lcout => \ALU.madd_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKFBA7_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000000000"
        )
    port map (
            in0 => \N__23918\,
            in1 => \N__24013\,
            in2 => \N__26599\,
            in3 => \N__37994\,
            lcout => \ALU.a0_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIR5FE6_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__37995\,
            in1 => \_gnd_net_\,
            in2 => \N__37425\,
            in3 => \N__43684\,
            lcout => \ALU.N_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILPO64_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__23456\,
            in1 => \_gnd_net_\,
            in2 => \N__26600\,
            in3 => \N__23568\,
            lcout => \ALU.N_231_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI35AS3_3_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__24015\,
            in1 => \N__26549\,
            in2 => \_gnd_net_\,
            in3 => \N__23919\,
            lcout => \ALU.N_237_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICVFN6_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__43683\,
            in1 => \N__37372\,
            in2 => \N__39140\,
            in3 => \N__37996\,
            lcout => \ALU.rshift_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9GDQS_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38726\,
            in1 => \N__23105\,
            in2 => \_gnd_net_\,
            in3 => \N__23090\,
            lcout => \ALU.N_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI1FPGN1_10_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23078\,
            in1 => \_gnd_net_\,
            in2 => \N__44218\,
            in3 => \N__23258\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI5V90O2_10_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23069\,
            in2 => \N__23057\,
            in3 => \N__46382\,
            lcout => \c_RNI5V90O2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIJQBMC_10_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111010100"
        )
    port map (
            in0 => \N__23252\,
            in1 => \N__27550\,
            in2 => \N__39606\,
            in3 => \N__47279\,
            lcout => \ALU.a_15_m2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_10_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__47278\,
            in1 => \N__44188\,
            in2 => \N__43938\,
            in3 => \N__43729\,
            lcout => \ALU.a_15_m2_ns_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_9_c_RNI8H83V_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__42522\,
            in1 => \N__39488\,
            in2 => \_gnd_net_\,
            in3 => \N__23246\,
            lcout => OPEN,
            ltout => \un9_addsub_cry_9_c_RNI8H83V_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNINNN4N3_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48329\,
            in2 => \N__23237\,
            in3 => \N__23234\,
            lcout => \aluOperation_RNINNN4N3_0\,
            ltout => \aluOperation_RNINNN4N3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_10_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48330\,
            in1 => \N__45967\,
            in2 => \N__23228\,
            in3 => \N__34411\,
            lcout => \ALU.aZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47656\,
            ce => \N__44837\,
            sr => \_gnd_net_\
        );

    \ALU.b_RNIM5AD1_11_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__35906\,
            in1 => \N__28475\,
            in2 => \N__35582\,
            in3 => \N__28457\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRII02_11_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__31136\,
            in1 => \N__35374\,
            in2 => \N__23225\,
            in3 => \N__31157\,
            lcout => \ALU.N_758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI41LF1_11_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__30830\,
            in1 => \N__35996\,
            in2 => \N__35911\,
            in3 => \N__32489\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI76HQ1_11_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__34112\,
            in1 => \N__35375\,
            in2 => \N__23222\,
            in3 => \N__31307\,
            lcout => OPEN,
            ltout => \ALU.N_710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI64TU3_11_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23378\,
            in2 => \N__23372\,
            in3 => \N__35222\,
            lcout => \ALU.aluOut_11\,
            ltout => \ALU.aluOut_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_484_6_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011010010"
        )
    port map (
            in0 => \N__27499\,
            in1 => \N__28089\,
            in2 => \N__23369\,
            in3 => \N__42644\,
            lcout => \ALU.madd_484_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJM067_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__37348\,
            in1 => \N__43933\,
            in2 => \_gnd_net_\,
            in3 => \N__37716\,
            lcout => \ALU.d_RNIJM067Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI80E86_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001100011"
        )
    port map (
            in0 => \N__23338\,
            in1 => \N__37347\,
            in2 => \N__26642\,
            in3 => \N__23300\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC4AT9_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23354\,
            in3 => \N__23278\,
            lcout => \ALU.d_RNIC4AT9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI5NDI1_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__27377\,
            in1 => \N__35224\,
            in2 => \N__35385\,
            in3 => \N__26945\,
            lcout => OPEN,
            ltout => \ALU.dout_7_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID01L2_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__28826\,
            in1 => \N__35225\,
            in2 => \N__23345\,
            in3 => \N__31724\,
            lcout => \ALU.aluOut_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI44SK3_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__30049\,
            in1 => \N__23337\,
            in2 => \_gnd_net_\,
            in3 => \N__23299\,
            lcout => \ALU.N_249_0\,
            ltout => \ALU.N_249_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI61SHA_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010001100"
        )
    port map (
            in0 => \N__37349\,
            in1 => \N__24594\,
            in2 => \N__23261\,
            in3 => \N__37717\,
            lcout => OPEN,
            ltout => \ALU.d_RNI61SHAZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9CMFI_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47277\,
            in2 => \N__23648\,
            in3 => \N__23645\,
            lcout => \ALU.a_15_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIK6LL_4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32081\,
            in1 => \N__31861\,
            in2 => \_gnd_net_\,
            in3 => \N__29047\,
            lcout => OPEN,
            ltout => \ALU.g_RNIK6LLZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI5F2S1_4_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__31261\,
            in1 => \N__35027\,
            in2 => \N__23627\,
            in3 => \N__23624\,
            lcout => \ALU.operand2_7_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIGQ8H_4_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32080\,
            in1 => \N__27941\,
            in2 => \_gnd_net_\,
            in3 => \N__26963\,
            lcout => \ALU.e_RNIGQ8HZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAS7T6_4_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23487\,
            in1 => \N__37318\,
            in2 => \N__24290\,
            in3 => \N__23523\,
            lcout => \ALU.a1_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3GJL7_4_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__23524\,
            in1 => \N__24253\,
            in2 => \N__23489\,
            in3 => \N__36813\,
            lcout => \ALU.a2_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1LUH3_4_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__24389\,
            in1 => \N__45389\,
            in2 => \N__33104\,
            in3 => \N__23579\,
            lcout => \ALU.operand2_4\,
            ltout => \ALU.operand2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITR684_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23488\,
            in2 => \N__23396\,
            in3 => \N__24249\,
            lcout => \ALU.N_231_0\,
            ltout => \ALU.N_231_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_168_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__39751\,
            in1 => \N__46648\,
            in2 => \N__23393\,
            in3 => \N__37715\,
            lcout => \ALU.madd_93_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIGOP81_10_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__28593\,
            in1 => \N__23706\,
            in2 => \N__27337\,
            in3 => \N__27129\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1PNQ1_10_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35709\,
            in1 => \N__34283\,
            in2 => \N__23678\,
            in3 => \N__34933\,
            lcout => \ALU.N_709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI471O1_10_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__26828\,
            in1 => \N__28526\,
            in2 => \N__35985\,
            in3 => \N__35876\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7I9B2_10_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__28426\,
            in1 => \N__35352\,
            in2 => \N__23675\,
            in3 => \N__24423\,
            lcout => OPEN,
            ltout => \ALU.N_757_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNICMQ94_10_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35207\,
            in1 => \_gnd_net_\,
            in2 => \N__23672\,
            in3 => \N__23669\,
            lcout => \ALU.aluOut_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_2_rep1_e_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27185\,
            lcout => \aluOperand1_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47680\,
            ce => \N__27697\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIQ5T31_5_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__27321\,
            in1 => \N__48965\,
            in2 => \N__36440\,
            in3 => \N__27128\,
            lcout => \ALU.dout_6_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGUO51_6_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__35013\,
            in1 => \N__43373\,
            in2 => \N__45622\,
            in3 => \N__23720\,
            lcout => OPEN,
            ltout => \ALU.N_865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDHB63_6_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32995\,
            in2 => \N__23651\,
            in3 => \N__23789\,
            lcout => \ALU.operand2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIKC1M_6_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__27897\,
            in1 => \N__28622\,
            in2 => \N__31044\,
            in3 => \N__32049\,
            lcout => OPEN,
            ltout => \ALU.operand2_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIBICH1_6_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__28975\,
            in1 => \N__29015\,
            in2 => \N__23792\,
            in3 => \N__35012\,
            lcout => \ALU.N_817\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDTEA7_6_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__26690\,
            in1 => \N__26279\,
            in2 => \N__24315\,
            in3 => \N__46622\,
            lcout => \ALU.a6_b_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKTLA7_6_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__26278\,
            in1 => \N__41809\,
            in2 => \N__24313\,
            in3 => \N__26689\,
            lcout => \ALU.a3_b_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNINI7O_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__36419\,
            in1 => \N__45129\,
            in2 => \N__31045\,
            in3 => \N__48815\,
            lcout => \ALU.operand2_6_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNII4LL_3_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29072\,
            in1 => \N__31879\,
            in2 => \_gnd_net_\,
            in3 => \N__32069\,
            lcout => \ALU.g_RNII4LLZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID7IK1_3_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__35671\,
            in1 => \N__45158\,
            in2 => \N__45185\,
            in3 => \N__27365\,
            lcout => OPEN,
            ltout => \ALU.N_750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI932E3_3_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__23825\,
            in1 => \_gnd_net_\,
            in2 => \N__23714\,
            in3 => \N__35221\,
            lcout => \ALU.aluOut_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7PG73_3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__44987\,
            in1 => \N__43247\,
            in2 => \N__33103\,
            in3 => \N__23810\,
            lcout => \ALU.operand2_3\,
            ltout => \ALU.operand2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1CMM3_3_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__23938\,
            in1 => \_gnd_net_\,
            in2 => \N__23711\,
            in3 => \N__25221\,
            lcout => \ALU.N_237_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKAQB7_3_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__23974\,
            in1 => \N__23940\,
            in2 => \N__24316\,
            in3 => \N__41861\,
            lcout => \ALU.a3_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHR4B7_3_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__23937\,
            in1 => \N__36844\,
            in2 => \N__24314\,
            in3 => \N__23972\,
            lcout => \ALU.a2_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC8CA7_3_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011000101"
        )
    port map (
            in0 => \N__23973\,
            in1 => \N__23939\,
            in2 => \N__26641\,
            in3 => \N__41860\,
            lcout => \ALU.un2_addsub_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDK21B_3_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23852\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41667\,
            lcout => \ALU.d_RNIDK21BZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI3H7N_3_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__44908\,
            in1 => \N__27029\,
            in2 => \N__27120\,
            in3 => \N__28637\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIOGML1_3_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__31883\,
            in1 => \N__35706\,
            in2 => \N__23828\,
            in3 => \N__29071\,
            lcout => \ALU.N_702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNITOVJ_3_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44907\,
            in1 => \N__28636\,
            in2 => \_gnd_net_\,
            in3 => \N__34891\,
            lcout => OPEN,
            ltout => \ALU.e_RNITOVJZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIGBPU1_3_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__31264\,
            in1 => \N__23819\,
            in2 => \N__23813\,
            in3 => \N__35028\,
            lcout => \ALU.operand2_7_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_6_c_RNIUKMKR_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42530\,
            in1 => \N__40145\,
            in2 => \_gnd_net_\,
            in3 => \N__23804\,
            lcout => \ALU.un9_addsub_cry_6_c_RNIUKMKRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_63_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010001000"
        )
    port map (
            in0 => \N__24545\,
            in1 => \N__24533\,
            in2 => \N__46682\,
            in3 => \N__37718\,
            lcout => \ALU.madd_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_2_l_fx_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24500\,
            in1 => \N__24488\,
            in2 => \N__25838\,
            in3 => \N__24470\,
            lcout => \ALU.madd_axb_2_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_9_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48597\,
            in1 => \N__36275\,
            in2 => \N__46162\,
            in3 => \N__36205\,
            lcout => \ALU.hZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47690\,
            ce => \N__45574\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2B0L_9_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32817\,
            in1 => \N__32798\,
            in2 => \_gnd_net_\,
            in3 => \N__45338\,
            lcout => \ALU.d_RNI2B0LZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIORSD1_15_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25912\,
            in1 => \N__28495\,
            in2 => \_gnd_net_\,
            in3 => \N__45337\,
            lcout => \ALU.b_RNIORSD1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNII1LU_10_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45336\,
            in1 => \N__24431\,
            in2 => \_gnd_net_\,
            in3 => \N__28427\,
            lcout => \ALU.d_RNII1LUZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO00L_4_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36535\,
            in1 => \N__45335\,
            in2 => \_gnd_net_\,
            in3 => \N__28990\,
            lcout => \ALU.d_RNIO00LZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_8_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48105\,
            in1 => \N__47888\,
            in2 => \_gnd_net_\,
            in3 => \N__47778\,
            lcout => \ALU.dZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47606\,
            ce => \N__43324\,
            sr => \_gnd_net_\
        );

    \FTDI.gap_0_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29206\,
            in2 => \_gnd_net_\,
            in3 => \N__29195\,
            lcout => \FTDI.gapZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_2_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29570\,
            in1 => \N__29587\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => \FTDI.baudAccZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNO_0_0_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110100"
        )
    port map (
            in0 => \N__24627\,
            in1 => \N__24776\,
            in2 => \N__29266\,
            in3 => \N__24722\,
            lcout => OPEN,
            ltout => \FTDI.N_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_0_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110001000"
        )
    port map (
            in0 => \N__29262\,
            in1 => \N__24632\,
            in2 => \N__24746\,
            in3 => \N__24681\,
            lcout => \FTDI.RXstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_1_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000010000000"
        )
    port map (
            in0 => \N__24682\,
            in1 => \N__29261\,
            in2 => \N__24645\,
            in3 => \N__24723\,
            lcout => \FTDI.RXstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_3_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110011101110"
        )
    port map (
            in0 => \N__24701\,
            in1 => \N__24631\,
            in2 => \N__29267\,
            in3 => \N__24680\,
            lcout => \FTDI.RXstateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2s2_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38973\,
            in2 => \_gnd_net_\,
            in3 => \N__44121\,
            lcout => \ALU.a_15_sm0\,
            ltout => \ALU.a_15_sm0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_12_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110101"
        )
    port map (
            in0 => \N__24596\,
            in1 => \_gnd_net_\,
            in2 => \N__24602\,
            in3 => \N__43900\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNISG1SC_12_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011110000110"
        )
    port map (
            in0 => \N__25378\,
            in1 => \N__47220\,
            in2 => \N__24599\,
            in3 => \N__40849\,
            lcout => \ALU.a_15_m2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m4_bm_1_2_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__24595\,
            in1 => \N__47210\,
            in2 => \_gnd_net_\,
            in3 => \N__43899\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_bm_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIII58A_2_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011110000110"
        )
    port map (
            in0 => \N__47211\,
            in1 => \N__36937\,
            in2 => \N__24833\,
            in3 => \N__37256\,
            lcout => \ALU.d_RNIII58AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITBSF7_3_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__36936\,
            in1 => \N__39005\,
            in2 => \N__43727\,
            in3 => \N__42014\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI870EE_5_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__39006\,
            in1 => \N__40429\,
            in2 => \N__24821\,
            in3 => \N__42998\,
            lcout => \ALU.N_470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFE9GA_0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38974\,
            in1 => \N__27235\,
            in2 => \_gnd_net_\,
            in3 => \N__24809\,
            lcout => \ALU.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3DJU7_14_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43676\,
            in1 => \N__40627\,
            in2 => \_gnd_net_\,
            in3 => \N__40747\,
            lcout => \ALU.N_589\,
            ltout => \ALU.N_589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI72MIC_0_15_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__39017\,
            in1 => \N__38730\,
            in2 => \N__24797\,
            in3 => \N__30478\,
            lcout => OPEN,
            ltout => \ALU.rshift_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI6PLSH_13_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111010001"
        )
    port map (
            in0 => \N__25235\,
            in1 => \N__43150\,
            in2 => \N__24794\,
            in3 => \N__44518\,
            lcout => \ALU.a_15_m3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI6KSGG_11_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39016\,
            in1 => \N__30495\,
            in2 => \_gnd_net_\,
            in3 => \N__25241\,
            lcout => \ALU.N_576\,
            ltout => \ALU.N_576_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIA9V4L_0_15_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__30479\,
            in1 => \N__38731\,
            in2 => \N__24779\,
            in3 => \N__39018\,
            lcout => OPEN,
            ltout => \ALU.N_636_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNILI6TQ_11_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110011"
        )
    port map (
            in0 => \N__44519\,
            in1 => \N__43151\,
            in2 => \N__25418\,
            in3 => \N__25415\,
            lcout => \ALU.a_15_m3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIT87FA1_7_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__43152\,
            in1 => \N__27383\,
            in2 => \_gnd_net_\,
            in3 => \N__25394\,
            lcout => \ALU.d_RNIT87FA1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIID898_11_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43707\,
            in1 => \N__39390\,
            in2 => \_gnd_net_\,
            in3 => \N__25377\,
            lcout => \ALU.N_462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5RLE5_13_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__25010\,
            in1 => \_gnd_net_\,
            in2 => \N__26601\,
            in3 => \N__25039\,
            lcout => \ALU.N_177_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIURPF4_13_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__40752\,
            in1 => \_gnd_net_\,
            in2 => \N__25052\,
            in3 => \N__29412\,
            lcout => \ALU.N_270_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m174_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001111111"
        )
    port map (
            in0 => \N__30211\,
            in1 => \N__25204\,
            in2 => \N__30238\,
            in3 => \N__29741\,
            lcout => \ALU.N_175_0\,
            ltout => \ALU.N_175_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISHKD9_13_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101001011001"
        )
    port map (
            in0 => \N__40751\,
            in1 => \N__26553\,
            in2 => \N__25013\,
            in3 => \N__25009\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9FOTE_13_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24980\,
            in3 => \N__24977\,
            lcout => \ALU.d_RNI9FOTEZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEG675_11_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100110011"
        )
    port map (
            in0 => \N__24905\,
            in1 => \N__31181\,
            in2 => \N__29438\,
            in3 => \N__26554\,
            lcout => \ALU.N_186_0_i\,
            ltout => \ALU.N_186_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIA7OEE_11_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__39388\,
            in1 => \_gnd_net_\,
            in2 => \N__25574\,
            in3 => \N__39472\,
            lcout => \ALU.c_RNIA7OEEZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_29_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__41359\,
            in1 => \N__41214\,
            in2 => \N__25556\,
            in3 => \N__30234\,
            lcout => \ctrlOut_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47625\,
            ce => \N__41062\,
            sr => \_gnd_net_\
        );

    \ALU.h_12_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48436\,
            in1 => \N__34076\,
            in2 => \N__45991\,
            in3 => \N__34030\,
            lcout => \ALU.hZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47632\,
            ce => \N__45498\,
            sr => \_gnd_net_\
        );

    \ALU.a_RNIFPBO_12_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45126\,
            in1 => \N__28561\,
            in2 => \_gnd_net_\,
            in3 => \N__28207\,
            lcout => \ALU.a_RNIFPBOZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIM5LU_12_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25492\,
            in1 => \N__45333\,
            in2 => \_gnd_net_\,
            in3 => \N__28390\,
            lcout => \ALU.d_RNIM5LUZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJ949_12_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45127\,
            in1 => \N__33958\,
            in2 => \_gnd_net_\,
            in3 => \N__31282\,
            lcout => OPEN,
            ltout => \ALU.c_RNIJ949Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI693U1_12_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__33084\,
            in1 => \N__34494\,
            in2 => \N__25481\,
            in3 => \N__25478\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI05RP4_12_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__32991\,
            in1 => \N__25472\,
            in2 => \N__25466\,
            in3 => \N__28328\,
            lcout => \ALU.operand2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7GCMD22_8_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__25664\,
            in1 => \N__26108\,
            in2 => \N__45989\,
            in3 => \N__26132\,
            lcout => \ALU.d_RNI7GCMD22Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPCSJD1_8_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44187\,
            in1 => \N__25712\,
            in2 => \_gnd_net_\,
            in3 => \N__25697\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIM0ETK2_8_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25685\,
            in1 => \_gnd_net_\,
            in2 => \N__25667\,
            in3 => \N__46394\,
            lcout => \ALU.a_15_m5_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIRM7O_8_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__47720\,
            in1 => \N__31043\,
            in2 => \N__25658\,
            in3 => \N__45122\,
            lcout => OPEN,
            ltout => \ALU.operand2_6_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQU7D1_8_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__25585\,
            in1 => \N__25627\,
            in2 => \N__25607\,
            in3 => \N__34496\,
            lcout => \ALU.N_867\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_8_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48434\,
            in1 => \N__47864\,
            in2 => \_gnd_net_\,
            in3 => \N__47756\,
            lcout => \ALU.hZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47638\,
            ce => \N__45525\,
            sr => \_gnd_net_\
        );

    \ALU.f_10_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48635\,
            in1 => \N__34310\,
            in2 => \N__46076\,
            in3 => \N__34404\,
            lcout => \ALU.fZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.f_11_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48638\,
            in1 => \N__34245\,
            in2 => \N__46080\,
            in3 => \N__34174\,
            lcout => \ALU.fZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.f_12_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101000101"
        )
    port map (
            in0 => \N__34086\,
            in1 => \N__48641\,
            in2 => \N__46077\,
            in3 => \N__34021\,
            lcout => \ALU.fZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.f_14_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48640\,
            in1 => \N__33816\,
            in2 => \N__46082\,
            in3 => \N__33749\,
            lcout => \ALU.fZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.f_15_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48636\,
            in1 => \N__33655\,
            in2 => \N__46078\,
            in3 => \N__33602\,
            lcout => \ALU.fZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.f_13_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48639\,
            in1 => \N__33935\,
            in2 => \N__46081\,
            in3 => \N__33873\,
            lcout => \ALU.fZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.f_9_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48637\,
            in1 => \N__36268\,
            in2 => \N__46079\,
            in3 => \N__36194\,
            lcout => \ALU.fZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47644\,
            ce => \N__36376\,
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_0_0_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25892\,
            in2 => \N__36662\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \ALU.madd_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_1_0_s_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33113\,
            in2 => \N__25877\,
            in3 => \N__25856\,
            lcout => \ALU.mult_2\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_0\,
            carryout => \ALU.madd_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_2_s_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25853\,
            in2 => \N__25831\,
            in3 => \N__25796\,
            lcout => \ALU.mult_3\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_1\,
            carryout => \ALU.madd_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_3_s_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25793\,
            in2 => \N__25781\,
            in3 => \N__25760\,
            lcout => \ALU.mult_4\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_2\,
            carryout => \ALU.madd_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_4_s_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25757\,
            in2 => \N__25742\,
            in3 => \N__25715\,
            lcout => \ALU.mult_5\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_3\,
            carryout => \ALU.madd_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_5_s_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26179\,
            in2 => \N__26159\,
            in3 => \N__26138\,
            lcout => \ALU.mult_6\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_4\,
            carryout => \ALU.madd_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_5_THRU_LUT4_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42349\,
            in2 => \_gnd_net_\,
            in3 => \N__26135\,
            lcout => \ALU.madd_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_5\,
            carryout => \ALU.madd_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_6_THRU_LUT4_0_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26128\,
            in2 => \_gnd_net_\,
            in3 => \N__26099\,
            lcout => \ALU.madd_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_6\,
            carryout => \ALU.madd_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_8_s_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26096\,
            in2 => \N__26078\,
            in3 => \N__26054\,
            lcout => \ALU.mult_9\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \ALU.madd_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_9_0_s_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26051\,
            in2 => \N__26039\,
            in3 => \N__26018\,
            lcout => \ALU.mult_10\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_8\,
            carryout => \ALU.madd_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_10_0_s_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26015\,
            in2 => \N__25997\,
            in3 => \N__25982\,
            lcout => \ALU.mult_11\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_9\,
            carryout => \ALU.madd_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_11_s_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25979\,
            in3 => \N__25964\,
            lcout => \ALU.mult_12\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_10\,
            carryout => \ALU.madd_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_12_s_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25961\,
            in2 => \N__25943\,
            in3 => \N__25919\,
            lcout => \ALU.mult_13\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_11\,
            carryout => \ALU.madd_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_13_0_s_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26786\,
            in2 => \N__26771\,
            in3 => \N__26753\,
            lcout => \ALU.mult_14\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_12\,
            carryout => \ALU.madd_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_s_14_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26750\,
            in2 => \_gnd_net_\,
            in3 => \N__26735\,
            lcout => \ALU.mult_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3O5R3_6_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__26728\,
            in1 => \N__26650\,
            in2 => \_gnd_net_\,
            in3 => \N__26253\,
            lcout => \ALU.N_219_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIS5U41_15_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__35871\,
            in1 => \N__31361\,
            in2 => \N__35554\,
            in3 => \N__31745\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI7JQF1_15_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35299\,
            in1 => \N__33539\,
            in2 => \N__26192\,
            in3 => \N__31523\,
            lcout => \ALU.N_714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_e_0_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27195\,
            lcout => \aluOperand1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47664\,
            ce => \N__27723\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIM2101_2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__31963\,
            in1 => \N__35870\,
            in2 => \N__35531\,
            in3 => \N__36458\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIR8K91_2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__31427\,
            in1 => \N__35298\,
            in2 => \N__26189\,
            in3 => \N__42038\,
            lcout => OPEN,
            ltout => \ALU.N_749_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6KCD3_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35202\,
            in2 => \N__26186\,
            in3 => \N__26918\,
            lcout => \ALU.aluOut_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNI70VV1_2_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001010101"
        )
    port map (
            in0 => \N__26912\,
            in1 => \N__31901\,
            in2 => \N__29096\,
            in3 => \N__35297\,
            lcout => \ALU.N_701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI40I81_2_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__35853\,
            in1 => \N__28758\,
            in2 => \N__35966\,
            in3 => \N__28781\,
            lcout => \ALU.dout_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_2_rep2_e_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27196\,
            lcout => \aluOperand1_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47671\,
            ce => \N__27719\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIGGOA1_7_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__35852\,
            in1 => \N__36391\,
            in2 => \N__35965\,
            in3 => \N__48655\,
            lcout => \ALU.dout_6_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_1_rep1_e_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aluOperand1_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47671\,
            ce => \N__27719\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIDCNA1_6_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__27336\,
            in1 => \N__36415\,
            in2 => \N__35875\,
            in3 => \N__48811\,
            lcout => \ALU.dout_6_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIQQJ01_7_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__48656\,
            in1 => \_gnd_net_\,
            in2 => \N__36395\,
            in3 => \N__45313\,
            lcout => \ALU.f_RNIQQJ01Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_e_0_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26880\,
            lcout => \aluOperand1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47671\,
            ce => \N__27719\,
            sr => \_gnd_net_\
        );

    \ALU.b_RNIEHSD1_10_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26826\,
            in1 => \N__28518\,
            in2 => \_gnd_net_\,
            in3 => \N__45314\,
            lcout => \ALU.b_RNIEHSD1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48618\,
            in1 => \N__42311\,
            in2 => \_gnd_net_\,
            in3 => \N__42233\,
            lcout => a_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.a_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48615\,
            in1 => \N__40994\,
            in2 => \_gnd_net_\,
            in3 => \N__36605\,
            lcout => a_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.a_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42163\,
            in1 => \N__48616\,
            in2 => \_gnd_net_\,
            in3 => \N__42079\,
            lcout => a_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.a_4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49281\,
            in1 => \N__49220\,
            in2 => \_gnd_net_\,
            in3 => \N__48617\,
            lcout => a_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.a_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49101\,
            in1 => \N__48620\,
            in2 => \_gnd_net_\,
            in3 => \N__49046\,
            lcout => a_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.a_6_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48619\,
            in1 => \N__48891\,
            in2 => \_gnd_net_\,
            in3 => \N__48942\,
            lcout => a_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.a_7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48770\,
            in1 => \N__48716\,
            in2 => \_gnd_net_\,
            in3 => \N__48621\,
            lcout => a_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47675\,
            ce => \N__44870\,
            sr => \_gnd_net_\
        );

    \ALU.e_RNI5J7N_4_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__27131\,
            in1 => \N__27924\,
            in2 => \N__27028\,
            in3 => \N__26959\,
            lcout => \ALU.dout_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_4_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48420\,
            in1 => \N__49286\,
            in2 => \_gnd_net_\,
            in3 => \N__49217\,
            lcout => \ALU.eZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47681\,
            ce => \N__32444\,
            sr => \_gnd_net_\
        );

    \ALU.e_RNIS97J_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27011\,
            in1 => \N__44586\,
            in2 => \_gnd_net_\,
            in3 => \N__26932\,
            lcout => \ALU.e_RNIS97JZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_1_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48419\,
            in1 => \N__40998\,
            in2 => \_gnd_net_\,
            in3 => \N__36614\,
            lcout => \ALU.eZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47681\,
            ce => \N__32444\,
            sr => \_gnd_net_\
        );

    \ALU.g_RNI0MJN_1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29110\,
            in1 => \_gnd_net_\,
            in2 => \N__27027\,
            in3 => \N__31921\,
            lcout => \ALU.g_RNI0MJNZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIM1T31_3_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__27338\,
            in1 => \N__49310\,
            in2 => \N__43268\,
            in3 => \N__27130\,
            lcout => \ALU.dout_6_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIO3T31_4_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__27132\,
            in1 => \N__45410\,
            in2 => \N__27348\,
            in3 => \N__49151\,
            lcout => \ALU.dout_6_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIE5EP3_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__27275\,
            in1 => \N__35135\,
            in2 => \N__43769\,
            in3 => \N__27263\,
            lcout => \ALU.N_404_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQQAK1_6_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__45623\,
            in1 => \N__43372\,
            in2 => \N__27212\,
            in3 => \N__35356\,
            lcout => OPEN,
            ltout => \ALU.N_753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI23RD3_6_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35134\,
            in2 => \N__27200\,
            in3 => \N__27764\,
            lcout => \ALU.aluOut_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_fast_e_2_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27197\,
            lcout => \aluOperand1_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47684\,
            ce => \N__27728\,
            sr => \_gnd_net_\
        );

    \ALU.e_RNI9N7N_6_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__28621\,
            in1 => \N__27127\,
            in2 => \N__27026\,
            in3 => \N__27898\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNI4TML1_6_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__35713\,
            in1 => \N__28976\,
            in2 => \N__27767\,
            in3 => \N__29011\,
            lcout => \ALU.N_705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_e_0_0_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27758\,
            lcout => \aluOperand1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47684\,
            ce => \N__27728\,
            sr => \_gnd_net_\
        );

    \ALU.c_8_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48074\,
            in1 => \N__47887\,
            in2 => \_gnd_net_\,
            in3 => \N__47798\,
            lcout => \ALU.cZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47600\,
            ce => \N__31498\,
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_0_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__29522\,
            in1 => \_gnd_net_\,
            in2 => \N__44749\,
            in3 => \N__30380\,
            lcout => \FTDI.TXstate_e_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI72MIC_15_LC_10_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__39022\,
            in1 => \N__30477\,
            in2 => \N__38734\,
            in3 => \N__30503\,
            lcout => OPEN,
            ltout => \ALU.c_RNI72MICZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBHJVC1_15_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44479\,
            in2 => \N__27620\,
            in3 => \N__27617\,
            lcout => \ALU.rshift_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_0_LC_10_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29586\,
            in2 => \_gnd_net_\,
            in3 => \N__30418\,
            lcout => \FTDI.baudAccZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6QT5G_9_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__27809\,
            in1 => \N__39860\,
            in2 => \N__39084\,
            in3 => \N__27607\,
            lcout => \ALU.N_475\,
            ltout => \ALU.N_475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIGVM161_15_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__44395\,
            in1 => \N__27827\,
            in2 => \N__27386\,
            in3 => \N__27803\,
            lcout => \ALU.rshift_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI4JFV4_15_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__30469\,
            in1 => \N__44394\,
            in2 => \N__38714\,
            in3 => \N__39011\,
            lcout => \ALU.rshift_15_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI83IG7_0_3_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__43690\,
            in1 => \N__42013\,
            in2 => \N__39069\,
            in3 => \N__42991\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4MEEE_6_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__39061\,
            in1 => \N__40428\,
            in2 => \N__27821\,
            in3 => \N__46716\,
            lcout => OPEN,
            ltout => \ALU.N_471_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9DPVU_6_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38648\,
            in2 => \N__27818\,
            in3 => \N__27815\,
            lcout => \ALU.d_RNI9DPVUZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIT1MQ7_7_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__43689\,
            in1 => \N__40119\,
            in2 => \N__39083\,
            in3 => \N__46975\,
            lcout => \ALU.rshift_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIA9V4L_15_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__39010\,
            in1 => \N__30470\,
            in2 => \N__38715\,
            in3 => \N__27802\,
            lcout => \ALU.c_RNIA9V4LZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6I9AJ2_5_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46363\,
            in1 => \N__27947\,
            in2 => \_gnd_net_\,
            in3 => \N__29528\,
            lcout => OPEN,
            ltout => \ALU.a_15_m5_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIH1NE6F_5_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45923\,
            in2 => \N__27794\,
            in3 => \N__27791\,
            lcout => \ALU.d_RNIH1NE6FZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRCOSL2_9_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46362\,
            in1 => \N__30428\,
            in2 => \_gnd_net_\,
            in3 => \N__27776\,
            lcout => \ALU.a_15_m5_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_5_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__47178\,
            in1 => \N__44151\,
            in2 => \N__43929\,
            in3 => \N__43726\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISQNAA_5_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001100111"
        )
    port map (
            in0 => \N__47179\,
            in1 => \N__40401\,
            in2 => \N__28100\,
            in3 => \N__28097\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQO6O01_5_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__44500\,
            in1 => \N__44152\,
            in2 => \N__27968\,
            in3 => \N__27965\,
            lcout => \ALU.a_15_m4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28937\,
            lcout => \TXbufferZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47613\,
            ce => \N__44551\,
            sr => \_gnd_net_\
        );

    \TXbuffer_2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28769\,
            lcout => \TXbufferZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47613\,
            ce => \N__44551\,
            sr => \_gnd_net_\
        );

    \TXbuffer_3_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44915\,
            lcout => \TXbufferZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47613\,
            ce => \N__44551\,
            sr => \_gnd_net_\
        );

    \TXbuffer_4_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27940\,
            lcout => \TXbufferZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47613\,
            ce => \N__44551\,
            sr => \_gnd_net_\
        );

    \TXbuffer_6_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27908\,
            lcout => \TXbufferZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47613\,
            ce => \N__44551\,
            sr => \_gnd_net_\
        );

    \TXbuffer_7_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27874\,
            lcout => \TXbufferZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47613\,
            ce => \N__44551\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1BC602_12_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44228\,
            in1 => \N__27836\,
            in2 => \_gnd_net_\,
            in3 => \N__28166\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIC8RDN2_12_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46383\,
            in2 => \N__28238\,
            in3 => \N__28187\,
            lcout => \c_RNIC8RDN2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_11_c_RNIQ9LMU_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__42459\,
            in1 => \N__40787\,
            in2 => \_gnd_net_\,
            in3 => \N__28235\,
            lcout => OPEN,
            ltout => \un2_addsub_cry_11_c_RNIQ9LMU_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNIGPL5M3_0_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48339\,
            in2 => \N__28223\,
            in3 => \N__28220\,
            lcout => \aluOperation_RNIGPL5M3_0\,
            ltout => \aluOperation_RNIGPL5M3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_12_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48340\,
            in1 => \N__45836\,
            in2 => \N__28214\,
            in3 => \N__34031\,
            lcout => \ALU.aZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47619\,
            ce => \N__44849\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIC6T9M_12_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100000011"
        )
    port map (
            in0 => \N__44437\,
            in1 => \N__28196\,
            in2 => \N__43189\,
            in3 => \N__43231\,
            lcout => \ALU.a_15_m3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6VHRI1_0_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44520\,
            in1 => \N__44959\,
            in2 => \_gnd_net_\,
            in3 => \N__28181\,
            lcout => \ALU.lshift_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_m2_1_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__45281\,
            in1 => \N__28126\,
            in2 => \N__28159\,
            in3 => \N__35033\,
            lcout => \ALU.g0_0_0_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_9_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48435\,
            in1 => \N__36257\,
            in2 => \N__46084\,
            in3 => \N__36204\,
            lcout => \ALU.bZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47626\,
            ce => \N__47393\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIUUJ01_9_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45284\,
            in2 => \N__28158\,
            in3 => \N__28125\,
            lcout => \ALU.f_RNIUUJ01Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_11_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101000101"
        )
    port map (
            in0 => \N__34246\,
            in1 => \N__48411\,
            in2 => \N__46083\,
            in3 => \N__34175\,
            lcout => \ALU.bZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47626\,
            ce => \N__47393\,
            sr => \_gnd_net_\
        );

    \ALU.b_12_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48409\,
            in1 => \N__45993\,
            in2 => \N__34088\,
            in3 => \N__34026\,
            lcout => \ALU.bZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47626\,
            ce => \N__47393\,
            sr => \_gnd_net_\
        );

    \ALU.b_RNIILSD1_12_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__45283\,
            in1 => \N__28363\,
            in2 => \_gnd_net_\,
            in3 => \N__28342\,
            lcout => \ALU.b_RNIILSD1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_14_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48410\,
            in1 => \N__33815\,
            in2 => \N__46118\,
            in3 => \N__33756\,
            lcout => \ALU.bZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47626\,
            ce => \N__47393\,
            sr => \_gnd_net_\
        );

    \ALU.b_RNIMPSD1_14_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28309\,
            in1 => \N__28288\,
            in2 => \_gnd_net_\,
            in3 => \N__45282\,
            lcout => \ALU.b_RNIMPSD1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8DRP4_13_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001010"
        )
    port map (
            in0 => \N__32983\,
            in1 => \N__28256\,
            in2 => \N__28250\,
            in3 => \N__31096\,
            lcout => OPEN,
            ltout => \ALU.g0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA7959_13_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__29612\,
            in1 => \N__29966\,
            in2 => \N__28277\,
            in3 => \N__38041\,
            lcout => \ALU.N_703_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIKNSD1_0_13_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45279\,
            in1 => \_gnd_net_\,
            in2 => \N__35614\,
            in3 => \N__35783\,
            lcout => \ALU.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO7LU_0_13_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35424\,
            in1 => \N__35461\,
            in2 => \_gnd_net_\,
            in3 => \N__45278\,
            lcout => \ALU.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__34799\,
            in1 => \N__32213\,
            in2 => \N__34721\,
            in3 => \N__45280\,
            lcout => \aluOperand2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIGJSD1_11_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45276\,
            in1 => \N__28468\,
            in2 => \_gnd_net_\,
            in3 => \N__28450\,
            lcout => \ALU.b_RNIGJSD1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIKNSD1_13_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35782\,
            in1 => \N__35607\,
            in2 => \_gnd_net_\,
            in3 => \N__45277\,
            lcout => \ALU.b_RNIKNSD1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_10_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48344\,
            in1 => \N__34343\,
            in2 => \N__46189\,
            in3 => \N__34395\,
            lcout => \ALU.dZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.d_11_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101010001"
        )
    port map (
            in0 => \N__34250\,
            in1 => \N__46163\,
            in2 => \N__48575\,
            in3 => \N__34160\,
            lcout => \ALU.dZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.d_12_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48345\,
            in1 => \N__34087\,
            in2 => \N__46190\,
            in3 => \N__34010\,
            lcout => \ALU.dZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.d_14_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101010001"
        )
    port map (
            in0 => \N__33812\,
            in1 => \N__46165\,
            in2 => \N__48576\,
            in3 => \N__33740\,
            lcout => \ALU.dZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.d_15_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48346\,
            in1 => \N__33659\,
            in2 => \N__46191\,
            in3 => \N__33591\,
            lcout => \ALU.dZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.d_13_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48412\,
            in1 => \N__46164\,
            in2 => \N__33941\,
            in3 => \N__33864\,
            lcout => \ALU.dZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.d_9_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48347\,
            in1 => \N__36260\,
            in2 => \N__46192\,
            in3 => \N__36178\,
            lcout => \ALU.dZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47639\,
            ce => \N__43345\,
            sr => \_gnd_net_\
        );

    \ALU.e_10_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111000101"
        )
    port map (
            in0 => \N__34344\,
            in1 => \N__34384\,
            in2 => \N__46147\,
            in3 => \N__48560\,
            lcout => \ALU.eZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => \N__32457\,
            sr => \_gnd_net_\
        );

    \ALU.e_11_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101010001"
        )
    port map (
            in0 => \N__34247\,
            in1 => \N__46060\,
            in2 => \N__48634\,
            in3 => \N__34147\,
            lcout => \ALU.eZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => \N__32457\,
            sr => \_gnd_net_\
        );

    \ALU.e_12_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48572\,
            in1 => \N__34090\,
            in2 => \N__46148\,
            in3 => \N__34000\,
            lcout => \ALU.eZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => \N__32457\,
            sr => \_gnd_net_\
        );

    \ALU.e_13_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48555\,
            in1 => \N__33934\,
            in2 => \N__46150\,
            in3 => \N__33853\,
            lcout => \ALU.eZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => \N__32457\,
            sr => \_gnd_net_\
        );

    \ALU.e_14_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48573\,
            in1 => \N__33814\,
            in2 => \N__46149\,
            in3 => \N__33727\,
            lcout => \ALU.eZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => \N__32457\,
            sr => \_gnd_net_\
        );

    \ALU.e_15_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48556\,
            in1 => \N__33660\,
            in2 => \N__46151\,
            in3 => \N__33589\,
            lcout => \ALU.eZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47645\,
            ce => \N__32457\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPER7_5_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45063\,
            in1 => \N__31396\,
            in2 => \_gnd_net_\,
            in3 => \N__43396\,
            lcout => \ALU.d_RNIPER7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_10_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48076\,
            in1 => \N__34345\,
            in2 => \N__46193\,
            in3 => \N__34394\,
            lcout => \ALU.bZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47402\,
            sr => \_gnd_net_\
        );

    \ALU.b_15_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48092\,
            in1 => \N__33661\,
            in2 => \N__46122\,
            in3 => \N__33590\,
            lcout => \ALU.bZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47402\,
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_12_c_RNIG3PMU_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__42518\,
            in1 => \N__40649\,
            in2 => \_gnd_net_\,
            in3 => \N__28700\,
            lcout => OPEN,
            ltout => \un2_addsub_cry_12_c_RNIG3PMU_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNI2J9SL3_0_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48075\,
            in2 => \N__28688\,
            in3 => \N__28685\,
            lcout => \aluOperation_RNI2J9SL3_0\,
            ltout => \aluOperation_RNI2J9SL3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_13_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48077\,
            in1 => \N__46046\,
            in2 => \N__28670\,
            in3 => \N__33863\,
            lcout => \ALU.bZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47402\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIFMN04_2_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46045\,
            in1 => \N__28667\,
            in2 => \_gnd_net_\,
            in3 => \N__28655\,
            lcout => \ALU.d_RNIIFMN04Z0Z_2\,
            ltout => \ALU.d_RNIIFMN04Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_2_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42151\,
            in2 => \N__28640\,
            in3 => \N__48093\,
            lcout => \ALU.bZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47651\,
            ce => \N__47402\,
            sr => \_gnd_net_\
        );

    \ALU.e_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48430\,
            in1 => \N__42321\,
            in2 => \_gnd_net_\,
            in3 => \N__42252\,
            lcout => \ALU.eZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => \N__32468\,
            sr => \_gnd_net_\
        );

    \ALU.e_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48567\,
            in1 => \N__42162\,
            in2 => \_gnd_net_\,
            in3 => \N__42078\,
            lcout => \ALU.eZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => \N__32468\,
            sr => \_gnd_net_\
        );

    \ALU.e_3_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48431\,
            in1 => \N__49468\,
            in2 => \_gnd_net_\,
            in3 => \N__49387\,
            lcout => \ALU.eZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => \N__32468\,
            sr => \_gnd_net_\
        );

    \ALU.e_6_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48932\,
            in1 => \N__48432\,
            in2 => \_gnd_net_\,
            in3 => \N__48881\,
            lcout => \ALU.eZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => \N__32468\,
            sr => \_gnd_net_\
        );

    \ALU.e_7_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48713\,
            in1 => \N__48569\,
            in2 => \_gnd_net_\,
            in3 => \N__48777\,
            lcout => \ALU.eZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => \N__32468\,
            sr => \_gnd_net_\
        );

    \ALU.e_8_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48568\,
            in1 => \N__47886\,
            in2 => \_gnd_net_\,
            in3 => \N__47794\,
            lcout => \ALU.eZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47657\,
            ce => \N__32468\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_fast_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__34764\,
            in1 => \N__31014\,
            in2 => \N__34709\,
            in3 => \N__34566\,
            lcout => \aluOperand2_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_1_rep1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__34567\,
            in1 => \N__34765\,
            in2 => \N__34708\,
            in3 => \N__34994\,
            lcout => \aluOperand2_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_fast_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__34867\,
            in1 => \N__32224\,
            in2 => \N__34787\,
            in3 => \N__34685\,
            lcout => \aluOperand2_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIRMVJ_2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__28780\,
            in1 => \N__28759\,
            in2 => \N__34868\,
            in3 => \_gnd_net_\,
            lcout => \ALU.e_RNIRMVJZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIV2CO_2_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29089\,
            in1 => \N__34855\,
            in2 => \_gnd_net_\,
            in3 => \N__31894\,
            lcout => OPEN,
            ltout => \ALU.g_RNIV2COZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIPKSL1_2_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__31013\,
            in1 => \N__31577\,
            in2 => \N__28742\,
            in3 => \N__28739\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAUJU2_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__33089\,
            in1 => \N__28811\,
            in2 => \N__28733\,
            in3 => \N__31949\,
            lcout => \ALU.operand2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNINIVJ_0_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34854\,
            in1 => \N__28948\,
            in2 => \_gnd_net_\,
            in3 => \N__28926\,
            lcout => \ALU.e_RNINIVJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIM8LL_5_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32025\,
            in1 => \N__31825\,
            in2 => \_gnd_net_\,
            in3 => \N__29026\,
            lcout => \ALU.g_RNIM8LLZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI1TVJ_5_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34863\,
            in1 => \N__44628\,
            in2 => \_gnd_net_\,
            in3 => \N__28861\,
            lcout => OPEN,
            ltout => \ALU.e_RNI1TVJZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIOJPU1_5_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__28892\,
            in1 => \N__34993\,
            in2 => \N__28886\,
            in3 => \N__31263\,
            lcout => \ALU.operand2_7_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_5_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48426\,
            in1 => \N__49130\,
            in2 => \_gnd_net_\,
            in3 => \N__49045\,
            lcout => \ALU.eZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47672\,
            ce => \N__32467\,
            sr => \_gnd_net_\
        );

    \ALU.g_RNIRUBO_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29134\,
            in1 => \N__34862\,
            in2 => \_gnd_net_\,
            in3 => \N__31933\,
            lcout => \ALU.g_RNIRUBOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIG6R7_1_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31441\,
            in1 => \N__32027\,
            in2 => \_gnd_net_\,
            in3 => \N__36553\,
            lcout => \ALU.d_RNIG6R7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI45J9_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36554\,
            in1 => \_gnd_net_\,
            in2 => \N__35586\,
            in3 => \N__31442\,
            lcout => \ALU.d_RNI45J9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNII8R7_2_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31423\,
            in1 => \N__32026\,
            in2 => \_gnd_net_\,
            in3 => \N__42034\,
            lcout => \ALU.d_RNII8R7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48631\,
            in1 => \N__42322\,
            in2 => \_gnd_net_\,
            in3 => \N__42254\,
            lcout => \ALU.cZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48421\,
            in1 => \N__41000\,
            in2 => \_gnd_net_\,
            in3 => \N__36613\,
            lcout => \ALU.cZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48632\,
            in1 => \N__42164\,
            in2 => \_gnd_net_\,
            in3 => \N__42092\,
            lcout => \ALU.cZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_3_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48422\,
            in1 => \N__49467\,
            in2 => \_gnd_net_\,
            in3 => \N__49388\,
            lcout => \ALU.cZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_4_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49218\,
            in1 => \N__48424\,
            in2 => \_gnd_net_\,
            in3 => \N__49285\,
            lcout => \ALU.cZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_5_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48423\,
            in1 => \N__49112\,
            in2 => \_gnd_net_\,
            in3 => \N__49047\,
            lcout => \ALU.cZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_6_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48943\,
            in1 => \N__48425\,
            in2 => \_gnd_net_\,
            in3 => \N__48892\,
            lcout => \ALU.cZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.c_7_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48715\,
            in1 => \N__48633\,
            in2 => \_gnd_net_\,
            in3 => \N__48749\,
            lcout => \ALU.cZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47676\,
            ce => \N__31502\,
            sr => \_gnd_net_\
        );

    \ALU.d_4_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48629\,
            in1 => \N__49287\,
            in2 => \_gnd_net_\,
            in3 => \N__49219\,
            lcout => \ALU.dZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47682\,
            ce => \N__43346\,
            sr => \_gnd_net_\
        );

    \ALU.g_6_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48630\,
            in1 => \N__48893\,
            in2 => \_gnd_net_\,
            in3 => \N__48947\,
            lcout => \ALU.gZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47685\,
            ce => \N__36104\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_2_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__29194\,
            in1 => \_gnd_net_\,
            in2 => \N__29219\,
            in3 => \N__29168\,
            lcout => \FTDI.gapZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_1_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__29167\,
            in1 => \N__29215\,
            in2 => \_gnd_net_\,
            in3 => \N__29193\,
            lcout => \FTDI.gapZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNICVLM_0_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30377\,
            in2 => \_gnd_net_\,
            in3 => \N__29518\,
            lcout => \FTDI.N_169_0\,
            ltout => \FTDI.N_169_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_0_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100000011"
        )
    port map (
            in0 => \N__32322\,
            in1 => \N__29159\,
            in2 => \N__29153\,
            in3 => \N__29494\,
            lcout => \FTDI.TXstateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_1_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001001000"
        )
    port map (
            in0 => \N__29495\,
            in1 => \N__44744\,
            in2 => \N__29150\,
            in3 => \N__29597\,
            lcout => \FTDI.TXstateZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_2_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011100000111"
        )
    port map (
            in0 => \N__44719\,
            in1 => \N__29467\,
            in2 => \N__32327\,
            in3 => \N__30379\,
            lcout => OPEN,
            ltout => \FTDI.TXstate_cnst_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_2_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30410\,
            in2 => \N__29141\,
            in3 => \N__30341\,
            lcout => \FTDI.un3_TX_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_1_1_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32321\,
            in2 => \_gnd_net_\,
            in3 => \N__29517\,
            lcout => OPEN,
            ltout => \FTDI.N_217_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_1_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__30378\,
            in1 => \N__44718\,
            in2 => \N__29600\,
            in3 => \N__29493\,
            lcout => \FTDI.N_216_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNINQ101_0_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30384\,
            in1 => \N__29519\,
            in2 => \_gnd_net_\,
            in3 => \N__29490\,
            lcout => \FTDI.N_170_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNIEFF51_0_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29520\,
            in1 => \N__29492\,
            in2 => \N__44748\,
            in3 => \N__32319\,
            lcout => \FTDI.TXready\,
            ltout => \FTDI.TXready_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_1_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29563\,
            in2 => \N__29591\,
            in3 => \N__29588\,
            lcout => \FTDI.baudAccZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID2HKH1_5_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43179\,
            in1 => \N__29552\,
            in2 => \_gnd_net_\,
            in3 => \N__29534\,
            lcout => \ALU.a_15_m3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_3_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30385\,
            in1 => \N__29521\,
            in2 => \_gnd_net_\,
            in3 => \N__29491\,
            lcout => OPEN,
            ltout => \FTDI.TXstate_e_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_3_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001010101010"
        )
    port map (
            in0 => \N__44717\,
            in1 => \N__29468\,
            in2 => \N__29456\,
            in3 => \N__32320\,
            lcout => \FTDI.TXstateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1OCN4_15_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__29453\,
            in1 => \N__32666\,
            in2 => \_gnd_net_\,
            in3 => \N__29437\,
            lcout => OPEN,
            ltout => \ALU.c_RNI1OCN4Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI68L5A_15_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43172\,
            in2 => \N__30560\,
            in3 => \N__30443\,
            lcout => \ALU.a_15_m3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIKUKV3_15_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__30557\,
            in1 => \N__30535\,
            in2 => \N__43747\,
            in3 => \N__35223\,
            lcout => \ALU.N_621_1\,
            ltout => \ALU.N_621_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI8597C_15_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39151\,
            in2 => \N__30506\,
            in3 => \N__30502\,
            lcout => \ALU.N_578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI4JFV4_0_15_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__38713\,
            in1 => \N__39152\,
            in2 => \N__44525\,
            in3 => \N__30471\,
            lcout => \ALU.c_RNI4JFV4_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI36KJ21_9_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100000011"
        )
    port map (
            in0 => \N__44499\,
            in1 => \N__30437\,
            in2 => \N__43184\,
            in3 => \N__31751\,
            lcout => \ALU.d_RNI36KJ21Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_RNINKH42_2_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__30417\,
            in1 => \N__30336\,
            in2 => \N__44768\,
            in3 => \N__30386\,
            lcout => \FTDI.un1_TXstate_0_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXstart_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111010101000"
        )
    port map (
            in0 => \N__30337\,
            in1 => \N__30808\,
            in2 => \N__30322\,
            in3 => \N__41413\,
            lcout => \TXstartZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m326dup_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30807\,
            in1 => \N__41409\,
            in2 => \_gnd_net_\,
            in3 => \N__30315\,
            lcout => m326dup,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g0_7_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30239\,
            in1 => \N__30218\,
            in2 => \N__30025\,
            in3 => \N__29754\,
            lcout => \ALU.N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_RNIB7C_2_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30806\,
            lcout => \testState_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIJTBO_14_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30721\,
            in1 => \N__31378\,
            in2 => \_gnd_net_\,
            in3 => \N__45128\,
            lcout => \ALU.a_RNIJTBOZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_13_c_RNI2LH1U_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__42458\,
            in1 => \N__40538\,
            in2 => \_gnd_net_\,
            in3 => \N__30704\,
            lcout => OPEN,
            ltout => \un2_addsub_cry_13_c_RNI2LH1U_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNIR872K3_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48271\,
            in2 => \N__30686\,
            in3 => \N__30683\,
            lcout => \aluOperation_RNIR872K3_0\,
            ltout => \aluOperation_RNIR872K3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_14_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48272\,
            in1 => \N__45930\,
            in2 => \N__30668\,
            in3 => \N__33757\,
            lcout => \ALU.hZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47614\,
            ce => \N__45567\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIEH3U1_14_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__34495\,
            in1 => \N__31532\,
            in2 => \N__30665\,
            in3 => \N__33065\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGLRP4_14_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__32971\,
            in1 => \N__30566\,
            in2 => \N__30656\,
            in3 => \N__30653\,
            lcout => \ALU.operand2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQ9LU_14_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30610\,
            in1 => \N__30589\,
            in2 => \_gnd_net_\,
            in3 => \N__45322\,
            lcout => \ALU.d_RNIQ9LUZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_8_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48267\,
            in1 => \N__47827\,
            in2 => \_gnd_net_\,
            in3 => \N__47777\,
            lcout => \ALU.aZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47620\,
            ce => \N__44871\,
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_7_c_RNIQIKVO_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42463\,
            in1 => \N__39875\,
            in2 => \_gnd_net_\,
            in3 => \N__31082\,
            lcout => \ALU.un9_addsub_cry_7_c_RNIQIKVOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIOG1M_8_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__31060\,
            in1 => \N__31042\,
            in2 => \N__30973\,
            in3 => \N__32073\,
            lcout => OPEN,
            ltout => \ALU.operand2_3_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIJQCH1_8_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__30937\,
            in1 => \N__30901\,
            in2 => \N__30878\,
            in3 => \N__35030\,
            lcout => \ALU.N_819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m715_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__48265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43728\,
            lcout => \ALU.addsub_0_sqmuxa\,
            ltout => \ALU.addsub_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_8_c_RNIKTS9S_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39623\,
            in1 => \_gnd_net_\,
            in2 => \N__30860\,
            in3 => \N__30857\,
            lcout => OPEN,
            ltout => \ALU.un9_addsub_cry_8_c_RNIKTS9SZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_8_c_RNIPHQ7I3_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__48266\,
            in1 => \_gnd_net_\,
            in2 => \N__30845\,
            in3 => \N__30842\,
            lcout => \ALU.a_15_ns_1_9\,
            ltout => \ALU.a_15_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_9_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100001101"
        )
    port map (
            in0 => \N__45990\,
            in1 => \N__48268\,
            in2 => \N__30833\,
            in3 => \N__36203\,
            lcout => \ALU.aZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47620\,
            ce => \N__44871\,
            sr => \_gnd_net_\
        );

    \ALU.a_RNICNBO_11_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32067\,
            in1 => \N__32482\,
            in2 => \_gnd_net_\,
            in3 => \N__30826\,
            lcout => OPEN,
            ltout => \ALU.a_RNICNBOZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITCKM1_11_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__35031\,
            in1 => \N__31249\,
            in2 => \N__31193\,
            in3 => \N__31118\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJ4CI4_11_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__32902\,
            in1 => \N__31142\,
            in2 => \N__31190\,
            in3 => \N__31187\,
            lcout => \ALU.operand2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIK3LU_11_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45275\,
            in1 => \N__31129\,
            in2 => \_gnd_net_\,
            in3 => \N__31153\,
            lcout => \ALU.d_RNIK3LUZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_11_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48348\,
            in1 => \N__34248\,
            in2 => \N__46117\,
            in3 => \N__34180\,
            lcout => \ALU.hZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47627\,
            ce => \N__45538\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIG749_11_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34105\,
            in1 => \N__32066\,
            in2 => \_gnd_net_\,
            in3 => \N__31300\,
            lcout => \ALU.c_RNIG749Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNILB49_13_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35809\,
            in1 => \N__35794\,
            in2 => \_gnd_net_\,
            in3 => \N__45076\,
            lcout => \ALU.c_RNILB49Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIHRBO_13_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45077\,
            in1 => \N__36031\,
            in2 => \_gnd_net_\,
            in3 => \N__36020\,
            lcout => OPEN,
            ltout => \ALU.a_RNIHRBOZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIAD3U1_13_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__33063\,
            in1 => \N__34468\,
            in2 => \N__31112\,
            in3 => \N__31109\,
            lcout => \ALU.operand2_7_ns_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_2_rep2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__45080\,
            in1 => \N__32214\,
            in2 => \N__34720\,
            in3 => \N__34797\,
            lcout => \aluOperand2_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47634\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIPF49_15_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31522\,
            in1 => \N__45078\,
            in2 => \_gnd_net_\,
            in3 => \N__33535\,
            lcout => \ALU.c_RNIPF49Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNILVBO_15_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45079\,
            in1 => \N__31360\,
            in2 => \_gnd_net_\,
            in3 => \N__31741\,
            lcout => OPEN,
            ltout => \ALU.a_RNILVBOZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIIL3U1_15_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__33064\,
            in1 => \N__34469\,
            in2 => \N__31349\,
            in3 => \N__31346\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIOTRP4_15_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__32946\,
            in1 => \N__33449\,
            in2 => \N__31340\,
            in3 => \N__31337\,
            lcout => \ALU.operand2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_10_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48561\,
            in1 => \N__34346\,
            in2 => \N__46152\,
            in3 => \N__34402\,
            lcout => \ALU.cZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.c_11_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48483\,
            in1 => \N__34249\,
            in2 => \N__46156\,
            in3 => \N__34167\,
            lcout => \ALU.cZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.c_12_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101000101"
        )
    port map (
            in0 => \N__34089\,
            in1 => \N__48485\,
            in2 => \N__46153\,
            in3 => \N__34020\,
            lcout => \ALU.cZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.c_13_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48484\,
            in1 => \N__33921\,
            in2 => \N__46157\,
            in3 => \N__33871\,
            lcout => \ALU.cZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.c_14_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48562\,
            in1 => \N__33813\,
            in2 => \N__46154\,
            in3 => \N__33747\,
            lcout => \ALU.cZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIND49_14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33685\,
            in1 => \N__31543\,
            in2 => \_gnd_net_\,
            in3 => \N__45081\,
            lcout => \ALU.c_RNIND49Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_15_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48563\,
            in1 => \N__33654\,
            in2 => \N__46155\,
            in3 => \N__33601\,
            lcout => \ALU.cZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.c_9_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000011111101"
        )
    port map (
            in0 => \N__46098\,
            in1 => \N__48564\,
            in2 => \N__36202\,
            in3 => \N__36259\,
            lcout => \ALU.cZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47640\,
            ce => \N__31497\,
            sr => \_gnd_net_\
        );

    \ALU.h_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36606\,
            in1 => \N__48095\,
            in2 => \_gnd_net_\,
            in3 => \N__40981\,
            lcout => \ALU.hZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47646\,
            ce => \N__45568\,
            sr => \_gnd_net_\
        );

    \ALU.h_2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48094\,
            in1 => \N__42150\,
            in2 => \_gnd_net_\,
            in3 => \N__42072\,
            lcout => \ALU.hZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47646\,
            ce => \N__45568\,
            sr => \_gnd_net_\
        );

    \ALU.h_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49460\,
            in1 => \N__48096\,
            in2 => \_gnd_net_\,
            in3 => \N__49382\,
            lcout => \ALU.hZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47646\,
            ce => \N__45568\,
            sr => \_gnd_net_\
        );

    \ALU.h_7_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48788\,
            in1 => \N__48700\,
            in2 => \_gnd_net_\,
            in3 => \N__48571\,
            lcout => \ALU.hZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47646\,
            ce => \N__45568\,
            sr => \_gnd_net_\
        );

    \ALU.h_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48570\,
            in1 => \N__49122\,
            in2 => \_gnd_net_\,
            in3 => \N__49027\,
            lcout => \ALU.hZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47646\,
            ce => \N__45568\,
            sr => \_gnd_net_\
        );

    \ALU.a_13_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48565\,
            in1 => \N__33920\,
            in2 => \N__46201\,
            in3 => \N__33880\,
            lcout => \ALU.aZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47652\,
            ce => \N__44884\,
            sr => \_gnd_net_\
        );

    \ALU.a_14_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48574\,
            in1 => \N__33817\,
            in2 => \N__46200\,
            in3 => \N__33758\,
            lcout => \ALU.aZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47652\,
            ce => \N__44884\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48566\,
            in1 => \N__33662\,
            in2 => \N__46202\,
            in3 => \N__33603\,
            lcout => \ALU.aZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47652\,
            ce => \N__44884\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNI0P6L_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36623\,
            in1 => \_gnd_net_\,
            in2 => \N__35581\,
            in3 => \N__36467\,
            lcout => \ALU.f_RNI0P6LZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNICQEJ_1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36466\,
            in1 => \N__36622\,
            in2 => \_gnd_net_\,
            in3 => \N__32015\,
            lcout => \ALU.f_RNICQEJZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_RNIQCLL_7_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32014\,
            in1 => \N__31807\,
            in2 => \_gnd_net_\,
            in3 => \N__31690\,
            lcout => \ALU.g_RNIQCLLZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIL2FJ_5_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36433\,
            in1 => \N__48964\,
            in2 => \_gnd_net_\,
            in3 => \N__45103\,
            lcout => \ALU.f_RNIL2FJZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.m286_ns_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31646\,
            in1 => \N__33359\,
            in2 => \_gnd_net_\,
            in3 => \N__31628\,
            lcout => \N_287_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_2_rep1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34686\,
            in1 => \N__34769\,
            in2 => \N__32065\,
            in3 => \N__32228\,
            lcout => \aluOperand2_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIAOEJ_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35044\,
            in1 => \N__36286\,
            in2 => \_gnd_net_\,
            in3 => \N__32040\,
            lcout => \ALU.f_RNIAOEJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_fast_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34687\,
            in1 => \N__34770\,
            in2 => \N__31593\,
            in3 => \N__41114\,
            lcout => \aluOperand2_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_RNIESEJ_2_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32039\,
            in1 => \N__36451\,
            in2 => \_gnd_net_\,
            in3 => \N__31964\,
            lcout => \ALU.f_RNIESEJZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48622\,
            in1 => \N__42298\,
            in2 => \_gnd_net_\,
            in3 => \N__42265\,
            lcout => \ALU.gZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.g_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40999\,
            in1 => \N__48624\,
            in2 => \_gnd_net_\,
            in3 => \N__36592\,
            lcout => \ALU.gZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.g_2_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42161\,
            in1 => \N__48628\,
            in2 => \_gnd_net_\,
            in3 => \N__42097\,
            lcout => \ALU.gZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.g_3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48626\,
            in1 => \N__49469\,
            in2 => \_gnd_net_\,
            in3 => \N__49383\,
            lcout => \ALU.gZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.g_4_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48623\,
            in1 => \N__49288\,
            in2 => \_gnd_net_\,
            in3 => \N__49204\,
            lcout => \ALU.gZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.g_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48627\,
            in1 => \N__49123\,
            in2 => \_gnd_net_\,
            in3 => \N__49048\,
            lcout => \ALU.gZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.g_7_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48787\,
            in1 => \N__48625\,
            in2 => \_gnd_net_\,
            in3 => \N__48714\,
            lcout => \ALU.gZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47666\,
            ce => \N__36100\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJ17GT_15_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38735\,
            in1 => \N__31783\,
            in2 => \_gnd_net_\,
            in3 => \N__31772\,
            lcout => \ALU.N_634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_2_c_inv_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__32363\,
            in1 => \N__36517\,
            in2 => \_gnd_net_\,
            in3 => \N__32326\,
            lcout => \FTDI.un3_TX_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_12_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__32294\,
            in1 => \N__41467\,
            in2 => \N__32184\,
            in3 => \N__41220\,
            lcout => \testWordZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47605\,
            ce => \N__41063\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44754\,
            in1 => \N__44675\,
            in2 => \_gnd_net_\,
            in3 => \N__32153\,
            lcout => \FTDI.TXshiftZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_5_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__44612\,
            in2 => \_gnd_net_\,
            in3 => \N__44758\,
            lcout => \FTDI.TXshiftZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_3_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32120\,
            in1 => \N__32144\,
            in2 => \_gnd_net_\,
            in3 => \N__44756\,
            lcout => \FTDI.TXshiftZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44757\,
            in1 => \N__32135\,
            in2 => \_gnd_net_\,
            in3 => \N__32129\,
            lcout => \FTDI.TXshiftZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_2_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32111\,
            in1 => \N__32105\,
            in2 => \_gnd_net_\,
            in3 => \N__44755\,
            lcout => \FTDI.TXshiftZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44759\,
            in1 => \N__32558\,
            in2 => \_gnd_net_\,
            in3 => \N__32096\,
            lcout => \FTDI.TXshiftZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32567\,
            in2 => \_gnd_net_\,
            in3 => \N__44753\,
            lcout => \FTDI.TXshiftZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__44659\,
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_10_c_RNIEBKOT_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__42517\,
            in1 => \N__39212\,
            in2 => \_gnd_net_\,
            in3 => \N__32552\,
            lcout => \un2_addsub_cry_10_c_RNIEBKOT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_11_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__43754\,
            in1 => \N__47259\,
            in2 => \N__43939\,
            in3 => \N__44203\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI55HKC_11_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011110000110"
        )
    port map (
            in0 => \N__47260\,
            in1 => \N__39368\,
            in2 => \N__32537\,
            in3 => \N__39476\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIPTRDR1_11_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44204\,
            in2 => \N__32534\,
            in3 => \N__32531\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNID7K8N2_11_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46353\,
            in2 => \N__32516\,
            in3 => \N__32513\,
            lcout => OPEN,
            ltout => \c_RNID7K8N2_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNI5QD2L3_0_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48269\,
            in2 => \N__32501\,
            in3 => \N__32498\,
            lcout => \aluOperation_RNI5QD2L3_0\,
            ltout => \aluOperation_RNI5QD2L3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_11_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__48270\,
            in1 => \N__46040\,
            in2 => \N__32492\,
            in3 => \N__34181\,
            lcout => \ALU.aZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47611\,
            ce => \N__44872\,
            sr => \_gnd_net_\
        );

    \ALU.e_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000011111101"
        )
    port map (
            in0 => \N__45992\,
            in1 => \N__48328\,
            in2 => \N__36209\,
            in3 => \N__36258\,
            lcout => \ALU.eZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47615\,
            ce => \N__32435\,
            sr => \_gnd_net_\
        );

    \ALU.g_RNIVGLL_9_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36123\,
            in1 => \N__32715\,
            in2 => \_gnd_net_\,
            in3 => \N__45112\,
            lcout => OPEN,
            ltout => \ALU.g_RNIVGLLZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIURH32_9_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__33062\,
            in1 => \N__34475\,
            in2 => \N__32852\,
            in3 => \N__38345\,
            lcout => \ALU.operand2_7_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_m2_0_1_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__45321\,
            in1 => \N__38364\,
            in2 => \N__38401\,
            in3 => \N__35032\,
            lcout => \ALU.g0_0_0_m2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_m2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__32840\,
            in1 => \N__32796\,
            in2 => \N__32759\,
            in3 => \N__34474\,
            lcout => OPEN,
            ltout => \ALU.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_m4_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32684\,
            in1 => \_gnd_net_\,
            in2 => \N__32741\,
            in3 => \N__32970\,
            lcout => \ALU.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_0_m2_0_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__32716\,
            in1 => \N__34473\,
            in2 => \N__32693\,
            in3 => \N__36124\,
            lcout => \ALU.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_15_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100111111"
        )
    port map (
            in0 => \N__44205\,
            in1 => \N__43937\,
            in2 => \N__47321\,
            in3 => \N__43675\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIMPCHC_15_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011110000110"
        )
    port map (
            in0 => \N__47314\,
            in1 => \N__32674\,
            in2 => \N__32618\,
            in3 => \N__32615\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIM5JEB2_15_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__44206\,
            in1 => \_gnd_net_\,
            in2 => \N__32585\,
            in3 => \N__32582\,
            lcout => OPEN,
            ltout => \ALU.a_15_m4_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIR4QHM2_15_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46352\,
            in2 => \N__33521\,
            in3 => \N__33518\,
            lcout => OPEN,
            ltout => \ALU.c_RNIR4QHM2Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_14_c_RNI1G6N93_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48273\,
            in2 => \N__33506\,
            in3 => \N__40487\,
            lcout => \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93\,
            ltout => \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_15_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48274\,
            in1 => \N__45903\,
            in2 => \N__33503\,
            in3 => \N__33604\,
            lcout => \ALU.hZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47621\,
            ce => \N__45572\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNISBLU_15_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33487\,
            in1 => \N__33472\,
            in2 => \_gnd_net_\,
            in3 => \N__45299\,
            lcout => \ALU.d_RNISBLUZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperationZ0Z_5_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001001110"
        )
    port map (
            in0 => \N__33443\,
            in1 => \N__33163\,
            in2 => \N__33395\,
            in3 => \N__33354\,
            lcout => \aluOperation_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47628\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_1_l_ofx_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__37796\,
            in1 => \N__33149\,
            in2 => \N__37786\,
            in3 => \N__37479\,
            lcout => \ALU.madd_axb_1_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_0_rep2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34714\,
            in1 => \N__34796\,
            in2 => \N__41113\,
            in3 => \N__33048\,
            lcout => \aluOperand2_0_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47628\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__34794\,
            in1 => \N__34715\,
            in2 => \N__32959\,
            in3 => \N__41107\,
            lcout => \aluOperand2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47628\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIEFIJ_10_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__35029\,
            in1 => \N__34917\,
            in2 => \N__34269\,
            in3 => \N__34882\,
            lcout => \ALU.g0_7_m4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__34795\,
            in1 => \N__34716\,
            in2 => \N__34568\,
            in3 => \N__34488\,
            lcout => \aluOperand2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47628\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_10_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011101111"
        )
    port map (
            in0 => \N__48486\,
            in1 => \N__34403\,
            in2 => \N__46158\,
            in3 => \N__34342\,
            lcout => \ALU.gZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.g_11_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48490\,
            in1 => \N__34214\,
            in2 => \N__46000\,
            in3 => \N__34179\,
            lcout => \ALU.gZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.g_12_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48487\,
            in1 => \N__34091\,
            in2 => \N__46159\,
            in3 => \N__34025\,
            lcout => \ALU.gZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.g_13_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48491\,
            in1 => \N__33939\,
            in2 => \N__46001\,
            in3 => \N__33872\,
            lcout => \ALU.gZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.g_14_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48488\,
            in1 => \N__33818\,
            in2 => \N__46160\,
            in3 => \N__33748\,
            lcout => \ALU.gZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.g_15_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__48492\,
            in1 => \N__33653\,
            in2 => \N__46002\,
            in3 => \N__33605\,
            lcout => \ALU.gZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.g_9_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__48489\,
            in1 => \N__36264\,
            in2 => \N__46161\,
            in3 => \N__36195\,
            lcout => \ALU.gZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47635\,
            ce => \N__36093\,
            sr => \_gnd_net_\
        );

    \ALU.a_RNI85LF1_13_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__36038\,
            in1 => \N__36019\,
            in2 => \N__36003\,
            in3 => \N__35898\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFEHQ1_13_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__35810\,
            in1 => \N__35377\,
            in2 => \N__35798\,
            in3 => \N__35795\,
            lcout => \ALU.N_712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIRBBD1_13_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__35781\,
            in1 => \N__35752\,
            in2 => \N__35615\,
            in3 => \N__35532\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4TJ02_13_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__35462\,
            in1 => \N__35434\,
            in2 => \N__35405\,
            in3 => \N__35378\,
            lcout => OPEN,
            ltout => \ALU.N_760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINMUU3_13_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35252\,
            in2 => \N__35246\,
            in3 => \N__35229\,
            lcout => \ALU.aluOut_13\,
            ltout => \ALU.aluOut_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI7KNC7_13_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35072\,
            in3 => \N__38325\,
            lcout => \ALU.a13_b_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48493\,
            in1 => \N__42296\,
            in2 => \_gnd_net_\,
            in3 => \N__42266\,
            lcout => \ALU.fZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48582\,
            in1 => \N__40959\,
            in2 => \_gnd_net_\,
            in3 => \N__36591\,
            lcout => \ALU.fZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48494\,
            in1 => \N__42146\,
            in2 => \_gnd_net_\,
            in3 => \N__42096\,
            lcout => \ALU.fZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49361\,
            in1 => \N__48496\,
            in2 => \_gnd_net_\,
            in3 => \N__49442\,
            lcout => \ALU.fZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_4_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49212\,
            in1 => \N__48584\,
            in2 => \_gnd_net_\,
            in3 => \N__49262\,
            lcout => \ALU.fZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_5_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49090\,
            in1 => \N__48497\,
            in2 => \_gnd_net_\,
            in3 => \N__49043\,
            lcout => \ALU.fZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48495\,
            in1 => \N__48867\,
            in2 => \_gnd_net_\,
            in3 => \N__48931\,
            lcout => \ALU.fZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.f_7_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48583\,
            in1 => \N__48789\,
            in2 => \_gnd_net_\,
            in3 => \N__48696\,
            lcout => \ALU.fZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47647\,
            ce => \N__36380\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO75MA_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100110101001"
        )
    port map (
            in0 => \N__38037\,
            in1 => \N__36329\,
            in2 => \N__42526\,
            in3 => \N__38248\,
            lcout => \ALU.d_RNIO75MAZ0Z_0\,
            ltout => \ALU.d_RNIO75MAZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__48590\,
            in1 => \_gnd_net_\,
            in2 => \N__36302\,
            in3 => \N__42253\,
            lcout => \ALU.bZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => \N__47397\,
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_0_l_ofx_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__38249\,
            in1 => \N__38036\,
            in2 => \N__37502\,
            in3 => \N__37762\,
            lcout => \ALU.madd_axb_0_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__37763\,
            in1 => \N__37480\,
            in2 => \N__38047\,
            in3 => \N__38247\,
            lcout => OPEN,
            ltout => \ALU.mult_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEICQ63_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46004\,
            in2 => \N__36647\,
            in3 => \N__36644\,
            lcout => \ALU.d_RNIEICQ63Z0Z_1\,
            ltout => \ALU.d_RNIEICQ63Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48589\,
            in2 => \N__36626\,
            in3 => \N__40979\,
            lcout => \ALU.bZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47653\,
            ce => \N__47397\,
            sr => \_gnd_net_\
        );

    \ALU.d_1_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48591\,
            in1 => \N__40980\,
            in2 => \_gnd_net_\,
            in3 => \N__36590\,
            lcout => \ALU.dZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47659\,
            ce => \N__43344\,
            sr => \_gnd_net_\
        );

    \ALU.h_4_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__49213\,
            in1 => \N__48588\,
            in2 => \_gnd_net_\,
            in3 => \N__49289\,
            lcout => \ALU.hZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47673\,
            ce => \N__45573\,
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_2_c_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36518\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_2_0_\,
            carryout => \FTDI.un3_TX_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_3_c_inv_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36506\,
            in2 => \_gnd_net_\,
            in3 => \N__44771\,
            lcout => \FTDI.un3_TX_axb_3\,
            ltout => OPEN,
            carryin => \FTDI.un3_TX_cry_2\,
            carryout => \FTDI.un3_TX_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__44770\,
            in1 => \N__36500\,
            in2 => \_gnd_net_\,
            in3 => \N__36488\,
            lcout => \FTDI_TX_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIU2HCP_0_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38744\,
            in1 => \N__39199\,
            in2 => \_gnd_net_\,
            in3 => \N__39181\,
            lcout => \ALU.N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIMGKHG_13_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__39070\,
            in1 => \N__38765\,
            in2 => \N__38739\,
            in3 => \N__38444\,
            lcout => \ALU.rshift_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIR49H_9_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__38391\,
            in1 => \N__38371\,
            in2 => \N__45135\,
            in3 => \_gnd_net_\,
            lcout => \ALU.e_RNIR49HZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKQQR6_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38338\,
            in2 => \N__38051\,
            in3 => \N__37254\,
            lcout => \ALU.a0_b_2\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \ALU.un9_addsub_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_0_c_RNI2U096_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37787\,
            in2 => \N__37501\,
            in3 => \N__37259\,
            lcout => \ALU.un9_addsub_cry_0_c_RNI2UZ0Z096\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_0\,
            carryout => \ALU.un9_addsub_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_1_c_RNI6TD17_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37255\,
            in2 => \N__37001\,
            in3 => \N__36698\,
            lcout => \ALU.un9_addsub_cry_1_c_RNI6TDZ0Z17\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_1\,
            carryout => \ALU.un9_addsub_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_2_c_RNIA3LG7_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41974\,
            in2 => \N__36695\,
            in3 => \N__36680\,
            lcout => \ALU.un9_addsub_cry_2_c_RNIA3LGZ0Z7\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_2\,
            carryout => \ALU.un9_addsub_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_3_c_RNI525R7_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42992\,
            in2 => \N__36677\,
            in3 => \N__36665\,
            lcout => \ALU.un9_addsub_cry_3_c_RNI525RZ0Z7\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_3\,
            carryout => \ALU.un9_addsub_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_4_c_RNIL4N97_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40391\,
            in2 => \N__40223\,
            in3 => \N__40196\,
            lcout => \ALU.un9_addsub_cry_4_c_RNIL4NZ0Z97\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_4\,
            carryout => \ALU.un9_addsub_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_5_c_RNI6SCF7_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46733\,
            in2 => \N__40193\,
            in3 => \N__40175\,
            lcout => \ALU.un9_addsub_cry_5_c_RNI6SCFZ0Z7\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_5\,
            carryout => \ALU.un9_addsub_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_6_c_RNI2EFH8_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46976\,
            in2 => \N__40172\,
            in3 => \N__40124\,
            lcout => \ALU.un9_addsub_cry_6_c_RNI2EFHZ0Z8\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_6\,
            carryout => \ALU.un9_addsub_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_7_c_RNIU7F18_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40121\,
            in2 => \N__39890\,
            in3 => \N__39863\,
            lcout => \ALU.un9_addsub_cry_7_c_RNIU7FZ0Z18\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \ALU.un9_addsub_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_8_c_RNIPV1S8_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39859\,
            in2 => \N__39641\,
            in3 => \N__39611\,
            lcout => \ALU.un9_addsub_cry_8_c_RNIPV1SZ0Z8\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_8\,
            carryout => \ALU.un9_addsub_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_9_c_RNI22U6K_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39605\,
            in2 => \N__39506\,
            in3 => \N__39479\,
            lcout => \ALU.un9_addsub_cry_9_c_RNI22U6KZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_9\,
            carryout => \ALU.un9_addsub_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_10_c_RNI9C0K9_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39467\,
            in2 => \N__39398\,
            in3 => \N__39203\,
            lcout => \ALU.un9_addsub_cry_10_c_RNI9C0KZ0Z9\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_10\,
            carryout => \ALU.un9_addsub_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_11_c_RNI10BQK_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40853\,
            in2 => \N__40805\,
            in3 => \N__40775\,
            lcout => \ALU.un9_addsub_cry_11_c_RNI10BQKZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_11\,
            carryout => \ALU.un9_addsub_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_12_c_RNIBB5Q9_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40711\,
            in2 => \N__40664\,
            in3 => \N__40637\,
            lcout => \ALU.un9_addsub_cry_12_c_RNIBB5QZ0Z9\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_12\,
            carryout => \ALU.un9_addsub_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_13_c_RNI4JGF9_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40634\,
            in2 => \N__40559\,
            in3 => \N__40526\,
            lcout => \ALU.un9_addsub_cry_13_c_RNI4JGFZ0Z9\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_13\,
            carryout => \ALU.un9_addsub_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_14_c_RNIS374J_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__42495\,
            in1 => \N__40523\,
            in2 => \N__40508\,
            in3 => \N__40490\,
            lcout => \ALU.un9_addsub_cry_14_c_RNIS374JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_3_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__47303\,
            in1 => \N__44198\,
            in2 => \N__43952\,
            in3 => \N__43761\,
            lcout => \ALU.a_15_m2_ns_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJK5GK1_15_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44527\,
            in1 => \N__40481\,
            in2 => \_gnd_net_\,
            in3 => \N__40466\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3V2CP1_3_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__43185\,
            in1 => \_gnd_net_\,
            in2 => \N__40454\,
            in3 => \N__40451\,
            lcout => OPEN,
            ltout => \ALU.d_RNI3V2CP1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBRAVJ2_3_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46391\,
            in2 => \N__40436\,
            in3 => \N__41588\,
            lcout => \ALU.a_15_m5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJTNHA_3_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001100111"
        )
    port map (
            in0 => \N__47304\,
            in1 => \N__42005\,
            in2 => \N__41747\,
            in3 => \N__41735\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI95MLP_3_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__44526\,
            in1 => \N__44202\,
            in2 => \N__41609\,
            in3 => \N__41606\,
            lcout => \ALU.d_RNI95MLPZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIE8SJN5_3_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45893\,
            in1 => \N__41582\,
            in2 => \_gnd_net_\,
            in3 => \N__41573\,
            lcout => \ALU.d_RNIE8SJN5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testWord_10_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__41567\,
            in1 => \N__41500\,
            in2 => \N__41108\,
            in3 => \N__41231\,
            lcout => \testWordZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47629\,
            ce => \N__41061\,
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_0_c_RNIEMTLK_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42502\,
            in1 => \N__41021\,
            in2 => \_gnd_net_\,
            in3 => \N__41012\,
            lcout => \ALU.un9_addsub_cry_0_c_RNIEMTLKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_1_c_RNIM56UL_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42506\,
            in1 => \N__40925\,
            in2 => \_gnd_net_\,
            in3 => \N__40916\,
            lcout => \ALU.un9_addsub_cry_1_c_RNIM56ULZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_2_c_RNIMN63N_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40901\,
            in1 => \N__42507\,
            in2 => \_gnd_net_\,
            in3 => \N__40892\,
            lcout => \ALU.un9_addsub_cry_2_c_RNIMN63NZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_3_c_RNI4L7RO_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40877\,
            in1 => \N__42503\,
            in2 => \_gnd_net_\,
            in3 => \N__40862\,
            lcout => \ALU.un9_addsub_cry_3_c_RNI4L7ROZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_4_c_RNIUEDLM_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42504\,
            in1 => \N__42563\,
            in2 => \_gnd_net_\,
            in3 => \N__42554\,
            lcout => \ALU.un9_addsub_cry_4_c_RNIUEDLMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_5_c_RNI26HCN_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42539\,
            in1 => \N__42505\,
            in2 => \_gnd_net_\,
            in3 => \N__42419\,
            lcout => \ALU.un9_addsub_cry_5_c_RNI26HCNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_7_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__44226\,
            in1 => \N__47320\,
            in2 => \N__43963\,
            in3 => \N__43767\,
            lcout => \ALU.a_15_m2_ns_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIP43E91_7_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__42404\,
            in1 => \N__44537\,
            in2 => \N__46748\,
            in3 => \N__44227\,
            lcout => OPEN,
            ltout => \ALU.d_RNIP43E91Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIL4SQK2_7_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46393\,
            in1 => \_gnd_net_\,
            in2 => \N__42389\,
            in3 => \N__42386\,
            lcout => OPEN,
            ltout => \ALU.a_15_m5_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIIPM081_7_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__46003\,
            in1 => \N__42371\,
            in2 => \N__42356\,
            in3 => \N__42353\,
            lcout => \ALU.d_RNIIIPM081Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48578\,
            in1 => \N__42297\,
            in2 => \_gnd_net_\,
            in3 => \N__42264\,
            lcout => \ALU.dZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => \N__43340\,
            sr => \_gnd_net_\
        );

    \ALU.d_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48579\,
            in1 => \N__42126\,
            in2 => \_gnd_net_\,
            in3 => \N__42098\,
            lcout => \ALU.dZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => \N__43340\,
            sr => \_gnd_net_\
        );

    \ALU.d_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49441\,
            in1 => \N__48580\,
            in2 => \_gnd_net_\,
            in3 => \N__49360\,
            lcout => \ALU.dZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => \N__43340\,
            sr => \_gnd_net_\
        );

    \ALU.d_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48585\,
            in1 => \N__49044\,
            in2 => \_gnd_net_\,
            in3 => \N__49089\,
            lcout => \ALU.dZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => \N__43340\,
            sr => \_gnd_net_\
        );

    \ALU.d_6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48917\,
            in1 => \N__48587\,
            in2 => \_gnd_net_\,
            in3 => \N__48863\,
            lcout => \ALU.dZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => \N__43340\,
            sr => \_gnd_net_\
        );

    \ALU.d_7_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48586\,
            in1 => \N__48790\,
            in2 => \_gnd_net_\,
            in3 => \N__48684\,
            lcout => \ALU.dZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47641\,
            ce => \N__43340\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIHUEJ_3_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43261\,
            in1 => \N__49303\,
            in2 => \_gnd_net_\,
            in3 => \N__45119\,
            lcout => \ALU.f_RNIHUEJZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_4_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__47323\,
            in1 => \N__44224\,
            in2 => \N__43967\,
            in3 => \N__43768\,
            lcout => \ALU.a_15_m2_ns_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISSLDG1_6_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44540\,
            in1 => \N__43232\,
            in2 => \_gnd_net_\,
            in3 => \N__43211\,
            lcout => OPEN,
            ltout => \ALU.rshift_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC1CRK1_4_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43193\,
            in2 => \N__43025\,
            in3 => \N__43022\,
            lcout => OPEN,
            ltout => \ALU.a_15_m3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBK80K2_4_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46384\,
            in1 => \_gnd_net_\,
            in2 => \N__43001\,
            in3 => \N__44942\,
            lcout => \ALU.a_15_m5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINL83B_4_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001100111"
        )
    port map (
            in0 => \N__47324\,
            in1 => \N__42993\,
            in2 => \N__42707\,
            in3 => \N__42697\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0SA7U_4_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__44225\,
            in1 => \N__44539\,
            in2 => \N__44972\,
            in3 => \N__44969\,
            lcout => \ALU.a_15_m4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMA3938_4_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46085\,
            in1 => \N__44936\,
            in2 => \_gnd_net_\,
            in3 => \N__44921\,
            lcout => \ALU.d_RNIMA3938Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_3_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48577\,
            in1 => \N__49450\,
            in2 => \_gnd_net_\,
            in3 => \N__49378\,
            lcout => a_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47660\,
            ce => \N__44888\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_1_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44780\,
            in1 => \N__44567\,
            in2 => \_gnd_net_\,
            in3 => \N__44769\,
            lcout => \FTDI.TXshiftZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__44666\,
            sr => \_gnd_net_\
        );

    \TXbuffer_5_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44645\,
            lcout => \TXbufferZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47608\,
            ce => \N__44558\,
            sr => \_gnd_net_\
        );

    \TXbuffer_1_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44600\,
            lcout => \TXbufferZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47608\,
            ce => \N__44558\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJ75U41_6_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__44219\,
            in1 => \N__46400\,
            in2 => \N__44538\,
            in3 => \N__44240\,
            lcout => \ALU.d_RNIJ75U41Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_ns_1_6_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__47309\,
            in1 => \N__44223\,
            in2 => \N__43962\,
            in3 => \N__43763\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_ns_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMBENA_6_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001100111"
        )
    port map (
            in0 => \N__47310\,
            in1 => \N__46727\,
            in2 => \N__46484\,
            in3 => \N__46481\,
            lcout => \ALU.a_15_m2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7VNOJ2_6_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46392\,
            in1 => \N__46229\,
            in2 => \_gnd_net_\,
            in3 => \N__46208\,
            lcout => OPEN,
            ltout => \ALU.a_15_m5_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILPR7TQ_6_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46033\,
            in2 => \N__45638\,
            in3 => \N__45635\,
            lcout => \ALU.d_RNILPR7TQZ0Z_6\,
            ltout => \ALU.d_RNILPR7TQZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_6_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48509\,
            in2 => \N__45626\,
            in3 => \N__48856\,
            lcout => \ALU.hZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47616\,
            ce => \N__45557\,
            sr => \_gnd_net_\
        );

    \ALU.f_RNIJ0FJ_4_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45121\,
            in1 => \N__45409\,
            in2 => \_gnd_net_\,
            in3 => \N__49144\,
            lcout => \ALU.f_RNIJ0FJZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIU60L_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45373\,
            in1 => \N__45349\,
            in2 => \_gnd_net_\,
            in3 => \N__45312\,
            lcout => \ALU.d_RNIU60LZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILAR7_3_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45175\,
            in1 => \N__45148\,
            in2 => \_gnd_net_\,
            in3 => \N__45120\,
            lcout => \ALU.d_RNILAR7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48592\,
            in1 => \N__49443\,
            in2 => \_gnd_net_\,
            in3 => \N__49368\,
            lcout => \ALU.bZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47636\,
            ce => \N__47401\,
            sr => \_gnd_net_\
        );

    \ALU.b_4_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49244\,
            in1 => \N__48595\,
            in2 => \_gnd_net_\,
            in3 => \N__49211\,
            lcout => \ALU.bZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47636\,
            ce => \N__47401\,
            sr => \_gnd_net_\
        );

    \ALU.b_5_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48593\,
            in1 => \N__49094\,
            in2 => \_gnd_net_\,
            in3 => \N__49049\,
            lcout => \ALU.bZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47636\,
            ce => \N__47401\,
            sr => \_gnd_net_\
        );

    \ALU.b_6_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48916\,
            in1 => \N__48596\,
            in2 => \_gnd_net_\,
            in3 => \N__48880\,
            lcout => \ALU.bZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47636\,
            ce => \N__47401\,
            sr => \_gnd_net_\
        );

    \ALU.b_7_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48594\,
            in1 => \N__48791\,
            in2 => \_gnd_net_\,
            in3 => \N__48695\,
            lcout => \ALU.bZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47636\,
            ce => \N__47401\,
            sr => \_gnd_net_\
        );

    \ALU.b_8_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48581\,
            in1 => \N__47892\,
            in2 => \_gnd_net_\,
            in3 => \N__47810\,
            lcout => \ALU.bZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47636\,
            ce => \N__47401\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHRFPB_7_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010100101011"
        )
    port map (
            in0 => \N__47322\,
            in1 => \N__47105\,
            in2 => \N__46991\,
            in3 => \N__46964\,
            lcout => \ALU.a_15_m2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
