// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Aug 14 2020 14:01:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    RX,
    GPIO3,
    TX,
    GPIO2,
    GPIO11,
    GPIO0,
    CLK,
    GPIO9,
    GPIO1);

    input RX;
    output GPIO3;
    output TX;
    output GPIO2;
    output GPIO11;
    output GPIO0;
    input CLK;
    output GPIO9;
    output GPIO1;

    wire N__16292;
    wire N__16291;
    wire N__16290;
    wire N__16281;
    wire N__16280;
    wire N__16279;
    wire N__16272;
    wire N__16271;
    wire N__16270;
    wire N__16263;
    wire N__16262;
    wire N__16261;
    wire N__16254;
    wire N__16253;
    wire N__16252;
    wire N__16245;
    wire N__16244;
    wire N__16243;
    wire N__16236;
    wire N__16235;
    wire N__16234;
    wire N__16227;
    wire N__16226;
    wire N__16225;
    wire N__16218;
    wire N__16217;
    wire N__16216;
    wire N__16199;
    wire N__16196;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16188;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16175;
    wire N__16174;
    wire N__16173;
    wire N__16172;
    wire N__16169;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16148;
    wire N__16145;
    wire N__16140;
    wire N__16133;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16116;
    wire N__16115;
    wire N__16114;
    wire N__16113;
    wire N__16112;
    wire N__16111;
    wire N__16110;
    wire N__16109;
    wire N__16108;
    wire N__16107;
    wire N__16106;
    wire N__16105;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16101;
    wire N__16100;
    wire N__16099;
    wire N__16098;
    wire N__16097;
    wire N__16096;
    wire N__16095;
    wire N__16094;
    wire N__16093;
    wire N__16092;
    wire N__16091;
    wire N__16090;
    wire N__16089;
    wire N__16088;
    wire N__16087;
    wire N__16086;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16082;
    wire N__16081;
    wire N__16080;
    wire N__16079;
    wire N__16078;
    wire N__16077;
    wire N__16076;
    wire N__16075;
    wire N__16074;
    wire N__16073;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15914;
    wire N__15913;
    wire N__15912;
    wire N__15911;
    wire N__15910;
    wire N__15909;
    wire N__15908;
    wire N__15907;
    wire N__15906;
    wire N__15903;
    wire N__15902;
    wire N__15895;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15881;
    wire N__15880;
    wire N__15879;
    wire N__15876;
    wire N__15873;
    wire N__15872;
    wire N__15867;
    wire N__15864;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15850;
    wire N__15849;
    wire N__15844;
    wire N__15841;
    wire N__15836;
    wire N__15829;
    wire N__15828;
    wire N__15827;
    wire N__15826;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15806;
    wire N__15799;
    wire N__15796;
    wire N__15785;
    wire N__15784;
    wire N__15783;
    wire N__15782;
    wire N__15779;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15761;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15735;
    wire N__15734;
    wire N__15733;
    wire N__15732;
    wire N__15731;
    wire N__15724;
    wire N__15717;
    wire N__15710;
    wire N__15703;
    wire N__15700;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15680;
    wire N__15679;
    wire N__15678;
    wire N__15677;
    wire N__15676;
    wire N__15675;
    wire N__15674;
    wire N__15671;
    wire N__15666;
    wire N__15663;
    wire N__15662;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15651;
    wire N__15650;
    wire N__15647;
    wire N__15646;
    wire N__15645;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15612;
    wire N__15607;
    wire N__15606;
    wire N__15605;
    wire N__15602;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15585;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15574;
    wire N__15573;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15556;
    wire N__15553;
    wire N__15546;
    wire N__15539;
    wire N__15536;
    wire N__15529;
    wire N__15518;
    wire N__15517;
    wire N__15516;
    wire N__15515;
    wire N__15510;
    wire N__15505;
    wire N__15504;
    wire N__15503;
    wire N__15502;
    wire N__15501;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15493;
    wire N__15486;
    wire N__15483;
    wire N__15478;
    wire N__15475;
    wire N__15470;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15436;
    wire N__15435;
    wire N__15430;
    wire N__15429;
    wire N__15428;
    wire N__15427;
    wire N__15426;
    wire N__15425;
    wire N__15424;
    wire N__15423;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15390;
    wire N__15389;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15381;
    wire N__15378;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15353;
    wire N__15348;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15275;
    wire N__15274;
    wire N__15273;
    wire N__15270;
    wire N__15265;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15250;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15224;
    wire N__15217;
    wire N__15214;
    wire N__15209;
    wire N__15206;
    wire N__15205;
    wire N__15204;
    wire N__15201;
    wire N__15200;
    wire N__15199;
    wire N__15196;
    wire N__15195;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15188;
    wire N__15183;
    wire N__15182;
    wire N__15181;
    wire N__15180;
    wire N__15179;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15161;
    wire N__15160;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15143;
    wire N__15142;
    wire N__15139;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15135;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15110;
    wire N__15107;
    wire N__15100;
    wire N__15099;
    wire N__15088;
    wire N__15079;
    wire N__15076;
    wire N__15071;
    wire N__15060;
    wire N__15057;
    wire N__15052;
    wire N__15041;
    wire N__15040;
    wire N__15039;
    wire N__15038;
    wire N__15037;
    wire N__15036;
    wire N__15033;
    wire N__15032;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15024;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15006;
    wire N__15005;
    wire N__15002;
    wire N__15001;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14988;
    wire N__14987;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14962;
    wire N__14957;
    wire N__14950;
    wire N__14945;
    wire N__14942;
    wire N__14933;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14899;
    wire N__14898;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14890;
    wire N__14889;
    wire N__14888;
    wire N__14887;
    wire N__14886;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14878;
    wire N__14877;
    wire N__14876;
    wire N__14875;
    wire N__14874;
    wire N__14869;
    wire N__14868;
    wire N__14867;
    wire N__14866;
    wire N__14863;
    wire N__14862;
    wire N__14861;
    wire N__14860;
    wire N__14857;
    wire N__14848;
    wire N__14847;
    wire N__14842;
    wire N__14841;
    wire N__14840;
    wire N__14833;
    wire N__14832;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14821;
    wire N__14820;
    wire N__14819;
    wire N__14816;
    wire N__14811;
    wire N__14808;
    wire N__14801;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14785;
    wire N__14782;
    wire N__14777;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14747;
    wire N__14742;
    wire N__14741;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14729;
    wire N__14724;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14706;
    wire N__14701;
    wire N__14696;
    wire N__14689;
    wire N__14684;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14659;
    wire N__14658;
    wire N__14657;
    wire N__14656;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14648;
    wire N__14645;
    wire N__14644;
    wire N__14641;
    wire N__14636;
    wire N__14631;
    wire N__14628;
    wire N__14623;
    wire N__14622;
    wire N__14617;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14579;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14571;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14560;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14543;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14515;
    wire N__14514;
    wire N__14511;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14472;
    wire N__14465;
    wire N__14464;
    wire N__14463;
    wire N__14460;
    wire N__14459;
    wire N__14458;
    wire N__14457;
    wire N__14456;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14448;
    wire N__14447;
    wire N__14446;
    wire N__14445;
    wire N__14444;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14427;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14412;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14369;
    wire N__14368;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14352;
    wire N__14349;
    wire N__14346;
    wire N__14339;
    wire N__14334;
    wire N__14331;
    wire N__14318;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14297;
    wire N__14296;
    wire N__14293;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14277;
    wire N__14274;
    wire N__14267;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14256;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14244;
    wire N__14243;
    wire N__14240;
    wire N__14235;
    wire N__14232;
    wire N__14225;
    wire N__14224;
    wire N__14223;
    wire N__14220;
    wire N__14219;
    wire N__14216;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14172;
    wire N__14169;
    wire N__14162;
    wire N__14161;
    wire N__14158;
    wire N__14157;
    wire N__14154;
    wire N__14153;
    wire N__14150;
    wire N__14149;
    wire N__14148;
    wire N__14145;
    wire N__14142;
    wire N__14139;
    wire N__14136;
    wire N__14131;
    wire N__14130;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14113;
    wire N__14112;
    wire N__14109;
    wire N__14102;
    wire N__14099;
    wire N__14092;
    wire N__14089;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14020;
    wire N__14019;
    wire N__14018;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14003;
    wire N__13994;
    wire N__13993;
    wire N__13992;
    wire N__13985;
    wire N__13982;
    wire N__13981;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13969;
    wire N__13968;
    wire N__13961;
    wire N__13958;
    wire N__13957;
    wire N__13956;
    wire N__13953;
    wire N__13952;
    wire N__13951;
    wire N__13950;
    wire N__13947;
    wire N__13938;
    wire N__13933;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13906;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13880;
    wire N__13879;
    wire N__13878;
    wire N__13875;
    wire N__13874;
    wire N__13873;
    wire N__13870;
    wire N__13869;
    wire N__13868;
    wire N__13867;
    wire N__13866;
    wire N__13865;
    wire N__13864;
    wire N__13863;
    wire N__13860;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13836;
    wire N__13833;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13808;
    wire N__13795;
    wire N__13784;
    wire N__13783;
    wire N__13782;
    wire N__13781;
    wire N__13780;
    wire N__13777;
    wire N__13776;
    wire N__13773;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13768;
    wire N__13767;
    wire N__13766;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13745;
    wire N__13744;
    wire N__13741;
    wire N__13736;
    wire N__13729;
    wire N__13728;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13718;
    wire N__13717;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13705;
    wire N__13702;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13676;
    wire N__13675;
    wire N__13674;
    wire N__13673;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13669;
    wire N__13664;
    wire N__13657;
    wire N__13652;
    wire N__13645;
    wire N__13644;
    wire N__13643;
    wire N__13642;
    wire N__13639;
    wire N__13632;
    wire N__13627;
    wire N__13616;
    wire N__13611;
    wire N__13602;
    wire N__13597;
    wire N__13594;
    wire N__13587;
    wire N__13582;
    wire N__13579;
    wire N__13574;
    wire N__13567;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13537;
    wire N__13536;
    wire N__13535;
    wire N__13534;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13523;
    wire N__13522;
    wire N__13521;
    wire N__13520;
    wire N__13519;
    wire N__13516;
    wire N__13515;
    wire N__13514;
    wire N__13513;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13499;
    wire N__13496;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13466;
    wire N__13465;
    wire N__13464;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13441;
    wire N__13440;
    wire N__13439;
    wire N__13438;
    wire N__13437;
    wire N__13436;
    wire N__13435;
    wire N__13434;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13411;
    wire N__13404;
    wire N__13401;
    wire N__13390;
    wire N__13377;
    wire N__13374;
    wire N__13365;
    wire N__13346;
    wire N__13345;
    wire N__13344;
    wire N__13343;
    wire N__13342;
    wire N__13339;
    wire N__13338;
    wire N__13335;
    wire N__13334;
    wire N__13331;
    wire N__13326;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13318;
    wire N__13317;
    wire N__13316;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13299;
    wire N__13298;
    wire N__13297;
    wire N__13296;
    wire N__13291;
    wire N__13288;
    wire N__13287;
    wire N__13286;
    wire N__13285;
    wire N__13282;
    wire N__13277;
    wire N__13270;
    wire N__13265;
    wire N__13264;
    wire N__13261;
    wire N__13256;
    wire N__13253;
    wire N__13252;
    wire N__13247;
    wire N__13244;
    wire N__13239;
    wire N__13234;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13218;
    wire N__13215;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13183;
    wire N__13182;
    wire N__13179;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13160;
    wire N__13157;
    wire N__13156;
    wire N__13155;
    wire N__13154;
    wire N__13153;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13149;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13137;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13115;
    wire N__13108;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13086;
    wire N__13085;
    wire N__13082;
    wire N__13081;
    wire N__13080;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13056;
    wire N__13055;
    wire N__13054;
    wire N__13049;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13043;
    wire N__13040;
    wire N__13039;
    wire N__13036;
    wire N__13033;
    wire N__13032;
    wire N__13027;
    wire N__13024;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__12994;
    wire N__12989;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12951;
    wire N__12950;
    wire N__12949;
    wire N__12948;
    wire N__12947;
    wire N__12946;
    wire N__12945;
    wire N__12942;
    wire N__12941;
    wire N__12940;
    wire N__12939;
    wire N__12938;
    wire N__12935;
    wire N__12934;
    wire N__12931;
    wire N__12930;
    wire N__12929;
    wire N__12928;
    wire N__12927;
    wire N__12926;
    wire N__12921;
    wire N__12914;
    wire N__12899;
    wire N__12894;
    wire N__12889;
    wire N__12886;
    wire N__12875;
    wire N__12866;
    wire N__12857;
    wire N__12856;
    wire N__12853;
    wire N__12852;
    wire N__12851;
    wire N__12846;
    wire N__12845;
    wire N__12844;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12832;
    wire N__12831;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12802;
    wire N__12801;
    wire N__12798;
    wire N__12789;
    wire N__12786;
    wire N__12781;
    wire N__12772;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12741;
    wire N__12738;
    wire N__12733;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12713;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12641;
    wire N__12640;
    wire N__12639;
    wire N__12638;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12608;
    wire N__12607;
    wire N__12604;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12552;
    wire N__12547;
    wire N__12544;
    wire N__12539;
    wire N__12530;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12453;
    wire N__12450;
    wire N__12445;
    wire N__12444;
    wire N__12443;
    wire N__12442;
    wire N__12437;
    wire N__12434;
    wire N__12429;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12413;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12379;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12371;
    wire N__12370;
    wire N__12369;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12351;
    wire N__12348;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12332;
    wire N__12327;
    wire N__12324;
    wire N__12319;
    wire N__12314;
    wire N__12311;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12286;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12271;
    wire N__12268;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12245;
    wire N__12244;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12217;
    wire N__12214;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12176;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12077;
    wire N__12068;
    wire N__12067;
    wire N__12066;
    wire N__12065;
    wire N__12064;
    wire N__12063;
    wire N__12062;
    wire N__12061;
    wire N__12058;
    wire N__12057;
    wire N__12054;
    wire N__12053;
    wire N__12050;
    wire N__12049;
    wire N__12048;
    wire N__12045;
    wire N__12040;
    wire N__12037;
    wire N__12036;
    wire N__12035;
    wire N__12034;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12026;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12014;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12000;
    wire N__11995;
    wire N__11994;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11976;
    wire N__11971;
    wire N__11970;
    wire N__11969;
    wire N__11968;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11952;
    wire N__11949;
    wire N__11948;
    wire N__11947;
    wire N__11946;
    wire N__11945;
    wire N__11944;
    wire N__11941;
    wire N__11940;
    wire N__11933;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11915;
    wire N__11908;
    wire N__11905;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11887;
    wire N__11884;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11866;
    wire N__11859;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11831;
    wire N__11828;
    wire N__11827;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11803;
    wire N__11800;
    wire N__11799;
    wire N__11798;
    wire N__11797;
    wire N__11794;
    wire N__11789;
    wire N__11786;
    wire N__11785;
    wire N__11784;
    wire N__11783;
    wire N__11782;
    wire N__11781;
    wire N__11776;
    wire N__11771;
    wire N__11766;
    wire N__11763;
    wire N__11758;
    wire N__11753;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11746;
    wire N__11743;
    wire N__11738;
    wire N__11731;
    wire N__11730;
    wire N__11729;
    wire N__11724;
    wire N__11719;
    wire N__11716;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11700;
    wire N__11695;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11654;
    wire N__11653;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11647;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11630;
    wire N__11627;
    wire N__11620;
    wire N__11617;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11607;
    wire N__11606;
    wire N__11603;
    wire N__11602;
    wire N__11595;
    wire N__11592;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11555;
    wire N__11550;
    wire N__11547;
    wire N__11542;
    wire N__11535;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11512;
    wire N__11511;
    wire N__11510;
    wire N__11509;
    wire N__11498;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11485;
    wire N__11484;
    wire N__11481;
    wire N__11476;
    wire N__11461;
    wire N__11456;
    wire N__11453;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11449;
    wire N__11444;
    wire N__11437;
    wire N__11432;
    wire N__11431;
    wire N__11428;
    wire N__11423;
    wire N__11420;
    wire N__11419;
    wire N__11418;
    wire N__11417;
    wire N__11416;
    wire N__11415;
    wire N__11410;
    wire N__11401;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11349;
    wire N__11346;
    wire N__11341;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11321;
    wire N__11320;
    wire N__11315;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11294;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11278;
    wire N__11277;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11271;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11257;
    wire N__11254;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11231;
    wire N__11230;
    wire N__11223;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11203;
    wire N__11202;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11186;
    wire N__11181;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11107;
    wire N__11106;
    wire N__11105;
    wire N__11100;
    wire N__11099;
    wire N__11096;
    wire N__11095;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11053;
    wire N__11050;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10943;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10917;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10852;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10844;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10833;
    wire N__10830;
    wire N__10829;
    wire N__10828;
    wire N__10827;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10819;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10803;
    wire N__10800;
    wire N__10793;
    wire N__10786;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10500;
    wire N__10499;
    wire N__10496;
    wire N__10495;
    wire N__10492;
    wire N__10491;
    wire N__10488;
    wire N__10477;
    wire N__10472;
    wire N__10471;
    wire N__10470;
    wire N__10467;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10420;
    wire N__10419;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10395;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10291;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10271;
    wire N__10268;
    wire N__10263;
    wire N__10262;
    wire N__10259;
    wire N__10258;
    wire N__10255;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10237;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9803;
    wire N__9802;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9773;
    wire N__9770;
    wire N__9769;
    wire N__9764;
    wire N__9759;
    wire N__9750;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9595;
    wire N__9594;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9577;
    wire N__9574;
    wire N__9565;
    wire N__9558;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8746;
    wire N__8745;
    wire N__8744;
    wire N__8743;
    wire N__8740;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8723;
    wire N__8720;
    wire N__8719;
    wire N__8716;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8696;
    wire N__8693;
    wire N__8692;
    wire N__8691;
    wire N__8686;
    wire N__8683;
    wire N__8678;
    wire N__8675;
    wire N__8662;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8321;
    wire N__8318;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8258;
    wire N__8255;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8169;
    wire N__8168;
    wire N__8165;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7977;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7963;
    wire N__7962;
    wire N__7957;
    wire N__7954;
    wire N__7949;
    wire N__7946;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7931;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7896;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7882;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7878;
    wire N__7877;
    wire N__7870;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7855;
    wire N__7852;
    wire N__7851;
    wire N__7848;
    wire N__7843;
    wire N__7840;
    wire N__7829;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7789;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7768;
    wire N__7767;
    wire N__7764;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7758;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7747;
    wire N__7744;
    wire N__7743;
    wire N__7740;
    wire N__7739;
    wire N__7736;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7714;
    wire N__7701;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7450;
    wire N__7447;
    wire N__7446;
    wire N__7445;
    wire N__7442;
    wire N__7437;
    wire N__7436;
    wire N__7435;
    wire N__7432;
    wire N__7427;
    wire N__7422;
    wire N__7421;
    wire N__7420;
    wire N__7419;
    wire N__7416;
    wire N__7411;
    wire N__7404;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7362;
    wire N__7361;
    wire N__7358;
    wire N__7357;
    wire N__7354;
    wire N__7353;
    wire N__7350;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7334;
    wire N__7329;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7294;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7265;
    wire N__7262;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7105;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6825;
    wire N__6818;
    wire N__6815;
    wire N__6814;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6796;
    wire N__6793;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6781;
    wire N__6776;
    wire N__6775;
    wire N__6772;
    wire N__6771;
    wire N__6770;
    wire N__6769;
    wire N__6768;
    wire N__6765;
    wire N__6758;
    wire N__6753;
    wire N__6746;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6731;
    wire N__6730;
    wire N__6729;
    wire N__6728;
    wire N__6727;
    wire N__6726;
    wire N__6725;
    wire N__6714;
    wire N__6709;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6565;
    wire N__6564;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6113;
    wire GNDG0;
    wire VCCG0;
    wire clkdivZ0Z_0;
    wire bfn_1_13_0_;
    wire clkdivZ0Z_1;
    wire clkdiv_cry_0;
    wire clkdivZ0Z_2;
    wire clkdiv_cry_1;
    wire clkdivZ0Z_3;
    wire clkdiv_cry_2;
    wire clkdivZ0Z_4;
    wire clkdiv_cry_3;
    wire clkdivZ0Z_5;
    wire clkdiv_cry_4;
    wire clkdivZ0Z_6;
    wire clkdiv_cry_5;
    wire clkdivZ0Z_7;
    wire clkdiv_cry_6;
    wire clkdiv_cry_7;
    wire clkdivZ0Z_8;
    wire bfn_1_14_0_;
    wire clkdivZ0Z_9;
    wire clkdiv_cry_8;
    wire clkdivZ0Z_10;
    wire clkdiv_cry_9;
    wire clkdivZ0Z_11;
    wire clkdiv_cry_10;
    wire clkdivZ0Z_12;
    wire clkdiv_cry_11;
    wire clkdivZ0Z_13;
    wire clkdiv_cry_12;
    wire clkdivZ0Z_14;
    wire clkdiv_cry_13;
    wire clkdivZ0Z_15;
    wire clkdiv_cry_14;
    wire clkdiv_cry_15;
    wire clkdivZ0Z_16;
    wire bfn_1_15_0_;
    wire clkdivZ0Z_17;
    wire clkdiv_cry_16;
    wire clkdivZ0Z_18;
    wire clkdiv_cry_17;
    wire clkdivZ0Z_19;
    wire clkdiv_cry_18;
    wire clkdivZ0Z_20;
    wire clkdiv_cry_19;
    wire clkdivZ0Z_21;
    wire clkdiv_cry_20;
    wire clkdivZ0Z_22;
    wire clkdiv_cry_21;
    wire clkdiv_cry_22;
    wire GPIO3_c;
    wire \ALU.regsA_result_cry_1_0_c_RNO_2 ;
    wire bfn_9_11_0_;
    wire \ALU.regsA_result_cry_1 ;
    wire bfn_9_12_0_;
    wire \ALU.regsA_result_cry_4 ;
    wire \ALU.regsA_result_cry_5 ;
    wire \ALU.regsA_result_cry_6 ;
    wire \ALU.regsA_result_cry_7 ;
    wire \ALU.regsA_result_cry_4_c_RNO ;
    wire \ALU.regsA_result_cry_1_0_c_RNIKGQO9 ;
    wire \FTDI.i2_mux_cascade_ ;
    wire \FTDI.TXstate_RNIE1MMZ0Z_2 ;
    wire \FTDI.TXstate_RNIE1MMZ0Z_2_cascade_ ;
    wire \INVFTDI.TXstate_0C_net ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_1 ;
    wire bfn_10_10_0_;
    wire \ALU.regsA_result_cry_2_ma_1 ;
    wire \ALU.regsA_result_cry_1_5 ;
    wire \ALU.regsA_result_cry_3_ma_1 ;
    wire \ALU.regsA_result_cry_2_7 ;
    wire \ALU.regsA_result_cry_4_ma_0 ;
    wire \ALU.regsA_result_cry_3_7 ;
    wire \ALU.regsA_result_cry_4_6 ;
    wire \ALU.regsA_result_cry_5_0 ;
    wire \ALU.regsA_result_axb_4_l_ofx_0 ;
    wire \ALU.regsA_result_cry_5_ma_0 ;
    wire bfn_10_11_0_;
    wire \ALU.mult_AdderTree2_bigtree_704 ;
    wire \ALU.regsA_result_cry_2_0 ;
    wire \ALU.mult_AdderTree2_bigtree_705 ;
    wire \ALU.regsA_result_cry_3_4 ;
    wire \ALU.mult_AdderTree2_bigtree_706 ;
    wire \ALU.mult_AdderTree2_bigtree_871 ;
    wire \ALU.regsA_result_cry_4_3 ;
    wire \ALU.mult_AdderTree2_bigtree_707 ;
    wire \ALU.mult_AdderTree2_bigtree_872 ;
    wire \ALU.regsA_result_cry_5_4 ;
    wire \ALU.mult_AdderTree2_bigtree_708 ;
    wire \ALU.regsA_result_cry_6_3 ;
    wire \ALU.regsA_result_cry_7_1 ;
    wire \ALU.regsA_result_cry_2_c_RNO ;
    wire bfn_10_12_0_;
    wire \ALU.mult_AdderTree2_bigtree_873 ;
    wire \ALU.regsA_result_cry_2_c_RNIC59KA ;
    wire \ALU.regsA_result_cry_2 ;
    wire \ALU.regsA_result_cry_3_0 ;
    wire \ALU.regsA_result_cry_3_0_THRU_CO ;
    wire \ALU.mult_AdderTree2_bigtree_739 ;
    wire \ALU.mult_AdderTree2_bigtree_774 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_3 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO ;
    wire bfn_10_13_0_;
    wire \ALU.regsA_result_axb_2_l_ofx_0 ;
    wire \ALU.mult_AdderTree2_bigtree_740 ;
    wire \ALU.regsA_result_cry_1_4 ;
    wire \ALU.mult_AdderTree2_bigtree_741 ;
    wire \ALU.regsA_result_cry_2_6 ;
    wire \ALU.regsA_result_axb_2 ;
    wire \ALU.regsA_result_cry_1_THRU_CO ;
    wire \ALU.regsA_result_cry_3 ;
    wire \ALU.regsA_result_axb_4_0 ;
    wire \ALU.regsA_result_axb_3_l_ofx_0 ;
    wire \ALU.regsA_result_axb_4 ;
    wire \FTDI.baudAccZ0Z_0 ;
    wire \FTDI.baudAccZ0Z_1 ;
    wire \INVFTDI.baudAcc_0C_net ;
    wire \FTDI.N_170_0_cascade_ ;
    wire \FTDI.TXstate_cnst_0_0_2_cascade_ ;
    wire \INVFTDI.TXstate_2C_net ;
    wire \ALU.mult_AdderTree2_bigtree_870 ;
    wire \FTDI.TXstateZ0Z_1 ;
    wire \FTDI.TXstate_fastZ0Z_3 ;
    wire \FTDI.TXstateZ0Z_0 ;
    wire FTDI_TXready_cascade_;
    wire un1_testState31_0_cascade_;
    wire bfn_10_16_0_;
    wire \ALU.mult_AdderTree2_bigtree_669 ;
    wire \ALU.regsA_result_cry_0_0 ;
    wire \ALU.regsA_result_cry_5_c_RNI073QE ;
    wire \ALU.regsA_result_cry_1_1 ;
    wire \ALU.regsA_result_cry_2_c_RNIHNOEF ;
    wire \ALU.regsA_result_cry_2_2 ;
    wire \ALU.regsA_result_cry_7_c_RNI8EG3H ;
    wire \ALU.regsA_result_cry_3_2 ;
    wire \ALU.regsA_result_cry_4_c_RNIA939H ;
    wire \ALU.regsA_result_cry_4_1 ;
    wire \ALU.regsA_result_cry_5_c_RNIKCNNP ;
    wire \ALU.regsA_result_cry_5_2 ;
    wire \ALU.regsA_result_cry_6_c_RNICICNO ;
    wire \ALU.regsA_result_cry_6_1 ;
    wire \ALU.regsA_result_cry_7_9 ;
    wire bfn_10_17_0_;
    wire a_fastZ0Z_10;
    wire \ALU.regsA_result_axb_2_l_ofx_1 ;
    wire \ALU.regsA_result_axb_3_l_ofx_1 ;
    wire \ALU.regsA_result_axb_5_l_ofx_0 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_1 ;
    wire bfn_11_11_0_;
    wire \ALU.regsA_result_axb_2_l_ofx_2 ;
    wire \ALU.regsA_result_cry_1_6 ;
    wire \ALU.regsA_result_axb_3_l_ofx_2 ;
    wire \ALU.mult_AdderTree2_bigtree_671 ;
    wire \ALU.regsA_result_cry_2_8 ;
    wire \ALU.regsA_result_axb_4_l_ofx_1 ;
    wire \ALU.mult_AdderTree2_bigtree_672 ;
    wire \ALU.regsA_result_cry_3_8 ;
    wire \ALU.regsA_result_axb_5_l_ofx_1 ;
    wire \ALU.mult_AdderTree2_bigtree_673 ;
    wire \ALU.regsA_result_cry_4_7 ;
    wire \ALU.regsA_result_axb_6_l_ofx_0 ;
    wire \ALU.mult_AdderTree2_bigtree_674 ;
    wire \ALU.regsA_result_cry_5_7 ;
    wire \ALU.mult_AdderTree2_bigtree_675 ;
    wire \ALU.regsA_result_cry_6_6 ;
    wire \ALU.regsA_result_cry_5_0_THRU_CO ;
    wire \ALU.regsA_result_cry_7_0 ;
    wire \ALU.regsA_result_axb_8_2 ;
    wire \ALU.regsA_result_cry_6_ma_0 ;
    wire \ALU.mult_AdderTree2_bigtree_670 ;
    wire \ALU.regsA_result_cry_2_c_RNO_0 ;
    wire \ALU.regsA_result_cry_3_ma_0 ;
    wire \ALU.regsA_result_axb_6 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_0 ;
    wire bfn_11_14_0_;
    wire \ALU.addsub_cry_0_c_THRU_CO ;
    wire \ALU.addsub_cry_0 ;
    wire \ALU.addsub_axb_2_l_ofxZ0 ;
    wire \ALU.addsub_cry_1 ;
    wire \ALU.addsub_cry_2 ;
    wire \ALU.addsub_cry_3 ;
    wire \ALU.addsub_cry_4 ;
    wire \ALU.addsub_cry_5 ;
    wire \ALU.addsub_cry_6 ;
    wire bfn_11_15_0_;
    wire \ALU.addsub_cry_7 ;
    wire \ALU.addsub_cry_8 ;
    wire aZ0Z_10;
    wire \ALU.addsub_axb_10_l_ofxZ0 ;
    wire \ALU.addsub_cry_9 ;
    wire \ALU.addsub_cry_10 ;
    wire aZ0Z_12;
    wire \ALU.addsub_axb_12_l_ofxZ0 ;
    wire \ALU.addsub_cry_11 ;
    wire \ALU.addsub_cry_12 ;
    wire \ALU.addsub_cry_13 ;
    wire \ALU.addsub_cry_14 ;
    wire aZ0Z_15;
    wire \ALU.addsub_axb_15_l_ofxZ0 ;
    wire bfn_11_16_0_;
    wire \ALU.mult_16 ;
    wire \ALU.addsub_cry_15 ;
    wire \ALU.addsub_14 ;
    wire \ALU.mult_14 ;
    wire \ALU.mult_ab_128 ;
    wire \ALU.addsub_8 ;
    wire res_8;
    wire \ALU.addsub_11 ;
    wire \ALU.mult_11 ;
    wire \ALU.addsub_0 ;
    wire GPIO0_c;
    wire \ALU.addsub_13 ;
    wire \ALU.mult_13 ;
    wire \ALU.addsub_12 ;
    wire \ALU.mult_12 ;
    wire \ALU.mult_1 ;
    wire \ALU.addsub_1 ;
    wire \ALU.addsub_9 ;
    wire \ALU.mult_9 ;
    wire \ALU.addsub_10 ;
    wire \ALU.mult_10 ;
    wire \ALU.addsub_15 ;
    wire \ALU.mult_15 ;
    wire \ALU.addsub_6 ;
    wire \ALU.mult_2_cascade_ ;
    wire \ALU.addsub_2 ;
    wire \ALU.regsA_result_cry_7_ma_0 ;
    wire \ALU.regsA_result_axb_7_l_ofx_0 ;
    wire \ALU.regsA_result_axb_8_1 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_2 ;
    wire \ALU.regsA_result_cry_2_ma_2 ;
    wire \ALU.regsA_result_cry_3_ma_2 ;
    wire \ALU.regsA_result_cry_4_ma_1 ;
    wire aZ0Z_14;
    wire \ALU.addsub_axb_14_l_ofxZ0 ;
    wire aZ0Z_8;
    wire \ALU.addsub_axb_8_l_ofxZ0 ;
    wire \ALU.addsub_axb_9_l_ofxZ0 ;
    wire aZ0Z_9;
    wire \ALU.regsA_result_cry_5_ma_1 ;
    wire \ALU.regsA_result_cry_0_0_c_RNO ;
    wire bfn_12_12_0_;
    wire \ALU.regsA_result_axb_1_l_ofx ;
    wire \ALU.regsA_result_cry_0_2 ;
    wire \ALU.regsA_result_axb_2_l_ofx ;
    wire \ALU.regsA_result_cry_1_3 ;
    wire \ALU.regsA_result_cry_3_ma ;
    wire \ALU.regsA_result_axb_3_l_ofx ;
    wire \ALU.regsA_result_cry_2_5 ;
    wire \ALU.regsA_result_axb_4_l_ofx ;
    wire \ALU.regsA_result_cry_3_6 ;
    wire \ALU.regsA_result_axb_5_l_ofx ;
    wire \ALU.regsA_result_cry_4_5 ;
    wire \ALU.regsA_result_cry_5_6 ;
    wire \ALU.regsA_result_axb_7_l_ofx ;
    wire \ALU.regsA_result_cry_6_5 ;
    wire \ALU.regsA_result_cry_7_5 ;
    wire bfn_12_13_0_;
    wire \ALU.regsA_result_cry_8_2 ;
    wire \ALU.regsA_result_cry_9_3 ;
    wire \ALU.regsA_result_cry_10_2 ;
    wire \ALU.regsA_result_cry_11_3 ;
    wire \ALU.regsA_result_cry_12_0 ;
    wire \ALU.regsA_result_cry_13_1 ;
    wire \ALU.regsA_result_cry_14 ;
    wire \ALU.regsA_result_axb_14_l_ofx ;
    wire \ALU.addsub_axb_7_l_ofxZ0 ;
    wire \ALU.regsA_result_cry_8_ma ;
    wire \ALU.regsA_result_axb_14_0 ;
    wire \ALU.regsA_result_cry_14_ma ;
    wire \ALU.addsub_axb_1_l_ofxZ0 ;
    wire bZ0Z_15;
    wire \ALU.overflow_RNOZ0Z_15 ;
    wire \ALU.addsub_axb_0_l_ofxZ0 ;
    wire bfn_12_15_0_;
    wire \ALU.regsA_result_cry_0 ;
    wire \ALU.mult_6 ;
    wire \ALU.regsA_result_cry_1_0 ;
    wire \ALU.regsA_result_cry_2_1 ;
    wire \ALU.mult_AdderTree2_bigtree_932 ;
    wire \ALU.regsA_result_cry_3_1 ;
    wire \ALU.mult_AdderTree2_bigtree_933 ;
    wire \ALU.regsA_result_cry_4_0 ;
    wire \ALU.mult_AdderTree2_bigtree_934 ;
    wire \ALU.regsA_result_cry_5_1 ;
    wire \ALU.mult_AdderTree2_bigtree_935 ;
    wire \ALU.regsA_result_cry_6_0 ;
    wire \ALU.regsA_result_cry_7_2 ;
    wire \ALU.mult_AdderTree2_bigtree_936 ;
    wire bfn_12_16_0_;
    wire \ALU.mult_AdderTree2_bigtree_937 ;
    wire \ALU.regsA_result_cry_8 ;
    wire \ALU.mult_AdderTree2_bigtree_938 ;
    wire \ALU.regsA_result_cry_9_0 ;
    wire \ALU.mult_AdderTree2_bigtree_939 ;
    wire \ALU.regsA_result_cry_10 ;
    wire \ALU.regsA_result_axb_8 ;
    wire \ALU.regsA_result_cry_7_THRU_CO ;
    wire \ALU.regsA_result_cry_11_0 ;
    wire \ALU.regsA_result_axb_8_0 ;
    wire \ALU.mult_5 ;
    wire \ALU.addsub_5 ;
    wire \ALU.addsub_7 ;
    wire \ALU.mult_7 ;
    wire overflow;
    wire N_91;
    wire res_13;
    wire res_5;
    wire GPIO2_c;
    wire res_10;
    wire res_6;
    wire res_14;
    wire res_15;
    wire res_7;
    wire aZ0Z_11;
    wire \ALU.addsub_axb_11_l_ofxZ0 ;
    wire \ALU.regsA_result_axb_12_l_ofx ;
    wire \ALU.regsA_result_cry_11_ma ;
    wire \ALU.regsA_result_cry_12_ma ;
    wire \ALU.regsA_result_axb_13_l_ofx ;
    wire bfn_13_11_0_;
    wire \ALU.regsA_result_cry_1_8 ;
    wire \ALU.regsA_result_cry_2_10 ;
    wire \ALU.regsA_result_cry_3_10 ;
    wire \ALU.regsA_result_cry_5_ma_3 ;
    wire \ALU.regsA_result_cry_4_9 ;
    wire \ALU.regsA_result_cry_5_9 ;
    wire \ALU.regsA_result_cry_6_8 ;
    wire \ALU.regsA_result_cry_7_7 ;
    wire \ALU.regsA_result_cry_8_4 ;
    wire bfn_13_12_0_;
    wire \ALU.regsA_result_cry_9_5 ;
    wire \ALU.regsA_result_cry_10_4 ;
    wire \ALU.regsA_result_cry_11_4 ;
    wire \ALU.regsA_result_cry_13_ma_0 ;
    wire \ALU.regsA_result_axb_13_l_ofx_0 ;
    wire \ALU.regsA_result_cry_12_1 ;
    wire \ALU.regsA_result_cry_13_0 ;
    wire \ALU.regsA_result_cry_13_0_THRU_CO ;
    wire \ALU.regsA_result_cry_12_ma_0 ;
    wire \ALU.regsA_result_cry_0_0_c_RNO_0 ;
    wire bfn_13_13_0_;
    wire \ALU.mult_AdderTree2_bigtree_531 ;
    wire \ALU.regsA_result_cry_0_1 ;
    wire \ALU.mult_AdderTree2_bigtree_532 ;
    wire \ALU.mult_AdderTree2_bigtree_565 ;
    wire \ALU.regsA_result_cry_1_2 ;
    wire \ALU.mult_AdderTree2_bigtree_533 ;
    wire \ALU.mult_AdderTree2_bigtree_566 ;
    wire \ALU.mult_AdderTree2_bigtree_797 ;
    wire \ALU.regsA_result_cry_2_3 ;
    wire \ALU.mult_AdderTree2_bigtree_534 ;
    wire \ALU.mult_AdderTree2_bigtree_567 ;
    wire \ALU.mult_AdderTree2_bigtree_798 ;
    wire \ALU.regsA_result_cry_3_3 ;
    wire \ALU.mult_AdderTree2_bigtree_535 ;
    wire \ALU.mult_AdderTree2_bigtree_568 ;
    wire \ALU.mult_AdderTree2_bigtree_799 ;
    wire \ALU.regsA_result_cry_4_2 ;
    wire \ALU.mult_AdderTree2_bigtree_536 ;
    wire \ALU.mult_AdderTree2_bigtree_569 ;
    wire \ALU.mult_AdderTree2_bigtree_800 ;
    wire \ALU.regsA_result_cry_5_3 ;
    wire \ALU.mult_AdderTree2_bigtree_537 ;
    wire \ALU.mult_AdderTree2_bigtree_570 ;
    wire \ALU.mult_AdderTree2_bigtree_801 ;
    wire \ALU.regsA_result_cry_6_2 ;
    wire \ALU.regsA_result_cry_7_3 ;
    wire \ALU.mult_AdderTree2_bigtree_538 ;
    wire \ALU.mult_AdderTree2_bigtree_571 ;
    wire \ALU.mult_AdderTree2_bigtree_802 ;
    wire bfn_13_14_0_;
    wire \ALU.mult_AdderTree2_bigtree_539 ;
    wire \ALU.mult_AdderTree2_bigtree_572 ;
    wire \ALU.mult_AdderTree2_bigtree_803 ;
    wire \ALU.regsA_result_cry_8_0 ;
    wire \ALU.mult_AdderTree2_bigtree_540 ;
    wire \ALU.mult_AdderTree2_bigtree_573 ;
    wire \ALU.mult_AdderTree2_bigtree_804 ;
    wire \ALU.regsA_result_cry_9_1 ;
    wire \ALU.mult_AdderTree2_bigtree_541 ;
    wire \ALU.mult_AdderTree2_bigtree_574 ;
    wire \ALU.mult_AdderTree2_bigtree_805 ;
    wire \ALU.regsA_result_cry_10_0 ;
    wire \ALU.mult_AdderTree2_bigtree_542 ;
    wire \ALU.mult_AdderTree2_bigtree_575 ;
    wire \ALU.mult_AdderTree2_bigtree_806 ;
    wire \ALU.regsA_result_cry_11_2 ;
    wire \ALU.mult_AdderTree2_bigtree_543 ;
    wire \ALU.mult_AdderTree2_bigtree_576 ;
    wire \ALU.mult_AdderTree2_bigtree_807 ;
    wire \ALU.regsA_result_cry_12 ;
    wire \ALU.regsA_result_axb_14 ;
    wire \ALU.regsA_result_cry_13 ;
    wire \ALU.regsA_result_axb_12_0 ;
    wire bfn_13_15_0_;
    wire \ALU.mult_AdderTree2_bigtree_832 ;
    wire \ALU.regsA_result_cry_2_4 ;
    wire \ALU.mult_AdderTree2_bigtree_833 ;
    wire \ALU.regsA_result_cry_3_5 ;
    wire \ALU.mult_AdderTree2_bigtree_834 ;
    wire \ALU.regsA_result_cry_4_4 ;
    wire \ALU.mult_AdderTree2_bigtree_835 ;
    wire \ALU.regsA_result_cry_5_5 ;
    wire \ALU.mult_AdderTree2_bigtree_836 ;
    wire \ALU.regsA_result_cry_6_4 ;
    wire \ALU.mult_AdderTree2_bigtree_837 ;
    wire \ALU.regsA_result_cry_7_4 ;
    wire \ALU.mult_AdderTree2_bigtree_838 ;
    wire \ALU.regsA_result_cry_8_1 ;
    wire \ALU.regsA_result_cry_9_2 ;
    wire \ALU.mult_AdderTree2_bigtree_839 ;
    wire bfn_13_16_0_;
    wire \ALU.mult_AdderTree2_bigtree_840 ;
    wire \ALU.regsA_result_cry_10_1 ;
    wire \ALU.regsA_result_cry_11 ;
    wire \ALU.regsA_result_cry_11_THRU_CO ;
    wire \ALU.regsA_result_axb_10_l_ofx ;
    wire \ALU.addsub_3 ;
    wire \ALU.mult_3 ;
    wire res_11;
    wire res_3;
    wire GPIO1_c;
    wire res_9;
    wire res_12;
    wire TXstate_fast_RNIP6NA1_3;
    wire \ALU.regsA_result_axb_11_l_ofx ;
    wire \ALU.regsA_result_cry_10_ma ;
    wire \ALU.regsA_result_axb_11_l_ofx_1 ;
    wire bZ0Z_12;
    wire \ALU.regsA_result_axb_12_l_ofx_0 ;
    wire \ALU.regsA_result_axb_10_l_ofx_1 ;
    wire \ALU.regsA_result_cry_11_ma_1 ;
    wire \ALU.regsA_result_axb_2_l_ofx_4 ;
    wire \ALU.regsA_result_axb_3_l_ofx_4 ;
    wire \ALU.regsA_result_axb_4_l_ofx_3 ;
    wire \ALU.regsA_result_axb_5_l_ofx_3 ;
    wire \ALU.mult_AdderTree2_bigtree_564 ;
    wire a_fastZ0Z_2;
    wire \ALU.regsA_result_cry_1_0_c_RNO_4 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_5 ;
    wire \ALU.regsA_result_cry_2_ma_4 ;
    wire \ALU.regsA_result_cry_3_ma_4 ;
    wire \ALU.regsA_result_cry_4_ma_3 ;
    wire \ALU.mult_AdderTree2_bigtree_831 ;
    wire \ALU.mult_AdderTree2_bigtree_530 ;
    wire a_2_repZ0Z1;
    wire \ALU.regsA_result_cry_0_c_RNO_0 ;
    wire \ALU.regsA_result_cry_4_ma ;
    wire \ALU.regsA_result_cry_6_ma_2 ;
    wire \ALU.regsA_result_axb_6_l_ofx ;
    wire \ALU.regsA_result_cry_5_ma ;
    wire \ALU.regsA_result_axb_6_l_ofx_2 ;
    wire \ALU.regsA_result_cry_7_ma_2 ;
    wire \ALU.regsA_result_axb_7_l_ofx_2 ;
    wire \ALU.regsA_result_cry_6_ma ;
    wire \ALU.regsA_result_cry_8_ma_1 ;
    wire bfn_14_15_0_;
    wire \ALU.regsA_result_cry_1_7 ;
    wire \ALU.mult_AdderTree2_bigtree_601 ;
    wire \ALU.regsA_result_cry_2_9 ;
    wire \ALU.mult_AdderTree2_bigtree_602 ;
    wire \ALU.regsA_result_cry_3_9 ;
    wire \ALU.mult_AdderTree2_bigtree_603 ;
    wire \ALU.regsA_result_cry_4_8 ;
    wire \ALU.regsA_result_axb_6_l_ofx_1 ;
    wire \ALU.mult_AdderTree2_bigtree_604 ;
    wire \ALU.regsA_result_cry_5_8 ;
    wire \ALU.regsA_result_axb_7_l_ofx_1 ;
    wire \ALU.mult_AdderTree2_bigtree_605 ;
    wire \ALU.regsA_result_cry_6_7 ;
    wire \ALU.regsA_result_axb_8_l_ofx_0 ;
    wire \ALU.regsA_result_cry_8_ma_0 ;
    wire \ALU.mult_AdderTree2_bigtree_606 ;
    wire \ALU.regsA_result_cry_7_6 ;
    wire \ALU.regsA_result_cry_8_3 ;
    wire \ALU.mult_AdderTree2_bigtree_607 ;
    wire bfn_14_16_0_;
    wire \ALU.mult_AdderTree2_bigtree_608 ;
    wire \ALU.regsA_result_cry_9_4 ;
    wire \ALU.mult_AdderTree2_bigtree_609 ;
    wire \ALU.regsA_result_cry_10_3 ;
    wire \ALU.regsA_result_axb_12_1 ;
    wire \ALU.regsA_result_cry_11_1 ;
    wire \ALU.regsA_result_axb_12 ;
    wire \ALU.regsA_result_axb_10_l_ofx_0 ;
    wire \ALU.regsA_result_cry_11_ma_0 ;
    wire bZ0Z_11;
    wire \ALU.regsA_result_axb_11_l_ofx_0 ;
    wire \ALU.regsA_result_cry_10_ma_0 ;
    wire TXbufferZ0Z_1;
    wire TXbufferZ0Z_2;
    wire \FTDI.TXshiftZ0Z_2 ;
    wire TXbufferZ0Z_6;
    wire TXbufferZ0Z_4;
    wire \FTDI.TXshiftZ0Z_1 ;
    wire TXbufferZ0Z_0;
    wire \FTDI.TXshiftZ0Z_4 ;
    wire TXbufferZ0Z_3;
    wire \FTDI.TXshiftZ0Z_3 ;
    wire \FTDI.TXshiftZ0Z_6 ;
    wire TXbufferZ0Z_5;
    wire \FTDI.TXshiftZ0Z_5 ;
    wire \INVFTDI.TXshift_1C_net ;
    wire \INVFTDI.RXbuffer_2C_net ;
    wire \INVFTDI.RXbuffer_5C_net ;
    wire RXbuffer_3;
    wire \ALU.mult_AdderTree2_bigtree_599 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_3 ;
    wire \ALU.regsA_result_axb_2_l_ofx_3 ;
    wire \ALU.regsA_result_axb_3_l_ofx_3 ;
    wire \ALU.regsA_result_cry_0_c_RNO ;
    wire a_fastZ0Z_4;
    wire \ALU.mult_AdderTree2_bigtree_796 ;
    wire \ALU.mult_AdderTree2_bigtree_634 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_5 ;
    wire bfn_15_13_0_;
    wire \ALU.regsA_result_axb_2_l_ofx_5 ;
    wire \ALU.mult_AdderTree2_bigtree_635 ;
    wire \ALU.regsA_result_cry_1_9 ;
    wire \ALU.regsA_result_axb_3_l_ofx_5 ;
    wire \ALU.mult_AdderTree2_bigtree_636 ;
    wire \ALU.regsA_result_cry_2_11 ;
    wire \ALU.regsA_result_axb_4_l_ofx_4 ;
    wire \ALU.mult_AdderTree2_bigtree_637 ;
    wire \ALU.regsA_result_cry_3_11 ;
    wire \ALU.regsA_result_axb_5_l_ofx_4 ;
    wire \ALU.mult_AdderTree2_bigtree_638 ;
    wire \ALU.regsA_result_cry_4_10 ;
    wire \ALU.regsA_result_axb_6_l_ofx_3 ;
    wire \ALU.mult_AdderTree2_bigtree_639 ;
    wire \ALU.regsA_result_cry_5_10 ;
    wire \ALU.regsA_result_axb_7_l_ofx_3 ;
    wire \ALU.mult_AdderTree2_bigtree_640 ;
    wire \ALU.regsA_result_cry_6_9 ;
    wire \ALU.mult_AdderTree2_bigtree_641 ;
    wire \ALU.regsA_result_cry_7_8 ;
    wire \ALU.regsA_result_cry_8_5 ;
    wire \ALU.mult_AdderTree2_bigtree_642 ;
    wire bfn_15_14_0_;
    wire \ALU.regsA_result_cry_9 ;
    wire \ALU.regsA_result_cry_9_THRU_CO ;
    wire \ALU.regsA_result_cry_9_ma_0 ;
    wire \ALU.regsA_result_cry_2_ma_3 ;
    wire \ALU.regsA_result_cry_7_ma_1 ;
    wire \ALU.regsA_result_axb_10 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_4 ;
    wire \ALU.regsA_result_cry_1_0_c_RNO_0_6 ;
    wire \ALU.regsA_result_axb_4_l_ofx_2 ;
    wire RXbuffer_4;
    wire \ALU.regsA_result_axb_5_l_ofx_2 ;
    wire \ALU.addsub_axb_4_l_ofxZ0 ;
    wire \ALU.regsA_result_cry_4_ma_2 ;
    wire \ALU.regsA_result_cry_5_ma_2 ;
    wire \ALU.regsA_result_cry_6_ma_1 ;
    wire \ALU.regsA_result_axb_9_l_ofx ;
    wire aZ0Z_4;
    wire \ALU.regsA_result_axb_9_l_ofx_0 ;
    wire \ALU.regsA_result_cry_10_ma_1 ;
    wire RXbuffer_2;
    wire TXbufferZ0Z_7;
    wire \FTDI.TXshiftZ0Z_7 ;
    wire \INVFTDI.TXshift_7C_net ;
    wire RX_c;
    wire \FTDI.m13_ns_1_cascade_ ;
    wire \FTDI.N_201_2 ;
    wire \FTDI.N_23_cascade_ ;
    wire \FTDI.RXstateZ0Z_0 ;
    wire \INVFTDI.RXstate_3C_net ;
    wire \FTDI.RXstateZ0Z_3 ;
    wire \FTDI.RXstateZ0Z_2 ;
    wire \FTDI.N_28 ;
    wire \FTDI.RXstateZ0Z_1 ;
    wire \INVFTDI.RXstate_2C_net ;
    wire RXready_RNIICV7_0;
    wire RXbuffer_1;
    wire opZ0Z_1;
    wire \ALU.addsub_4 ;
    wire \ALU.mult_4 ;
    wire res_4;
    wire \ALU.regsA_result_cry_2_ma_0 ;
    wire RXbuffer_5;
    wire RXready_RNIICV7_1;
    wire \ALU.regsA_result_cry_1_ma ;
    wire \ALU.regsA_result_cry_3_ma_3 ;
    wire \ALU.regsA_result_cry_2_ma ;
    wire RXbuffer_7;
    wire bZ0Z_1;
    wire \ALU.regsA_result_cry_2_ma_5 ;
    wire bZ0Z_2;
    wire \ALU.regsA_result_cry_3_ma_5 ;
    wire \ALU.regsA_result_cry_4_ma_4 ;
    wire bZ0Z_4;
    wire \ALU.regsA_result_cry_5_ma_4 ;
    wire \ALU.regsA_result_cry_6_ma_3 ;
    wire aZ0Z_1;
    wire \ALU.regsA_result_axb_8_l_ofx ;
    wire \ALU.regsA_result_cry_7_ma ;
    wire \ALU.regsA_result_axb_8_l_ofx_1 ;
    wire \ALU.regsA_result_cry_9_ma_1 ;
    wire aZ0Z_2;
    wire \ALU.regsA_result_axb_9_l_ofx_1 ;
    wire \ALU.regsA_result_axb_8_l_ofx_2 ;
    wire bZ0Z_9;
    wire \ALU.regsA_result_axb_9_l_ofx_2 ;
    wire \ALU.addsub_axb_6_l_ofxZ0 ;
    wire \ALU.mult_AdderTree2_bigtree_600 ;
    wire aZ0Z_6;
    wire bZ0Z_0;
    wire \ALU.regsA_result_cry_2_c_RNO_1 ;
    wire aZ0Z_3;
    wire bZ0Z_3;
    wire \ALU.addsub_axb_3_l_ofxZ0 ;
    wire bZ0Z_8;
    wire \ALU.regsA_result_cry_9_ma_2 ;
    wire bZ0Z_6;
    wire \ALU.regsA_result_cry_7_ma_3 ;
    wire aZ0Z_7;
    wire bZ0Z_7;
    wire \ALU.regsA_result_cry_8_ma_2 ;
    wire \FTDI.baudAccZ0Z_2 ;
    wire \FTDI.un1_TXstate_0_sqmuxa_0_i ;
    wire TXstartZ0;
    wire un1_testState31_0_0;
    wire bZ0Z_10;
    wire \ALU.regsA_result_cry_9_ma ;
    wire CONSTANT_ONE_NET;
    wire \FTDI.un3_TX_0 ;
    wire \FTDI.gap8 ;
    wire \FTDI.gapZ0Z_1 ;
    wire \FTDI.gapZ0Z_0 ;
    wire \FTDI.gapZ0Z_2 ;
    wire \INVFTDI.gap_1C_net ;
    wire m7_x1;
    wire m7_x0_cascade_;
    wire RXready_RNIICV7_2;
    wire testState30_testState30_1_cascade_;
    wire aZ0Z_5;
    wire bZ0Z_5;
    wire \ALU.addsub_axb_5_l_ofxZ0 ;
    wire aZ0Z_0;
    wire \ALU.regsA_result_cry_13_ma ;
    wire aZ0Z_13;
    wire bZ0Z_13;
    wire \ALU.addsub_axb_13_l_ofxZ0 ;
    wire RXbuffer_0;
    wire opZ0Z_0;
    wire RXbuffer_6;
    wire bZ0Z_14;
    wire RXready_RNIICV7;
    wire i3_mux_i_x0_cascade_;
    wire FTDI_TXready;
    wire CLK_c_g;
    wire testState27;
    wire testStateZ0Z_0;
    wire testStateZ0Z_2;
    wire testStateZ0Z_1;
    wire RXready;
    wire i3_mux_i_x1;
    wire \FTDI.un3_TX_0_i ;
    wire bfn_17_16_0_;
    wire \FTDI.un3_TX_axb_3 ;
    wire \FTDI.un3_TX_cry_2 ;
    wire \FTDI.TXstateZ0Z_3 ;
    wire \FTDI.TXshiftZ0Z_0 ;
    wire \FTDI.un3_TX_cry_3 ;
    wire FTDI_TX_0_i;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__16290),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__16292),
            .DIN(N__16291),
            .DOUT(N__16290),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__16292),
            .PADOUT(N__16291),
            .PADIN(N__16290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO1_obuf_iopad (
            .OE(N__16281),
            .DIN(N__16280),
            .DOUT(N__16279),
            .PACKAGEPIN(GPIO1));
    defparam GPIO1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO1_obuf_preio (
            .PADOEN(N__16281),
            .PADOUT(N__16280),
            .PADIN(N__16279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9440),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO3_obuf_iopad (
            .OE(N__16272),
            .DIN(N__16271),
            .DOUT(N__16270),
            .PACKAGEPIN(GPIO3));
    defparam GPIO3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO3_obuf_preio (
            .PADOEN(N__16272),
            .PADOUT(N__16271),
            .PADIN(N__16270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6281),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO0_obuf_iopad (
            .OE(N__16263),
            .DIN(N__16262),
            .DOUT(N__16261),
            .PACKAGEPIN(GPIO0));
    defparam GPIO0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO0_obuf_preio (
            .PADOEN(N__16263),
            .PADOUT(N__16262),
            .PADIN(N__16261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7550),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO2_obuf_iopad (
            .OE(N__16254),
            .DIN(N__16253),
            .DOUT(N__16252),
            .PACKAGEPIN(GPIO2));
    defparam GPIO2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO2_obuf_preio (
            .PADOEN(N__16254),
            .PADOUT(N__16253),
            .PADIN(N__16252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8456),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RX_ibuf_iopad (
            .OE(N__16245),
            .DIN(N__16244),
            .DOUT(N__16243),
            .PACKAGEPIN(RX));
    defparam RX_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RX_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RX_ibuf_preio (
            .PADOEN(N__16245),
            .PADOUT(N__16244),
            .PADIN(N__16243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RX_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO11_obuf_iopad (
            .OE(N__16236),
            .DIN(N__16235),
            .DOUT(N__16234),
            .PACKAGEPIN(GPIO11));
    defparam GPIO11_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO11_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO11_obuf_preio (
            .PADOEN(N__16236),
            .PADOUT(N__16235),
            .PADIN(N__16234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TX_obuf_iopad (
            .OE(N__16227),
            .DIN(N__16226),
            .DOUT(N__16225),
            .PACKAGEPIN(TX));
    defparam TX_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TX_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TX_obuf_preio (
            .PADOEN(N__16227),
            .PADOUT(N__16226),
            .PADIN(N__16225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15326),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO9_obuf_iopad (
            .OE(N__16218),
            .DIN(N__16217),
            .DOUT(N__16216),
            .PACKAGEPIN(GPIO9));
    defparam GPIO9_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO9_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO9_obuf_preio (
            .PADOEN(N__16218),
            .PADOUT(N__16217),
            .PADIN(N__16216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14056),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__3892 (
            .O(N__16199),
            .I(i3_mux_i_x0_cascade_));
    InMux I__3891 (
            .O(N__16196),
            .I(N__16192));
    InMux I__3890 (
            .O(N__16195),
            .I(N__16189));
    LocalMux I__3889 (
            .O(N__16192),
            .I(N__16182));
    LocalMux I__3888 (
            .O(N__16189),
            .I(N__16179));
    InMux I__3887 (
            .O(N__16188),
            .I(N__16176));
    InMux I__3886 (
            .O(N__16187),
            .I(N__16169));
    InMux I__3885 (
            .O(N__16186),
            .I(N__16164));
    InMux I__3884 (
            .O(N__16185),
            .I(N__16164));
    Span4Mux_h I__3883 (
            .O(N__16182),
            .I(N__16161));
    Span4Mux_v I__3882 (
            .O(N__16179),
            .I(N__16158));
    LocalMux I__3881 (
            .O(N__16176),
            .I(N__16155));
    InMux I__3880 (
            .O(N__16175),
            .I(N__16148));
    InMux I__3879 (
            .O(N__16174),
            .I(N__16148));
    InMux I__3878 (
            .O(N__16173),
            .I(N__16148));
    InMux I__3877 (
            .O(N__16172),
            .I(N__16145));
    LocalMux I__3876 (
            .O(N__16169),
            .I(N__16140));
    LocalMux I__3875 (
            .O(N__16164),
            .I(N__16140));
    Span4Mux_v I__3874 (
            .O(N__16161),
            .I(N__16133));
    Span4Mux_h I__3873 (
            .O(N__16158),
            .I(N__16133));
    Span4Mux_v I__3872 (
            .O(N__16155),
            .I(N__16133));
    LocalMux I__3871 (
            .O(N__16148),
            .I(FTDI_TXready));
    LocalMux I__3870 (
            .O(N__16145),
            .I(FTDI_TXready));
    Odrv12 I__3869 (
            .O(N__16140),
            .I(FTDI_TXready));
    Odrv4 I__3868 (
            .O(N__16133),
            .I(FTDI_TXready));
    ClkMux I__3867 (
            .O(N__16124),
            .I(N__15968));
    ClkMux I__3866 (
            .O(N__16123),
            .I(N__15968));
    ClkMux I__3865 (
            .O(N__16122),
            .I(N__15968));
    ClkMux I__3864 (
            .O(N__16121),
            .I(N__15968));
    ClkMux I__3863 (
            .O(N__16120),
            .I(N__15968));
    ClkMux I__3862 (
            .O(N__16119),
            .I(N__15968));
    ClkMux I__3861 (
            .O(N__16118),
            .I(N__15968));
    ClkMux I__3860 (
            .O(N__16117),
            .I(N__15968));
    ClkMux I__3859 (
            .O(N__16116),
            .I(N__15968));
    ClkMux I__3858 (
            .O(N__16115),
            .I(N__15968));
    ClkMux I__3857 (
            .O(N__16114),
            .I(N__15968));
    ClkMux I__3856 (
            .O(N__16113),
            .I(N__15968));
    ClkMux I__3855 (
            .O(N__16112),
            .I(N__15968));
    ClkMux I__3854 (
            .O(N__16111),
            .I(N__15968));
    ClkMux I__3853 (
            .O(N__16110),
            .I(N__15968));
    ClkMux I__3852 (
            .O(N__16109),
            .I(N__15968));
    ClkMux I__3851 (
            .O(N__16108),
            .I(N__15968));
    ClkMux I__3850 (
            .O(N__16107),
            .I(N__15968));
    ClkMux I__3849 (
            .O(N__16106),
            .I(N__15968));
    ClkMux I__3848 (
            .O(N__16105),
            .I(N__15968));
    ClkMux I__3847 (
            .O(N__16104),
            .I(N__15968));
    ClkMux I__3846 (
            .O(N__16103),
            .I(N__15968));
    ClkMux I__3845 (
            .O(N__16102),
            .I(N__15968));
    ClkMux I__3844 (
            .O(N__16101),
            .I(N__15968));
    ClkMux I__3843 (
            .O(N__16100),
            .I(N__15968));
    ClkMux I__3842 (
            .O(N__16099),
            .I(N__15968));
    ClkMux I__3841 (
            .O(N__16098),
            .I(N__15968));
    ClkMux I__3840 (
            .O(N__16097),
            .I(N__15968));
    ClkMux I__3839 (
            .O(N__16096),
            .I(N__15968));
    ClkMux I__3838 (
            .O(N__16095),
            .I(N__15968));
    ClkMux I__3837 (
            .O(N__16094),
            .I(N__15968));
    ClkMux I__3836 (
            .O(N__16093),
            .I(N__15968));
    ClkMux I__3835 (
            .O(N__16092),
            .I(N__15968));
    ClkMux I__3834 (
            .O(N__16091),
            .I(N__15968));
    ClkMux I__3833 (
            .O(N__16090),
            .I(N__15968));
    ClkMux I__3832 (
            .O(N__16089),
            .I(N__15968));
    ClkMux I__3831 (
            .O(N__16088),
            .I(N__15968));
    ClkMux I__3830 (
            .O(N__16087),
            .I(N__15968));
    ClkMux I__3829 (
            .O(N__16086),
            .I(N__15968));
    ClkMux I__3828 (
            .O(N__16085),
            .I(N__15968));
    ClkMux I__3827 (
            .O(N__16084),
            .I(N__15968));
    ClkMux I__3826 (
            .O(N__16083),
            .I(N__15968));
    ClkMux I__3825 (
            .O(N__16082),
            .I(N__15968));
    ClkMux I__3824 (
            .O(N__16081),
            .I(N__15968));
    ClkMux I__3823 (
            .O(N__16080),
            .I(N__15968));
    ClkMux I__3822 (
            .O(N__16079),
            .I(N__15968));
    ClkMux I__3821 (
            .O(N__16078),
            .I(N__15968));
    ClkMux I__3820 (
            .O(N__16077),
            .I(N__15968));
    ClkMux I__3819 (
            .O(N__16076),
            .I(N__15968));
    ClkMux I__3818 (
            .O(N__16075),
            .I(N__15968));
    ClkMux I__3817 (
            .O(N__16074),
            .I(N__15968));
    ClkMux I__3816 (
            .O(N__16073),
            .I(N__15968));
    GlobalMux I__3815 (
            .O(N__15968),
            .I(N__15965));
    gio2CtrlBuf I__3814 (
            .O(N__15965),
            .I(CLK_c_g));
    CascadeMux I__3813 (
            .O(N__15962),
            .I(N__15958));
    SRMux I__3812 (
            .O(N__15961),
            .I(N__15955));
    InMux I__3811 (
            .O(N__15958),
            .I(N__15951));
    LocalMux I__3810 (
            .O(N__15955),
            .I(N__15948));
    InMux I__3809 (
            .O(N__15954),
            .I(N__15944));
    LocalMux I__3808 (
            .O(N__15951),
            .I(N__15941));
    Span4Mux_h I__3807 (
            .O(N__15948),
            .I(N__15938));
    InMux I__3806 (
            .O(N__15947),
            .I(N__15935));
    LocalMux I__3805 (
            .O(N__15944),
            .I(N__15932));
    Span4Mux_v I__3804 (
            .O(N__15941),
            .I(N__15929));
    Span4Mux_h I__3803 (
            .O(N__15938),
            .I(N__15926));
    LocalMux I__3802 (
            .O(N__15935),
            .I(N__15923));
    Odrv4 I__3801 (
            .O(N__15932),
            .I(testState27));
    Odrv4 I__3800 (
            .O(N__15929),
            .I(testState27));
    Odrv4 I__3799 (
            .O(N__15926),
            .I(testState27));
    Odrv12 I__3798 (
            .O(N__15923),
            .I(testState27));
    InMux I__3797 (
            .O(N__15914),
            .I(N__15903));
    InMux I__3796 (
            .O(N__15913),
            .I(N__15895));
    InMux I__3795 (
            .O(N__15912),
            .I(N__15895));
    InMux I__3794 (
            .O(N__15911),
            .I(N__15895));
    InMux I__3793 (
            .O(N__15910),
            .I(N__15884));
    InMux I__3792 (
            .O(N__15909),
            .I(N__15884));
    InMux I__3791 (
            .O(N__15908),
            .I(N__15884));
    InMux I__3790 (
            .O(N__15907),
            .I(N__15884));
    InMux I__3789 (
            .O(N__15906),
            .I(N__15884));
    LocalMux I__3788 (
            .O(N__15903),
            .I(N__15876));
    InMux I__3787 (
            .O(N__15902),
            .I(N__15873));
    LocalMux I__3786 (
            .O(N__15895),
            .I(N__15867));
    LocalMux I__3785 (
            .O(N__15884),
            .I(N__15867));
    InMux I__3784 (
            .O(N__15883),
            .I(N__15864));
    InMux I__3783 (
            .O(N__15882),
            .I(N__15861));
    InMux I__3782 (
            .O(N__15881),
            .I(N__15858));
    InMux I__3781 (
            .O(N__15880),
            .I(N__15855));
    CascadeMux I__3780 (
            .O(N__15879),
            .I(N__15850));
    Span4Mux_v I__3779 (
            .O(N__15876),
            .I(N__15844));
    LocalMux I__3778 (
            .O(N__15873),
            .I(N__15844));
    InMux I__3777 (
            .O(N__15872),
            .I(N__15841));
    Span4Mux_v I__3776 (
            .O(N__15867),
            .I(N__15836));
    LocalMux I__3775 (
            .O(N__15864),
            .I(N__15836));
    LocalMux I__3774 (
            .O(N__15861),
            .I(N__15829));
    LocalMux I__3773 (
            .O(N__15858),
            .I(N__15829));
    LocalMux I__3772 (
            .O(N__15855),
            .I(N__15829));
    InMux I__3771 (
            .O(N__15854),
            .I(N__15819));
    InMux I__3770 (
            .O(N__15853),
            .I(N__15819));
    InMux I__3769 (
            .O(N__15850),
            .I(N__15819));
    InMux I__3768 (
            .O(N__15849),
            .I(N__15816));
    Span4Mux_h I__3767 (
            .O(N__15844),
            .I(N__15813));
    LocalMux I__3766 (
            .O(N__15841),
            .I(N__15806));
    Span4Mux_h I__3765 (
            .O(N__15836),
            .I(N__15806));
    Span4Mux_v I__3764 (
            .O(N__15829),
            .I(N__15806));
    InMux I__3763 (
            .O(N__15828),
            .I(N__15799));
    InMux I__3762 (
            .O(N__15827),
            .I(N__15799));
    InMux I__3761 (
            .O(N__15826),
            .I(N__15799));
    LocalMux I__3760 (
            .O(N__15819),
            .I(N__15796));
    LocalMux I__3759 (
            .O(N__15816),
            .I(testStateZ0Z_0));
    Odrv4 I__3758 (
            .O(N__15813),
            .I(testStateZ0Z_0));
    Odrv4 I__3757 (
            .O(N__15806),
            .I(testStateZ0Z_0));
    LocalMux I__3756 (
            .O(N__15799),
            .I(testStateZ0Z_0));
    Odrv12 I__3755 (
            .O(N__15796),
            .I(testStateZ0Z_0));
    CascadeMux I__3754 (
            .O(N__15785),
            .I(N__15779));
    CascadeMux I__3753 (
            .O(N__15784),
            .I(N__15775));
    CascadeMux I__3752 (
            .O(N__15783),
            .I(N__15772));
    CascadeMux I__3751 (
            .O(N__15782),
            .I(N__15769));
    InMux I__3750 (
            .O(N__15779),
            .I(N__15765));
    InMux I__3749 (
            .O(N__15778),
            .I(N__15762));
    InMux I__3748 (
            .O(N__15775),
            .I(N__15757));
    InMux I__3747 (
            .O(N__15772),
            .I(N__15754));
    InMux I__3746 (
            .O(N__15769),
            .I(N__15751));
    InMux I__3745 (
            .O(N__15768),
            .I(N__15748));
    LocalMux I__3744 (
            .O(N__15765),
            .I(N__15745));
    LocalMux I__3743 (
            .O(N__15762),
            .I(N__15742));
    CascadeMux I__3742 (
            .O(N__15761),
            .I(N__15739));
    CascadeMux I__3741 (
            .O(N__15760),
            .I(N__15736));
    LocalMux I__3740 (
            .O(N__15757),
            .I(N__15724));
    LocalMux I__3739 (
            .O(N__15754),
            .I(N__15724));
    LocalMux I__3738 (
            .O(N__15751),
            .I(N__15724));
    LocalMux I__3737 (
            .O(N__15748),
            .I(N__15717));
    Span4Mux_v I__3736 (
            .O(N__15745),
            .I(N__15717));
    Span4Mux_h I__3735 (
            .O(N__15742),
            .I(N__15717));
    InMux I__3734 (
            .O(N__15739),
            .I(N__15710));
    InMux I__3733 (
            .O(N__15736),
            .I(N__15710));
    InMux I__3732 (
            .O(N__15735),
            .I(N__15710));
    InMux I__3731 (
            .O(N__15734),
            .I(N__15703));
    InMux I__3730 (
            .O(N__15733),
            .I(N__15703));
    InMux I__3729 (
            .O(N__15732),
            .I(N__15703));
    InMux I__3728 (
            .O(N__15731),
            .I(N__15700));
    Span4Mux_v I__3727 (
            .O(N__15724),
            .I(N__15695));
    Span4Mux_h I__3726 (
            .O(N__15717),
            .I(N__15695));
    LocalMux I__3725 (
            .O(N__15710),
            .I(N__15692));
    LocalMux I__3724 (
            .O(N__15703),
            .I(N__15689));
    LocalMux I__3723 (
            .O(N__15700),
            .I(testStateZ0Z_2));
    Odrv4 I__3722 (
            .O(N__15695),
            .I(testStateZ0Z_2));
    Odrv4 I__3721 (
            .O(N__15692),
            .I(testStateZ0Z_2));
    Odrv12 I__3720 (
            .O(N__15689),
            .I(testStateZ0Z_2));
    CascadeMux I__3719 (
            .O(N__15680),
            .I(N__15671));
    InMux I__3718 (
            .O(N__15679),
            .I(N__15666));
    InMux I__3717 (
            .O(N__15678),
            .I(N__15666));
    InMux I__3716 (
            .O(N__15677),
            .I(N__15663));
    CascadeMux I__3715 (
            .O(N__15676),
            .I(N__15658));
    CascadeMux I__3714 (
            .O(N__15675),
            .I(N__15655));
    CascadeMux I__3713 (
            .O(N__15674),
            .I(N__15652));
    InMux I__3712 (
            .O(N__15671),
            .I(N__15647));
    LocalMux I__3711 (
            .O(N__15666),
            .I(N__15640));
    LocalMux I__3710 (
            .O(N__15663),
            .I(N__15640));
    InMux I__3709 (
            .O(N__15662),
            .I(N__15637));
    InMux I__3708 (
            .O(N__15661),
            .I(N__15634));
    InMux I__3707 (
            .O(N__15658),
            .I(N__15625));
    InMux I__3706 (
            .O(N__15655),
            .I(N__15625));
    InMux I__3705 (
            .O(N__15652),
            .I(N__15625));
    InMux I__3704 (
            .O(N__15651),
            .I(N__15625));
    CascadeMux I__3703 (
            .O(N__15650),
            .I(N__15622));
    LocalMux I__3702 (
            .O(N__15647),
            .I(N__15619));
    CascadeMux I__3701 (
            .O(N__15646),
            .I(N__15616));
    CascadeMux I__3700 (
            .O(N__15645),
            .I(N__15613));
    Span4Mux_v I__3699 (
            .O(N__15640),
            .I(N__15607));
    LocalMux I__3698 (
            .O(N__15637),
            .I(N__15607));
    LocalMux I__3697 (
            .O(N__15634),
            .I(N__15602));
    LocalMux I__3696 (
            .O(N__15625),
            .I(N__15598));
    InMux I__3695 (
            .O(N__15622),
            .I(N__15595));
    Span4Mux_v I__3694 (
            .O(N__15619),
            .I(N__15592));
    InMux I__3693 (
            .O(N__15616),
            .I(N__15585));
    InMux I__3692 (
            .O(N__15613),
            .I(N__15585));
    InMux I__3691 (
            .O(N__15612),
            .I(N__15585));
    Span4Mux_v I__3690 (
            .O(N__15607),
            .I(N__15581));
    InMux I__3689 (
            .O(N__15606),
            .I(N__15578));
    InMux I__3688 (
            .O(N__15605),
            .I(N__15575));
    Span4Mux_v I__3687 (
            .O(N__15602),
            .I(N__15569));
    InMux I__3686 (
            .O(N__15601),
            .I(N__15566));
    Span4Mux_v I__3685 (
            .O(N__15598),
            .I(N__15563));
    LocalMux I__3684 (
            .O(N__15595),
            .I(N__15556));
    Span4Mux_h I__3683 (
            .O(N__15592),
            .I(N__15556));
    LocalMux I__3682 (
            .O(N__15585),
            .I(N__15556));
    InMux I__3681 (
            .O(N__15584),
            .I(N__15553));
    Span4Mux_h I__3680 (
            .O(N__15581),
            .I(N__15546));
    LocalMux I__3679 (
            .O(N__15578),
            .I(N__15546));
    LocalMux I__3678 (
            .O(N__15575),
            .I(N__15546));
    InMux I__3677 (
            .O(N__15574),
            .I(N__15539));
    InMux I__3676 (
            .O(N__15573),
            .I(N__15539));
    InMux I__3675 (
            .O(N__15572),
            .I(N__15539));
    Span4Mux_h I__3674 (
            .O(N__15569),
            .I(N__15536));
    LocalMux I__3673 (
            .O(N__15566),
            .I(N__15529));
    Span4Mux_h I__3672 (
            .O(N__15563),
            .I(N__15529));
    Span4Mux_v I__3671 (
            .O(N__15556),
            .I(N__15529));
    LocalMux I__3670 (
            .O(N__15553),
            .I(testStateZ0Z_1));
    Odrv4 I__3669 (
            .O(N__15546),
            .I(testStateZ0Z_1));
    LocalMux I__3668 (
            .O(N__15539),
            .I(testStateZ0Z_1));
    Odrv4 I__3667 (
            .O(N__15536),
            .I(testStateZ0Z_1));
    Odrv4 I__3666 (
            .O(N__15529),
            .I(testStateZ0Z_1));
    InMux I__3665 (
            .O(N__15518),
            .I(N__15510));
    InMux I__3664 (
            .O(N__15517),
            .I(N__15510));
    InMux I__3663 (
            .O(N__15516),
            .I(N__15505));
    InMux I__3662 (
            .O(N__15515),
            .I(N__15505));
    LocalMux I__3661 (
            .O(N__15510),
            .I(N__15493));
    LocalMux I__3660 (
            .O(N__15505),
            .I(N__15493));
    InMux I__3659 (
            .O(N__15504),
            .I(N__15486));
    InMux I__3658 (
            .O(N__15503),
            .I(N__15486));
    InMux I__3657 (
            .O(N__15502),
            .I(N__15486));
    InMux I__3656 (
            .O(N__15501),
            .I(N__15483));
    InMux I__3655 (
            .O(N__15500),
            .I(N__15478));
    InMux I__3654 (
            .O(N__15499),
            .I(N__15478));
    InMux I__3653 (
            .O(N__15498),
            .I(N__15475));
    Span4Mux_v I__3652 (
            .O(N__15493),
            .I(N__15470));
    LocalMux I__3651 (
            .O(N__15486),
            .I(N__15470));
    LocalMux I__3650 (
            .O(N__15483),
            .I(RXready));
    LocalMux I__3649 (
            .O(N__15478),
            .I(RXready));
    LocalMux I__3648 (
            .O(N__15475),
            .I(RXready));
    Odrv4 I__3647 (
            .O(N__15470),
            .I(RXready));
    InMux I__3646 (
            .O(N__15461),
            .I(N__15458));
    LocalMux I__3645 (
            .O(N__15458),
            .I(i3_mux_i_x1));
    InMux I__3644 (
            .O(N__15455),
            .I(N__15451));
    InMux I__3643 (
            .O(N__15454),
            .I(N__15448));
    LocalMux I__3642 (
            .O(N__15451),
            .I(\FTDI.un3_TX_0_i ));
    LocalMux I__3641 (
            .O(N__15448),
            .I(\FTDI.un3_TX_0_i ));
    InMux I__3640 (
            .O(N__15443),
            .I(N__15440));
    LocalMux I__3639 (
            .O(N__15440),
            .I(\FTDI.un3_TX_axb_3 ));
    InMux I__3638 (
            .O(N__15437),
            .I(N__15430));
    InMux I__3637 (
            .O(N__15436),
            .I(N__15430));
    CascadeMux I__3636 (
            .O(N__15435),
            .I(N__15419));
    LocalMux I__3635 (
            .O(N__15430),
            .I(N__15416));
    InMux I__3634 (
            .O(N__15429),
            .I(N__15401));
    InMux I__3633 (
            .O(N__15428),
            .I(N__15401));
    InMux I__3632 (
            .O(N__15427),
            .I(N__15401));
    InMux I__3631 (
            .O(N__15426),
            .I(N__15401));
    InMux I__3630 (
            .O(N__15425),
            .I(N__15401));
    InMux I__3629 (
            .O(N__15424),
            .I(N__15401));
    InMux I__3628 (
            .O(N__15423),
            .I(N__15401));
    InMux I__3627 (
            .O(N__15422),
            .I(N__15398));
    InMux I__3626 (
            .O(N__15419),
            .I(N__15395));
    Span4Mux_v I__3625 (
            .O(N__15416),
            .I(N__15390));
    LocalMux I__3624 (
            .O(N__15401),
            .I(N__15390));
    LocalMux I__3623 (
            .O(N__15398),
            .I(N__15385));
    LocalMux I__3622 (
            .O(N__15395),
            .I(N__15382));
    Span4Mux_h I__3621 (
            .O(N__15390),
            .I(N__15378));
    CascadeMux I__3620 (
            .O(N__15389),
            .I(N__15374));
    CascadeMux I__3619 (
            .O(N__15388),
            .I(N__15371));
    Span4Mux_v I__3618 (
            .O(N__15385),
            .I(N__15366));
    Span4Mux_h I__3617 (
            .O(N__15382),
            .I(N__15366));
    InMux I__3616 (
            .O(N__15381),
            .I(N__15363));
    Span4Mux_h I__3615 (
            .O(N__15378),
            .I(N__15360));
    InMux I__3614 (
            .O(N__15377),
            .I(N__15353));
    InMux I__3613 (
            .O(N__15374),
            .I(N__15353));
    InMux I__3612 (
            .O(N__15371),
            .I(N__15353));
    Span4Mux_h I__3611 (
            .O(N__15366),
            .I(N__15348));
    LocalMux I__3610 (
            .O(N__15363),
            .I(N__15348));
    Odrv4 I__3609 (
            .O(N__15360),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__3608 (
            .O(N__15353),
            .I(\FTDI.TXstateZ0Z_3 ));
    Odrv4 I__3607 (
            .O(N__15348),
            .I(\FTDI.TXstateZ0Z_3 ));
    InMux I__3606 (
            .O(N__15341),
            .I(N__15338));
    LocalMux I__3605 (
            .O(N__15338),
            .I(N__15335));
    Span4Mux_v I__3604 (
            .O(N__15335),
            .I(N__15332));
    Odrv4 I__3603 (
            .O(N__15332),
            .I(\FTDI.TXshiftZ0Z_0 ));
    InMux I__3602 (
            .O(N__15329),
            .I(\FTDI.un3_TX_cry_3 ));
    IoInMux I__3601 (
            .O(N__15326),
            .I(N__15323));
    LocalMux I__3600 (
            .O(N__15323),
            .I(N__15320));
    Span4Mux_s1_v I__3599 (
            .O(N__15320),
            .I(N__15317));
    Sp12to4 I__3598 (
            .O(N__15317),
            .I(N__15314));
    Span12Mux_h I__3597 (
            .O(N__15314),
            .I(N__15311));
    Span12Mux_v I__3596 (
            .O(N__15311),
            .I(N__15308));
    Odrv12 I__3595 (
            .O(N__15308),
            .I(FTDI_TX_0_i));
    InMux I__3594 (
            .O(N__15305),
            .I(N__15302));
    LocalMux I__3593 (
            .O(N__15302),
            .I(m7_x1));
    CascadeMux I__3592 (
            .O(N__15299),
            .I(m7_x0_cascade_));
    CEMux I__3591 (
            .O(N__15296),
            .I(N__15292));
    CEMux I__3590 (
            .O(N__15295),
            .I(N__15289));
    LocalMux I__3589 (
            .O(N__15292),
            .I(N__15286));
    LocalMux I__3588 (
            .O(N__15289),
            .I(N__15282));
    Span4Mux_v I__3587 (
            .O(N__15286),
            .I(N__15279));
    CEMux I__3586 (
            .O(N__15285),
            .I(N__15276));
    Span4Mux_v I__3585 (
            .O(N__15282),
            .I(N__15270));
    Span4Mux_v I__3584 (
            .O(N__15279),
            .I(N__15265));
    LocalMux I__3583 (
            .O(N__15276),
            .I(N__15265));
    CEMux I__3582 (
            .O(N__15275),
            .I(N__15261));
    CEMux I__3581 (
            .O(N__15274),
            .I(N__15258));
    CEMux I__3580 (
            .O(N__15273),
            .I(N__15255));
    Span4Mux_h I__3579 (
            .O(N__15270),
            .I(N__15250));
    Span4Mux_v I__3578 (
            .O(N__15265),
            .I(N__15250));
    CEMux I__3577 (
            .O(N__15264),
            .I(N__15246));
    LocalMux I__3576 (
            .O(N__15261),
            .I(N__15243));
    LocalMux I__3575 (
            .O(N__15258),
            .I(N__15238));
    LocalMux I__3574 (
            .O(N__15255),
            .I(N__15238));
    Span4Mux_h I__3573 (
            .O(N__15250),
            .I(N__15235));
    CEMux I__3572 (
            .O(N__15249),
            .I(N__15232));
    LocalMux I__3571 (
            .O(N__15246),
            .I(N__15229));
    Span4Mux_h I__3570 (
            .O(N__15243),
            .I(N__15224));
    Span4Mux_v I__3569 (
            .O(N__15238),
            .I(N__15224));
    Sp12to4 I__3568 (
            .O(N__15235),
            .I(N__15217));
    LocalMux I__3567 (
            .O(N__15232),
            .I(N__15217));
    Sp12to4 I__3566 (
            .O(N__15229),
            .I(N__15217));
    Span4Mux_h I__3565 (
            .O(N__15224),
            .I(N__15214));
    Odrv12 I__3564 (
            .O(N__15217),
            .I(RXready_RNIICV7_2));
    Odrv4 I__3563 (
            .O(N__15214),
            .I(RXready_RNIICV7_2));
    CascadeMux I__3562 (
            .O(N__15209),
            .I(testState30_testState30_1_cascade_));
    CascadeMux I__3561 (
            .O(N__15206),
            .I(N__15201));
    CascadeMux I__3560 (
            .O(N__15205),
            .I(N__15196));
    InMux I__3559 (
            .O(N__15204),
            .I(N__15192));
    InMux I__3558 (
            .O(N__15201),
            .I(N__15183));
    InMux I__3557 (
            .O(N__15200),
            .I(N__15183));
    InMux I__3556 (
            .O(N__15199),
            .I(N__15174));
    InMux I__3555 (
            .O(N__15196),
            .I(N__15174));
    InMux I__3554 (
            .O(N__15195),
            .I(N__15171));
    LocalMux I__3553 (
            .O(N__15192),
            .I(N__15168));
    InMux I__3552 (
            .O(N__15191),
            .I(N__15165));
    CascadeMux I__3551 (
            .O(N__15190),
            .I(N__15162));
    InMux I__3550 (
            .O(N__15189),
            .I(N__15156));
    InMux I__3549 (
            .O(N__15188),
            .I(N__15153));
    LocalMux I__3548 (
            .O(N__15183),
            .I(N__15150));
    InMux I__3547 (
            .O(N__15182),
            .I(N__15143));
    InMux I__3546 (
            .O(N__15181),
            .I(N__15143));
    InMux I__3545 (
            .O(N__15180),
            .I(N__15143));
    CascadeMux I__3544 (
            .O(N__15179),
            .I(N__15139));
    LocalMux I__3543 (
            .O(N__15174),
            .I(N__15129));
    LocalMux I__3542 (
            .O(N__15171),
            .I(N__15126));
    Span4Mux_v I__3541 (
            .O(N__15168),
            .I(N__15123));
    LocalMux I__3540 (
            .O(N__15165),
            .I(N__15120));
    InMux I__3539 (
            .O(N__15162),
            .I(N__15117));
    InMux I__3538 (
            .O(N__15161),
            .I(N__15110));
    InMux I__3537 (
            .O(N__15160),
            .I(N__15110));
    InMux I__3536 (
            .O(N__15159),
            .I(N__15110));
    LocalMux I__3535 (
            .O(N__15156),
            .I(N__15107));
    LocalMux I__3534 (
            .O(N__15153),
            .I(N__15100));
    Span4Mux_v I__3533 (
            .O(N__15150),
            .I(N__15100));
    LocalMux I__3532 (
            .O(N__15143),
            .I(N__15100));
    InMux I__3531 (
            .O(N__15142),
            .I(N__15088));
    InMux I__3530 (
            .O(N__15139),
            .I(N__15088));
    InMux I__3529 (
            .O(N__15138),
            .I(N__15088));
    InMux I__3528 (
            .O(N__15137),
            .I(N__15088));
    InMux I__3527 (
            .O(N__15136),
            .I(N__15088));
    InMux I__3526 (
            .O(N__15135),
            .I(N__15079));
    InMux I__3525 (
            .O(N__15134),
            .I(N__15079));
    InMux I__3524 (
            .O(N__15133),
            .I(N__15079));
    InMux I__3523 (
            .O(N__15132),
            .I(N__15079));
    Span4Mux_v I__3522 (
            .O(N__15129),
            .I(N__15076));
    Span4Mux_v I__3521 (
            .O(N__15126),
            .I(N__15071));
    Span4Mux_h I__3520 (
            .O(N__15123),
            .I(N__15071));
    Span4Mux_v I__3519 (
            .O(N__15120),
            .I(N__15060));
    LocalMux I__3518 (
            .O(N__15117),
            .I(N__15060));
    LocalMux I__3517 (
            .O(N__15110),
            .I(N__15060));
    Span4Mux_v I__3516 (
            .O(N__15107),
            .I(N__15060));
    Span4Mux_v I__3515 (
            .O(N__15100),
            .I(N__15060));
    InMux I__3514 (
            .O(N__15099),
            .I(N__15057));
    LocalMux I__3513 (
            .O(N__15088),
            .I(N__15052));
    LocalMux I__3512 (
            .O(N__15079),
            .I(N__15052));
    Odrv4 I__3511 (
            .O(N__15076),
            .I(aZ0Z_5));
    Odrv4 I__3510 (
            .O(N__15071),
            .I(aZ0Z_5));
    Odrv4 I__3509 (
            .O(N__15060),
            .I(aZ0Z_5));
    LocalMux I__3508 (
            .O(N__15057),
            .I(aZ0Z_5));
    Odrv12 I__3507 (
            .O(N__15052),
            .I(aZ0Z_5));
    CascadeMux I__3506 (
            .O(N__15041),
            .I(N__15033));
    InMux I__3505 (
            .O(N__15040),
            .I(N__15028));
    InMux I__3504 (
            .O(N__15039),
            .I(N__15025));
    InMux I__3503 (
            .O(N__15038),
            .I(N__15019));
    InMux I__3502 (
            .O(N__15037),
            .I(N__15019));
    InMux I__3501 (
            .O(N__15036),
            .I(N__15014));
    InMux I__3500 (
            .O(N__15033),
            .I(N__15011));
    InMux I__3499 (
            .O(N__15032),
            .I(N__15006));
    InMux I__3498 (
            .O(N__15031),
            .I(N__15006));
    LocalMux I__3497 (
            .O(N__15028),
            .I(N__15002));
    LocalMux I__3496 (
            .O(N__15025),
            .I(N__14995));
    InMux I__3495 (
            .O(N__15024),
            .I(N__14992));
    LocalMux I__3494 (
            .O(N__15019),
            .I(N__14989));
    InMux I__3493 (
            .O(N__15018),
            .I(N__14982));
    InMux I__3492 (
            .O(N__15017),
            .I(N__14982));
    LocalMux I__3491 (
            .O(N__15014),
            .I(N__14979));
    LocalMux I__3490 (
            .O(N__15011),
            .I(N__14976));
    LocalMux I__3489 (
            .O(N__15006),
            .I(N__14973));
    InMux I__3488 (
            .O(N__15005),
            .I(N__14970));
    Span4Mux_v I__3487 (
            .O(N__15002),
            .I(N__14967));
    InMux I__3486 (
            .O(N__15001),
            .I(N__14962));
    InMux I__3485 (
            .O(N__15000),
            .I(N__14962));
    InMux I__3484 (
            .O(N__14999),
            .I(N__14957));
    InMux I__3483 (
            .O(N__14998),
            .I(N__14957));
    Span4Mux_h I__3482 (
            .O(N__14995),
            .I(N__14950));
    LocalMux I__3481 (
            .O(N__14992),
            .I(N__14950));
    Span4Mux_h I__3480 (
            .O(N__14989),
            .I(N__14950));
    InMux I__3479 (
            .O(N__14988),
            .I(N__14945));
    InMux I__3478 (
            .O(N__14987),
            .I(N__14945));
    LocalMux I__3477 (
            .O(N__14982),
            .I(N__14942));
    Span4Mux_v I__3476 (
            .O(N__14979),
            .I(N__14933));
    Span4Mux_h I__3475 (
            .O(N__14976),
            .I(N__14933));
    Span4Mux_h I__3474 (
            .O(N__14973),
            .I(N__14933));
    LocalMux I__3473 (
            .O(N__14970),
            .I(N__14933));
    Odrv4 I__3472 (
            .O(N__14967),
            .I(bZ0Z_5));
    LocalMux I__3471 (
            .O(N__14962),
            .I(bZ0Z_5));
    LocalMux I__3470 (
            .O(N__14957),
            .I(bZ0Z_5));
    Odrv4 I__3469 (
            .O(N__14950),
            .I(bZ0Z_5));
    LocalMux I__3468 (
            .O(N__14945),
            .I(bZ0Z_5));
    Odrv4 I__3467 (
            .O(N__14942),
            .I(bZ0Z_5));
    Odrv4 I__3466 (
            .O(N__14933),
            .I(bZ0Z_5));
    CascadeMux I__3465 (
            .O(N__14918),
            .I(N__14915));
    InMux I__3464 (
            .O(N__14915),
            .I(N__14912));
    LocalMux I__3463 (
            .O(N__14912),
            .I(N__14909));
    Span4Mux_h I__3462 (
            .O(N__14909),
            .I(N__14906));
    Span4Mux_h I__3461 (
            .O(N__14906),
            .I(N__14903));
    Odrv4 I__3460 (
            .O(N__14903),
            .I(\ALU.addsub_axb_5_l_ofxZ0 ));
    CascadeMux I__3459 (
            .O(N__14900),
            .I(N__14894));
    CascadeMux I__3458 (
            .O(N__14899),
            .I(N__14891));
    CascadeMux I__3457 (
            .O(N__14898),
            .I(N__14882));
    CascadeMux I__3456 (
            .O(N__14897),
            .I(N__14879));
    InMux I__3455 (
            .O(N__14894),
            .I(N__14869));
    InMux I__3454 (
            .O(N__14891),
            .I(N__14869));
    InMux I__3453 (
            .O(N__14890),
            .I(N__14863));
    InMux I__3452 (
            .O(N__14889),
            .I(N__14857));
    InMux I__3451 (
            .O(N__14888),
            .I(N__14848));
    InMux I__3450 (
            .O(N__14887),
            .I(N__14848));
    InMux I__3449 (
            .O(N__14886),
            .I(N__14848));
    InMux I__3448 (
            .O(N__14885),
            .I(N__14848));
    InMux I__3447 (
            .O(N__14882),
            .I(N__14842));
    InMux I__3446 (
            .O(N__14879),
            .I(N__14842));
    InMux I__3445 (
            .O(N__14878),
            .I(N__14833));
    InMux I__3444 (
            .O(N__14877),
            .I(N__14833));
    InMux I__3443 (
            .O(N__14876),
            .I(N__14833));
    InMux I__3442 (
            .O(N__14875),
            .I(N__14828));
    InMux I__3441 (
            .O(N__14874),
            .I(N__14825));
    LocalMux I__3440 (
            .O(N__14869),
            .I(N__14822));
    InMux I__3439 (
            .O(N__14868),
            .I(N__14816));
    InMux I__3438 (
            .O(N__14867),
            .I(N__14811));
    InMux I__3437 (
            .O(N__14866),
            .I(N__14811));
    LocalMux I__3436 (
            .O(N__14863),
            .I(N__14808));
    InMux I__3435 (
            .O(N__14862),
            .I(N__14801));
    InMux I__3434 (
            .O(N__14861),
            .I(N__14801));
    InMux I__3433 (
            .O(N__14860),
            .I(N__14801));
    LocalMux I__3432 (
            .O(N__14857),
            .I(N__14796));
    LocalMux I__3431 (
            .O(N__14848),
            .I(N__14796));
    InMux I__3430 (
            .O(N__14847),
            .I(N__14793));
    LocalMux I__3429 (
            .O(N__14842),
            .I(N__14790));
    InMux I__3428 (
            .O(N__14841),
            .I(N__14785));
    InMux I__3427 (
            .O(N__14840),
            .I(N__14785));
    LocalMux I__3426 (
            .O(N__14833),
            .I(N__14782));
    InMux I__3425 (
            .O(N__14832),
            .I(N__14777));
    InMux I__3424 (
            .O(N__14831),
            .I(N__14777));
    LocalMux I__3423 (
            .O(N__14828),
            .I(N__14770));
    LocalMux I__3422 (
            .O(N__14825),
            .I(N__14770));
    Span4Mux_h I__3421 (
            .O(N__14822),
            .I(N__14770));
    InMux I__3420 (
            .O(N__14821),
            .I(N__14767));
    InMux I__3419 (
            .O(N__14820),
            .I(N__14764));
    InMux I__3418 (
            .O(N__14819),
            .I(N__14761));
    LocalMux I__3417 (
            .O(N__14816),
            .I(N__14758));
    LocalMux I__3416 (
            .O(N__14811),
            .I(N__14755));
    Span4Mux_v I__3415 (
            .O(N__14808),
            .I(N__14747));
    LocalMux I__3414 (
            .O(N__14801),
            .I(N__14747));
    Span4Mux_h I__3413 (
            .O(N__14796),
            .I(N__14742));
    LocalMux I__3412 (
            .O(N__14793),
            .I(N__14742));
    Span4Mux_h I__3411 (
            .O(N__14790),
            .I(N__14737));
    LocalMux I__3410 (
            .O(N__14785),
            .I(N__14734));
    Span4Mux_h I__3409 (
            .O(N__14782),
            .I(N__14729));
    LocalMux I__3408 (
            .O(N__14777),
            .I(N__14729));
    Span4Mux_h I__3407 (
            .O(N__14770),
            .I(N__14724));
    LocalMux I__3406 (
            .O(N__14767),
            .I(N__14724));
    LocalMux I__3405 (
            .O(N__14764),
            .I(N__14717));
    LocalMux I__3404 (
            .O(N__14761),
            .I(N__14717));
    Span4Mux_v I__3403 (
            .O(N__14758),
            .I(N__14717));
    Span4Mux_h I__3402 (
            .O(N__14755),
            .I(N__14714));
    InMux I__3401 (
            .O(N__14754),
            .I(N__14711));
    InMux I__3400 (
            .O(N__14753),
            .I(N__14706));
    InMux I__3399 (
            .O(N__14752),
            .I(N__14706));
    Span4Mux_h I__3398 (
            .O(N__14747),
            .I(N__14701));
    Span4Mux_h I__3397 (
            .O(N__14742),
            .I(N__14701));
    InMux I__3396 (
            .O(N__14741),
            .I(N__14696));
    InMux I__3395 (
            .O(N__14740),
            .I(N__14696));
    Span4Mux_h I__3394 (
            .O(N__14737),
            .I(N__14689));
    Span4Mux_h I__3393 (
            .O(N__14734),
            .I(N__14689));
    Span4Mux_h I__3392 (
            .O(N__14729),
            .I(N__14689));
    Span4Mux_v I__3391 (
            .O(N__14724),
            .I(N__14684));
    Span4Mux_h I__3390 (
            .O(N__14717),
            .I(N__14684));
    Odrv4 I__3389 (
            .O(N__14714),
            .I(aZ0Z_0));
    LocalMux I__3388 (
            .O(N__14711),
            .I(aZ0Z_0));
    LocalMux I__3387 (
            .O(N__14706),
            .I(aZ0Z_0));
    Odrv4 I__3386 (
            .O(N__14701),
            .I(aZ0Z_0));
    LocalMux I__3385 (
            .O(N__14696),
            .I(aZ0Z_0));
    Odrv4 I__3384 (
            .O(N__14689),
            .I(aZ0Z_0));
    Odrv4 I__3383 (
            .O(N__14684),
            .I(aZ0Z_0));
    InMux I__3382 (
            .O(N__14669),
            .I(N__14666));
    LocalMux I__3381 (
            .O(N__14666),
            .I(N__14663));
    Odrv12 I__3380 (
            .O(N__14663),
            .I(\ALU.regsA_result_cry_13_ma ));
    InMux I__3379 (
            .O(N__14660),
            .I(N__14652));
    InMux I__3378 (
            .O(N__14659),
            .I(N__14649));
    CascadeMux I__3377 (
            .O(N__14658),
            .I(N__14645));
    InMux I__3376 (
            .O(N__14657),
            .I(N__14641));
    InMux I__3375 (
            .O(N__14656),
            .I(N__14636));
    InMux I__3374 (
            .O(N__14655),
            .I(N__14636));
    LocalMux I__3373 (
            .O(N__14652),
            .I(N__14631));
    LocalMux I__3372 (
            .O(N__14649),
            .I(N__14631));
    InMux I__3371 (
            .O(N__14648),
            .I(N__14628));
    InMux I__3370 (
            .O(N__14645),
            .I(N__14623));
    InMux I__3369 (
            .O(N__14644),
            .I(N__14623));
    LocalMux I__3368 (
            .O(N__14641),
            .I(N__14617));
    LocalMux I__3367 (
            .O(N__14636),
            .I(N__14617));
    Span4Mux_v I__3366 (
            .O(N__14631),
            .I(N__14610));
    LocalMux I__3365 (
            .O(N__14628),
            .I(N__14610));
    LocalMux I__3364 (
            .O(N__14623),
            .I(N__14610));
    InMux I__3363 (
            .O(N__14622),
            .I(N__14607));
    Span4Mux_v I__3362 (
            .O(N__14617),
            .I(N__14604));
    Span4Mux_h I__3361 (
            .O(N__14610),
            .I(N__14600));
    LocalMux I__3360 (
            .O(N__14607),
            .I(N__14597));
    Span4Mux_h I__3359 (
            .O(N__14604),
            .I(N__14594));
    InMux I__3358 (
            .O(N__14603),
            .I(N__14591));
    Span4Mux_h I__3357 (
            .O(N__14600),
            .I(N__14588));
    Odrv4 I__3356 (
            .O(N__14597),
            .I(aZ0Z_13));
    Odrv4 I__3355 (
            .O(N__14594),
            .I(aZ0Z_13));
    LocalMux I__3354 (
            .O(N__14591),
            .I(aZ0Z_13));
    Odrv4 I__3353 (
            .O(N__14588),
            .I(aZ0Z_13));
    InMux I__3352 (
            .O(N__14579),
            .I(N__14575));
    InMux I__3351 (
            .O(N__14578),
            .I(N__14572));
    LocalMux I__3350 (
            .O(N__14575),
            .I(N__14567));
    LocalMux I__3349 (
            .O(N__14572),
            .I(N__14564));
    CascadeMux I__3348 (
            .O(N__14571),
            .I(N__14561));
    InMux I__3347 (
            .O(N__14570),
            .I(N__14556));
    Span4Mux_h I__3346 (
            .O(N__14567),
            .I(N__14553));
    Span4Mux_v I__3345 (
            .O(N__14564),
            .I(N__14550));
    InMux I__3344 (
            .O(N__14561),
            .I(N__14543));
    InMux I__3343 (
            .O(N__14560),
            .I(N__14543));
    InMux I__3342 (
            .O(N__14559),
            .I(N__14543));
    LocalMux I__3341 (
            .O(N__14556),
            .I(bZ0Z_13));
    Odrv4 I__3340 (
            .O(N__14553),
            .I(bZ0Z_13));
    Odrv4 I__3339 (
            .O(N__14550),
            .I(bZ0Z_13));
    LocalMux I__3338 (
            .O(N__14543),
            .I(bZ0Z_13));
    CascadeMux I__3337 (
            .O(N__14534),
            .I(N__14531));
    InMux I__3336 (
            .O(N__14531),
            .I(N__14528));
    LocalMux I__3335 (
            .O(N__14528),
            .I(N__14525));
    Span4Mux_h I__3334 (
            .O(N__14525),
            .I(N__14522));
    Span4Mux_h I__3333 (
            .O(N__14522),
            .I(N__14519));
    Odrv4 I__3332 (
            .O(N__14519),
            .I(\ALU.addsub_axb_13_l_ofxZ0 ));
    InMux I__3331 (
            .O(N__14516),
            .I(N__14511));
    CascadeMux I__3330 (
            .O(N__14515),
            .I(N__14507));
    InMux I__3329 (
            .O(N__14514),
            .I(N__14504));
    LocalMux I__3328 (
            .O(N__14511),
            .I(N__14500));
    InMux I__3327 (
            .O(N__14510),
            .I(N__14497));
    InMux I__3326 (
            .O(N__14507),
            .I(N__14494));
    LocalMux I__3325 (
            .O(N__14504),
            .I(N__14491));
    InMux I__3324 (
            .O(N__14503),
            .I(N__14488));
    Span4Mux_h I__3323 (
            .O(N__14500),
            .I(N__14481));
    LocalMux I__3322 (
            .O(N__14497),
            .I(N__14481));
    LocalMux I__3321 (
            .O(N__14494),
            .I(N__14481));
    Span4Mux_h I__3320 (
            .O(N__14491),
            .I(N__14478));
    LocalMux I__3319 (
            .O(N__14488),
            .I(N__14475));
    Span4Mux_v I__3318 (
            .O(N__14481),
            .I(N__14472));
    Odrv4 I__3317 (
            .O(N__14478),
            .I(RXbuffer_0));
    Odrv4 I__3316 (
            .O(N__14475),
            .I(RXbuffer_0));
    Odrv4 I__3315 (
            .O(N__14472),
            .I(RXbuffer_0));
    CascadeMux I__3314 (
            .O(N__14465),
            .I(N__14460));
    InMux I__3313 (
            .O(N__14464),
            .I(N__14452));
    CascadeMux I__3312 (
            .O(N__14463),
            .I(N__14449));
    InMux I__3311 (
            .O(N__14460),
            .I(N__14440));
    InMux I__3310 (
            .O(N__14459),
            .I(N__14437));
    InMux I__3309 (
            .O(N__14458),
            .I(N__14434));
    InMux I__3308 (
            .O(N__14457),
            .I(N__14427));
    InMux I__3307 (
            .O(N__14456),
            .I(N__14427));
    InMux I__3306 (
            .O(N__14455),
            .I(N__14427));
    LocalMux I__3305 (
            .O(N__14452),
            .I(N__14423));
    InMux I__3304 (
            .O(N__14449),
            .I(N__14420));
    InMux I__3303 (
            .O(N__14448),
            .I(N__14417));
    InMux I__3302 (
            .O(N__14447),
            .I(N__14412));
    InMux I__3301 (
            .O(N__14446),
            .I(N__14412));
    InMux I__3300 (
            .O(N__14445),
            .I(N__14405));
    InMux I__3299 (
            .O(N__14444),
            .I(N__14405));
    InMux I__3298 (
            .O(N__14443),
            .I(N__14405));
    LocalMux I__3297 (
            .O(N__14440),
            .I(N__14402));
    LocalMux I__3296 (
            .O(N__14437),
            .I(N__14399));
    LocalMux I__3295 (
            .O(N__14434),
            .I(N__14396));
    LocalMux I__3294 (
            .O(N__14427),
            .I(N__14393));
    InMux I__3293 (
            .O(N__14426),
            .I(N__14390));
    Span4Mux_v I__3292 (
            .O(N__14423),
            .I(N__14379));
    LocalMux I__3291 (
            .O(N__14420),
            .I(N__14379));
    LocalMux I__3290 (
            .O(N__14417),
            .I(N__14379));
    LocalMux I__3289 (
            .O(N__14412),
            .I(N__14379));
    LocalMux I__3288 (
            .O(N__14405),
            .I(N__14379));
    Span4Mux_h I__3287 (
            .O(N__14402),
            .I(N__14376));
    Span4Mux_h I__3286 (
            .O(N__14399),
            .I(N__14373));
    Span4Mux_v I__3285 (
            .O(N__14396),
            .I(N__14363));
    Span4Mux_h I__3284 (
            .O(N__14393),
            .I(N__14363));
    LocalMux I__3283 (
            .O(N__14390),
            .I(N__14360));
    Span4Mux_h I__3282 (
            .O(N__14379),
            .I(N__14357));
    Span4Mux_h I__3281 (
            .O(N__14376),
            .I(N__14352));
    Span4Mux_h I__3280 (
            .O(N__14373),
            .I(N__14352));
    InMux I__3279 (
            .O(N__14372),
            .I(N__14349));
    InMux I__3278 (
            .O(N__14371),
            .I(N__14346));
    InMux I__3277 (
            .O(N__14370),
            .I(N__14339));
    InMux I__3276 (
            .O(N__14369),
            .I(N__14339));
    InMux I__3275 (
            .O(N__14368),
            .I(N__14339));
    Span4Mux_h I__3274 (
            .O(N__14363),
            .I(N__14334));
    Span4Mux_h I__3273 (
            .O(N__14360),
            .I(N__14334));
    Span4Mux_h I__3272 (
            .O(N__14357),
            .I(N__14331));
    Odrv4 I__3271 (
            .O(N__14352),
            .I(opZ0Z_0));
    LocalMux I__3270 (
            .O(N__14349),
            .I(opZ0Z_0));
    LocalMux I__3269 (
            .O(N__14346),
            .I(opZ0Z_0));
    LocalMux I__3268 (
            .O(N__14339),
            .I(opZ0Z_0));
    Odrv4 I__3267 (
            .O(N__14334),
            .I(opZ0Z_0));
    Odrv4 I__3266 (
            .O(N__14331),
            .I(opZ0Z_0));
    InMux I__3265 (
            .O(N__14318),
            .I(N__14314));
    InMux I__3264 (
            .O(N__14317),
            .I(N__14311));
    LocalMux I__3263 (
            .O(N__14314),
            .I(N__14308));
    LocalMux I__3262 (
            .O(N__14311),
            .I(N__14304));
    Span4Mux_v I__3261 (
            .O(N__14308),
            .I(N__14301));
    InMux I__3260 (
            .O(N__14307),
            .I(N__14298));
    Span4Mux_v I__3259 (
            .O(N__14304),
            .I(N__14293));
    Span4Mux_h I__3258 (
            .O(N__14301),
            .I(N__14288));
    LocalMux I__3257 (
            .O(N__14298),
            .I(N__14288));
    InMux I__3256 (
            .O(N__14297),
            .I(N__14285));
    InMux I__3255 (
            .O(N__14296),
            .I(N__14282));
    Span4Mux_v I__3254 (
            .O(N__14293),
            .I(N__14277));
    Span4Mux_v I__3253 (
            .O(N__14288),
            .I(N__14277));
    LocalMux I__3252 (
            .O(N__14285),
            .I(N__14274));
    LocalMux I__3251 (
            .O(N__14282),
            .I(RXbuffer_6));
    Odrv4 I__3250 (
            .O(N__14277),
            .I(RXbuffer_6));
    Odrv4 I__3249 (
            .O(N__14274),
            .I(RXbuffer_6));
    InMux I__3248 (
            .O(N__14267),
            .I(N__14263));
    InMux I__3247 (
            .O(N__14266),
            .I(N__14260));
    LocalMux I__3246 (
            .O(N__14263),
            .I(N__14257));
    LocalMux I__3245 (
            .O(N__14260),
            .I(N__14252));
    Span4Mux_v I__3244 (
            .O(N__14257),
            .I(N__14249));
    InMux I__3243 (
            .O(N__14256),
            .I(N__14244));
    InMux I__3242 (
            .O(N__14255),
            .I(N__14244));
    Span4Mux_h I__3241 (
            .O(N__14252),
            .I(N__14240));
    Sp12to4 I__3240 (
            .O(N__14249),
            .I(N__14235));
    LocalMux I__3239 (
            .O(N__14244),
            .I(N__14235));
    InMux I__3238 (
            .O(N__14243),
            .I(N__14232));
    Odrv4 I__3237 (
            .O(N__14240),
            .I(bZ0Z_14));
    Odrv12 I__3236 (
            .O(N__14235),
            .I(bZ0Z_14));
    LocalMux I__3235 (
            .O(N__14232),
            .I(bZ0Z_14));
    CEMux I__3234 (
            .O(N__14225),
            .I(N__14220));
    CEMux I__3233 (
            .O(N__14224),
            .I(N__14216));
    CEMux I__3232 (
            .O(N__14223),
            .I(N__14212));
    LocalMux I__3231 (
            .O(N__14220),
            .I(N__14209));
    CEMux I__3230 (
            .O(N__14219),
            .I(N__14206));
    LocalMux I__3229 (
            .O(N__14216),
            .I(N__14203));
    CEMux I__3228 (
            .O(N__14215),
            .I(N__14200));
    LocalMux I__3227 (
            .O(N__14212),
            .I(N__14196));
    Span4Mux_h I__3226 (
            .O(N__14209),
            .I(N__14193));
    LocalMux I__3225 (
            .O(N__14206),
            .I(N__14190));
    Span4Mux_h I__3224 (
            .O(N__14203),
            .I(N__14185));
    LocalMux I__3223 (
            .O(N__14200),
            .I(N__14185));
    CEMux I__3222 (
            .O(N__14199),
            .I(N__14182));
    Span4Mux_h I__3221 (
            .O(N__14196),
            .I(N__14179));
    Span4Mux_h I__3220 (
            .O(N__14193),
            .I(N__14172));
    Span4Mux_v I__3219 (
            .O(N__14190),
            .I(N__14172));
    Span4Mux_v I__3218 (
            .O(N__14185),
            .I(N__14172));
    LocalMux I__3217 (
            .O(N__14182),
            .I(N__14169));
    Odrv4 I__3216 (
            .O(N__14179),
            .I(RXready_RNIICV7));
    Odrv4 I__3215 (
            .O(N__14172),
            .I(RXready_RNIICV7));
    Odrv4 I__3214 (
            .O(N__14169),
            .I(RXready_RNIICV7));
    CascadeMux I__3213 (
            .O(N__14162),
            .I(N__14158));
    InMux I__3212 (
            .O(N__14161),
            .I(N__14154));
    InMux I__3211 (
            .O(N__14158),
            .I(N__14150));
    CascadeMux I__3210 (
            .O(N__14157),
            .I(N__14145));
    LocalMux I__3209 (
            .O(N__14154),
            .I(N__14142));
    CascadeMux I__3208 (
            .O(N__14153),
            .I(N__14139));
    LocalMux I__3207 (
            .O(N__14150),
            .I(N__14136));
    InMux I__3206 (
            .O(N__14149),
            .I(N__14131));
    InMux I__3205 (
            .O(N__14148),
            .I(N__14131));
    InMux I__3204 (
            .O(N__14145),
            .I(N__14124));
    Span4Mux_v I__3203 (
            .O(N__14142),
            .I(N__14121));
    InMux I__3202 (
            .O(N__14139),
            .I(N__14118));
    Span4Mux_h I__3201 (
            .O(N__14136),
            .I(N__14113));
    LocalMux I__3200 (
            .O(N__14131),
            .I(N__14113));
    InMux I__3199 (
            .O(N__14130),
            .I(N__14109));
    InMux I__3198 (
            .O(N__14129),
            .I(N__14102));
    InMux I__3197 (
            .O(N__14128),
            .I(N__14102));
    InMux I__3196 (
            .O(N__14127),
            .I(N__14102));
    LocalMux I__3195 (
            .O(N__14124),
            .I(N__14099));
    Span4Mux_h I__3194 (
            .O(N__14121),
            .I(N__14092));
    LocalMux I__3193 (
            .O(N__14118),
            .I(N__14092));
    Span4Mux_v I__3192 (
            .O(N__14113),
            .I(N__14092));
    InMux I__3191 (
            .O(N__14112),
            .I(N__14089));
    LocalMux I__3190 (
            .O(N__14109),
            .I(bZ0Z_10));
    LocalMux I__3189 (
            .O(N__14102),
            .I(bZ0Z_10));
    Odrv4 I__3188 (
            .O(N__14099),
            .I(bZ0Z_10));
    Odrv4 I__3187 (
            .O(N__14092),
            .I(bZ0Z_10));
    LocalMux I__3186 (
            .O(N__14089),
            .I(bZ0Z_10));
    InMux I__3185 (
            .O(N__14078),
            .I(N__14075));
    LocalMux I__3184 (
            .O(N__14075),
            .I(N__14072));
    Span4Mux_h I__3183 (
            .O(N__14072),
            .I(N__14069));
    Span4Mux_h I__3182 (
            .O(N__14069),
            .I(N__14066));
    Odrv4 I__3181 (
            .O(N__14066),
            .I(\ALU.regsA_result_cry_9_ma ));
    InMux I__3180 (
            .O(N__14063),
            .I(N__14060));
    LocalMux I__3179 (
            .O(N__14060),
            .I(N__14057));
    Span4Mux_h I__3178 (
            .O(N__14057),
            .I(N__14053));
    IoInMux I__3177 (
            .O(N__14056),
            .I(N__14050));
    Span4Mux_h I__3176 (
            .O(N__14053),
            .I(N__14047));
    LocalMux I__3175 (
            .O(N__14050),
            .I(N__14044));
    Sp12to4 I__3174 (
            .O(N__14047),
            .I(N__14041));
    IoSpan4Mux I__3173 (
            .O(N__14044),
            .I(N__14038));
    Span12Mux_v I__3172 (
            .O(N__14041),
            .I(N__14035));
    Span4Mux_s2_v I__3171 (
            .O(N__14038),
            .I(N__14032));
    Odrv12 I__3170 (
            .O(N__14035),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3169 (
            .O(N__14032),
            .I(CONSTANT_ONE_NET));
    InMux I__3168 (
            .O(N__14027),
            .I(N__14024));
    LocalMux I__3167 (
            .O(N__14024),
            .I(N__14021));
    Span12Mux_v I__3166 (
            .O(N__14021),
            .I(N__14014));
    InMux I__3165 (
            .O(N__14020),
            .I(N__14011));
    InMux I__3164 (
            .O(N__14019),
            .I(N__14008));
    InMux I__3163 (
            .O(N__14018),
            .I(N__14003));
    InMux I__3162 (
            .O(N__14017),
            .I(N__14003));
    Odrv12 I__3161 (
            .O(N__14014),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__3160 (
            .O(N__14011),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__3159 (
            .O(N__14008),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__3158 (
            .O(N__14003),
            .I(\FTDI.un3_TX_0 ));
    InMux I__3157 (
            .O(N__13994),
            .I(N__13985));
    InMux I__3156 (
            .O(N__13993),
            .I(N__13985));
    InMux I__3155 (
            .O(N__13992),
            .I(N__13985));
    LocalMux I__3154 (
            .O(N__13985),
            .I(\FTDI.gap8 ));
    InMux I__3153 (
            .O(N__13982),
            .I(N__13976));
    InMux I__3152 (
            .O(N__13981),
            .I(N__13976));
    LocalMux I__3151 (
            .O(N__13976),
            .I(\FTDI.gapZ0Z_1 ));
    CascadeMux I__3150 (
            .O(N__13973),
            .I(N__13970));
    InMux I__3149 (
            .O(N__13970),
            .I(N__13961));
    InMux I__3148 (
            .O(N__13969),
            .I(N__13961));
    InMux I__3147 (
            .O(N__13968),
            .I(N__13961));
    LocalMux I__3146 (
            .O(N__13961),
            .I(\FTDI.gapZ0Z_0 ));
    CascadeMux I__3145 (
            .O(N__13958),
            .I(N__13953));
    CascadeMux I__3144 (
            .O(N__13957),
            .I(N__13947));
    InMux I__3143 (
            .O(N__13956),
            .I(N__13938));
    InMux I__3142 (
            .O(N__13953),
            .I(N__13938));
    InMux I__3141 (
            .O(N__13952),
            .I(N__13938));
    InMux I__3140 (
            .O(N__13951),
            .I(N__13938));
    InMux I__3139 (
            .O(N__13950),
            .I(N__13933));
    InMux I__3138 (
            .O(N__13947),
            .I(N__13933));
    LocalMux I__3137 (
            .O(N__13938),
            .I(\FTDI.gapZ0Z_2 ));
    LocalMux I__3136 (
            .O(N__13933),
            .I(\FTDI.gapZ0Z_2 ));
    CascadeMux I__3135 (
            .O(N__13928),
            .I(N__13925));
    InMux I__3134 (
            .O(N__13925),
            .I(N__13922));
    LocalMux I__3133 (
            .O(N__13922),
            .I(N__13919));
    Span4Mux_h I__3132 (
            .O(N__13919),
            .I(N__13916));
    Odrv4 I__3131 (
            .O(N__13916),
            .I(\ALU.addsub_axb_6_l_ofxZ0 ));
    InMux I__3130 (
            .O(N__13913),
            .I(N__13910));
    LocalMux I__3129 (
            .O(N__13910),
            .I(N__13907));
    Span4Mux_v I__3128 (
            .O(N__13907),
            .I(N__13902));
    InMux I__3127 (
            .O(N__13906),
            .I(N__13899));
    CascadeMux I__3126 (
            .O(N__13905),
            .I(N__13896));
    Span4Mux_v I__3125 (
            .O(N__13902),
            .I(N__13893));
    LocalMux I__3124 (
            .O(N__13899),
            .I(N__13890));
    InMux I__3123 (
            .O(N__13896),
            .I(N__13887));
    Odrv4 I__3122 (
            .O(N__13893),
            .I(\ALU.mult_AdderTree2_bigtree_600 ));
    Odrv4 I__3121 (
            .O(N__13890),
            .I(\ALU.mult_AdderTree2_bigtree_600 ));
    LocalMux I__3120 (
            .O(N__13887),
            .I(\ALU.mult_AdderTree2_bigtree_600 ));
    CascadeMux I__3119 (
            .O(N__13880),
            .I(N__13875));
    InMux I__3118 (
            .O(N__13879),
            .I(N__13870));
    CascadeMux I__3117 (
            .O(N__13878),
            .I(N__13860));
    InMux I__3116 (
            .O(N__13875),
            .I(N__13855));
    InMux I__3115 (
            .O(N__13874),
            .I(N__13855));
    CascadeMux I__3114 (
            .O(N__13873),
            .I(N__13852));
    LocalMux I__3113 (
            .O(N__13870),
            .I(N__13849));
    InMux I__3112 (
            .O(N__13869),
            .I(N__13846));
    InMux I__3111 (
            .O(N__13868),
            .I(N__13843));
    InMux I__3110 (
            .O(N__13867),
            .I(N__13840));
    CascadeMux I__3109 (
            .O(N__13866),
            .I(N__13837));
    CascadeMux I__3108 (
            .O(N__13865),
            .I(N__13833));
    CascadeMux I__3107 (
            .O(N__13864),
            .I(N__13829));
    InMux I__3106 (
            .O(N__13863),
            .I(N__13823));
    InMux I__3105 (
            .O(N__13860),
            .I(N__13823));
    LocalMux I__3104 (
            .O(N__13855),
            .I(N__13820));
    InMux I__3103 (
            .O(N__13852),
            .I(N__13817));
    Span4Mux_h I__3102 (
            .O(N__13849),
            .I(N__13808));
    LocalMux I__3101 (
            .O(N__13846),
            .I(N__13808));
    LocalMux I__3100 (
            .O(N__13843),
            .I(N__13808));
    LocalMux I__3099 (
            .O(N__13840),
            .I(N__13808));
    InMux I__3098 (
            .O(N__13837),
            .I(N__13795));
    InMux I__3097 (
            .O(N__13836),
            .I(N__13795));
    InMux I__3096 (
            .O(N__13833),
            .I(N__13795));
    InMux I__3095 (
            .O(N__13832),
            .I(N__13795));
    InMux I__3094 (
            .O(N__13829),
            .I(N__13795));
    InMux I__3093 (
            .O(N__13828),
            .I(N__13795));
    LocalMux I__3092 (
            .O(N__13823),
            .I(aZ0Z_6));
    Odrv4 I__3091 (
            .O(N__13820),
            .I(aZ0Z_6));
    LocalMux I__3090 (
            .O(N__13817),
            .I(aZ0Z_6));
    Odrv4 I__3089 (
            .O(N__13808),
            .I(aZ0Z_6));
    LocalMux I__3088 (
            .O(N__13795),
            .I(aZ0Z_6));
    InMux I__3087 (
            .O(N__13784),
            .I(N__13777));
    CascadeMux I__3086 (
            .O(N__13783),
            .I(N__13773));
    InMux I__3085 (
            .O(N__13782),
            .I(N__13762));
    InMux I__3084 (
            .O(N__13781),
            .I(N__13759));
    InMux I__3083 (
            .O(N__13780),
            .I(N__13756));
    LocalMux I__3082 (
            .O(N__13777),
            .I(N__13752));
    InMux I__3081 (
            .O(N__13776),
            .I(N__13749));
    InMux I__3080 (
            .O(N__13773),
            .I(N__13745));
    InMux I__3079 (
            .O(N__13772),
            .I(N__13741));
    InMux I__3078 (
            .O(N__13771),
            .I(N__13736));
    InMux I__3077 (
            .O(N__13770),
            .I(N__13736));
    InMux I__3076 (
            .O(N__13769),
            .I(N__13729));
    InMux I__3075 (
            .O(N__13768),
            .I(N__13729));
    InMux I__3074 (
            .O(N__13767),
            .I(N__13729));
    CascadeMux I__3073 (
            .O(N__13766),
            .I(N__13718));
    InMux I__3072 (
            .O(N__13765),
            .I(N__13713));
    LocalMux I__3071 (
            .O(N__13762),
            .I(N__13710));
    LocalMux I__3070 (
            .O(N__13759),
            .I(N__13705));
    LocalMux I__3069 (
            .O(N__13756),
            .I(N__13705));
    InMux I__3068 (
            .O(N__13755),
            .I(N__13702));
    Span4Mux_v I__3067 (
            .O(N__13752),
            .I(N__13697));
    LocalMux I__3066 (
            .O(N__13749),
            .I(N__13697));
    InMux I__3065 (
            .O(N__13748),
            .I(N__13694));
    LocalMux I__3064 (
            .O(N__13745),
            .I(N__13691));
    InMux I__3063 (
            .O(N__13744),
            .I(N__13688));
    LocalMux I__3062 (
            .O(N__13741),
            .I(N__13683));
    LocalMux I__3061 (
            .O(N__13736),
            .I(N__13683));
    LocalMux I__3060 (
            .O(N__13729),
            .I(N__13680));
    InMux I__3059 (
            .O(N__13728),
            .I(N__13677));
    InMux I__3058 (
            .O(N__13727),
            .I(N__13664));
    InMux I__3057 (
            .O(N__13726),
            .I(N__13664));
    InMux I__3056 (
            .O(N__13725),
            .I(N__13657));
    InMux I__3055 (
            .O(N__13724),
            .I(N__13657));
    InMux I__3054 (
            .O(N__13723),
            .I(N__13657));
    InMux I__3053 (
            .O(N__13722),
            .I(N__13652));
    InMux I__3052 (
            .O(N__13721),
            .I(N__13652));
    InMux I__3051 (
            .O(N__13718),
            .I(N__13645));
    InMux I__3050 (
            .O(N__13717),
            .I(N__13645));
    InMux I__3049 (
            .O(N__13716),
            .I(N__13645));
    LocalMux I__3048 (
            .O(N__13713),
            .I(N__13639));
    Span4Mux_h I__3047 (
            .O(N__13710),
            .I(N__13632));
    Span4Mux_v I__3046 (
            .O(N__13705),
            .I(N__13632));
    LocalMux I__3045 (
            .O(N__13702),
            .I(N__13632));
    Span4Mux_h I__3044 (
            .O(N__13697),
            .I(N__13627));
    LocalMux I__3043 (
            .O(N__13694),
            .I(N__13627));
    Span4Mux_h I__3042 (
            .O(N__13691),
            .I(N__13616));
    LocalMux I__3041 (
            .O(N__13688),
            .I(N__13616));
    Span4Mux_v I__3040 (
            .O(N__13683),
            .I(N__13616));
    Span4Mux_v I__3039 (
            .O(N__13680),
            .I(N__13616));
    LocalMux I__3038 (
            .O(N__13677),
            .I(N__13616));
    InMux I__3037 (
            .O(N__13676),
            .I(N__13611));
    InMux I__3036 (
            .O(N__13675),
            .I(N__13611));
    InMux I__3035 (
            .O(N__13674),
            .I(N__13602));
    InMux I__3034 (
            .O(N__13673),
            .I(N__13602));
    InMux I__3033 (
            .O(N__13672),
            .I(N__13602));
    InMux I__3032 (
            .O(N__13671),
            .I(N__13602));
    InMux I__3031 (
            .O(N__13670),
            .I(N__13597));
    InMux I__3030 (
            .O(N__13669),
            .I(N__13597));
    LocalMux I__3029 (
            .O(N__13664),
            .I(N__13594));
    LocalMux I__3028 (
            .O(N__13657),
            .I(N__13587));
    LocalMux I__3027 (
            .O(N__13652),
            .I(N__13587));
    LocalMux I__3026 (
            .O(N__13645),
            .I(N__13587));
    InMux I__3025 (
            .O(N__13644),
            .I(N__13582));
    InMux I__3024 (
            .O(N__13643),
            .I(N__13582));
    InMux I__3023 (
            .O(N__13642),
            .I(N__13579));
    Span4Mux_h I__3022 (
            .O(N__13639),
            .I(N__13574));
    Span4Mux_h I__3021 (
            .O(N__13632),
            .I(N__13574));
    Span4Mux_h I__3020 (
            .O(N__13627),
            .I(N__13567));
    Span4Mux_h I__3019 (
            .O(N__13616),
            .I(N__13567));
    LocalMux I__3018 (
            .O(N__13611),
            .I(N__13567));
    LocalMux I__3017 (
            .O(N__13602),
            .I(bZ0Z_0));
    LocalMux I__3016 (
            .O(N__13597),
            .I(bZ0Z_0));
    Odrv12 I__3015 (
            .O(N__13594),
            .I(bZ0Z_0));
    Odrv12 I__3014 (
            .O(N__13587),
            .I(bZ0Z_0));
    LocalMux I__3013 (
            .O(N__13582),
            .I(bZ0Z_0));
    LocalMux I__3012 (
            .O(N__13579),
            .I(bZ0Z_0));
    Odrv4 I__3011 (
            .O(N__13574),
            .I(bZ0Z_0));
    Odrv4 I__3010 (
            .O(N__13567),
            .I(bZ0Z_0));
    InMux I__3009 (
            .O(N__13550),
            .I(N__13547));
    LocalMux I__3008 (
            .O(N__13547),
            .I(N__13544));
    Span4Mux_h I__3007 (
            .O(N__13544),
            .I(N__13541));
    Odrv4 I__3006 (
            .O(N__13541),
            .I(\ALU.regsA_result_cry_2_c_RNO_1 ));
    CascadeMux I__3005 (
            .O(N__13538),
            .I(N__13530));
    CascadeMux I__3004 (
            .O(N__13537),
            .I(N__13527));
    CascadeMux I__3003 (
            .O(N__13536),
            .I(N__13524));
    CascadeMux I__3002 (
            .O(N__13535),
            .I(N__13516));
    InMux I__3001 (
            .O(N__13534),
            .I(N__13509));
    InMux I__3000 (
            .O(N__13533),
            .I(N__13506));
    InMux I__2999 (
            .O(N__13530),
            .I(N__13499));
    InMux I__2998 (
            .O(N__13527),
            .I(N__13499));
    InMux I__2997 (
            .O(N__13524),
            .I(N__13499));
    InMux I__2996 (
            .O(N__13523),
            .I(N__13496));
    CascadeMux I__2995 (
            .O(N__13522),
            .I(N__13492));
    CascadeMux I__2994 (
            .O(N__13521),
            .I(N__13489));
    InMux I__2993 (
            .O(N__13520),
            .I(N__13485));
    InMux I__2992 (
            .O(N__13519),
            .I(N__13482));
    InMux I__2991 (
            .O(N__13516),
            .I(N__13475));
    InMux I__2990 (
            .O(N__13515),
            .I(N__13475));
    InMux I__2989 (
            .O(N__13514),
            .I(N__13475));
    InMux I__2988 (
            .O(N__13513),
            .I(N__13472));
    InMux I__2987 (
            .O(N__13512),
            .I(N__13469));
    LocalMux I__2986 (
            .O(N__13509),
            .I(N__13460));
    LocalMux I__2985 (
            .O(N__13506),
            .I(N__13457));
    LocalMux I__2984 (
            .O(N__13499),
            .I(N__13454));
    LocalMux I__2983 (
            .O(N__13496),
            .I(N__13451));
    InMux I__2982 (
            .O(N__13495),
            .I(N__13448));
    InMux I__2981 (
            .O(N__13492),
            .I(N__13441));
    InMux I__2980 (
            .O(N__13489),
            .I(N__13441));
    InMux I__2979 (
            .O(N__13488),
            .I(N__13441));
    LocalMux I__2978 (
            .O(N__13485),
            .I(N__13431));
    LocalMux I__2977 (
            .O(N__13482),
            .I(N__13428));
    LocalMux I__2976 (
            .O(N__13475),
            .I(N__13425));
    LocalMux I__2975 (
            .O(N__13472),
            .I(N__13422));
    LocalMux I__2974 (
            .O(N__13469),
            .I(N__13419));
    InMux I__2973 (
            .O(N__13468),
            .I(N__13416));
    InMux I__2972 (
            .O(N__13467),
            .I(N__13411));
    InMux I__2971 (
            .O(N__13466),
            .I(N__13411));
    InMux I__2970 (
            .O(N__13465),
            .I(N__13404));
    InMux I__2969 (
            .O(N__13464),
            .I(N__13404));
    InMux I__2968 (
            .O(N__13463),
            .I(N__13404));
    Span4Mux_v I__2967 (
            .O(N__13460),
            .I(N__13401));
    Span4Mux_v I__2966 (
            .O(N__13457),
            .I(N__13390));
    Span4Mux_h I__2965 (
            .O(N__13454),
            .I(N__13390));
    Span4Mux_h I__2964 (
            .O(N__13451),
            .I(N__13390));
    LocalMux I__2963 (
            .O(N__13448),
            .I(N__13390));
    LocalMux I__2962 (
            .O(N__13441),
            .I(N__13390));
    InMux I__2961 (
            .O(N__13440),
            .I(N__13377));
    InMux I__2960 (
            .O(N__13439),
            .I(N__13377));
    InMux I__2959 (
            .O(N__13438),
            .I(N__13377));
    InMux I__2958 (
            .O(N__13437),
            .I(N__13377));
    InMux I__2957 (
            .O(N__13436),
            .I(N__13377));
    InMux I__2956 (
            .O(N__13435),
            .I(N__13377));
    InMux I__2955 (
            .O(N__13434),
            .I(N__13374));
    Span4Mux_v I__2954 (
            .O(N__13431),
            .I(N__13365));
    Span4Mux_v I__2953 (
            .O(N__13428),
            .I(N__13365));
    Span4Mux_v I__2952 (
            .O(N__13425),
            .I(N__13365));
    Span4Mux_v I__2951 (
            .O(N__13422),
            .I(N__13365));
    Odrv12 I__2950 (
            .O(N__13419),
            .I(aZ0Z_3));
    LocalMux I__2949 (
            .O(N__13416),
            .I(aZ0Z_3));
    LocalMux I__2948 (
            .O(N__13411),
            .I(aZ0Z_3));
    LocalMux I__2947 (
            .O(N__13404),
            .I(aZ0Z_3));
    Odrv4 I__2946 (
            .O(N__13401),
            .I(aZ0Z_3));
    Odrv4 I__2945 (
            .O(N__13390),
            .I(aZ0Z_3));
    LocalMux I__2944 (
            .O(N__13377),
            .I(aZ0Z_3));
    LocalMux I__2943 (
            .O(N__13374),
            .I(aZ0Z_3));
    Odrv4 I__2942 (
            .O(N__13365),
            .I(aZ0Z_3));
    InMux I__2941 (
            .O(N__13346),
            .I(N__13339));
    InMux I__2940 (
            .O(N__13345),
            .I(N__13335));
    InMux I__2939 (
            .O(N__13344),
            .I(N__13331));
    InMux I__2938 (
            .O(N__13343),
            .I(N__13326));
    InMux I__2937 (
            .O(N__13342),
            .I(N__13326));
    LocalMux I__2936 (
            .O(N__13339),
            .I(N__13322));
    InMux I__2935 (
            .O(N__13338),
            .I(N__13319));
    LocalMux I__2934 (
            .O(N__13335),
            .I(N__13312));
    InMux I__2933 (
            .O(N__13334),
            .I(N__13309));
    LocalMux I__2932 (
            .O(N__13331),
            .I(N__13306));
    LocalMux I__2931 (
            .O(N__13326),
            .I(N__13303));
    InMux I__2930 (
            .O(N__13325),
            .I(N__13300));
    Span4Mux_v I__2929 (
            .O(N__13322),
            .I(N__13291));
    LocalMux I__2928 (
            .O(N__13319),
            .I(N__13291));
    InMux I__2927 (
            .O(N__13318),
            .I(N__13288));
    InMux I__2926 (
            .O(N__13317),
            .I(N__13282));
    InMux I__2925 (
            .O(N__13316),
            .I(N__13277));
    InMux I__2924 (
            .O(N__13315),
            .I(N__13277));
    Span4Mux_v I__2923 (
            .O(N__13312),
            .I(N__13270));
    LocalMux I__2922 (
            .O(N__13309),
            .I(N__13270));
    Span4Mux_h I__2921 (
            .O(N__13306),
            .I(N__13270));
    Span4Mux_h I__2920 (
            .O(N__13303),
            .I(N__13265));
    LocalMux I__2919 (
            .O(N__13300),
            .I(N__13265));
    InMux I__2918 (
            .O(N__13299),
            .I(N__13261));
    InMux I__2917 (
            .O(N__13298),
            .I(N__13256));
    InMux I__2916 (
            .O(N__13297),
            .I(N__13256));
    InMux I__2915 (
            .O(N__13296),
            .I(N__13253));
    Span4Mux_v I__2914 (
            .O(N__13291),
            .I(N__13247));
    LocalMux I__2913 (
            .O(N__13288),
            .I(N__13247));
    InMux I__2912 (
            .O(N__13287),
            .I(N__13244));
    InMux I__2911 (
            .O(N__13286),
            .I(N__13239));
    InMux I__2910 (
            .O(N__13285),
            .I(N__13239));
    LocalMux I__2909 (
            .O(N__13282),
            .I(N__13234));
    LocalMux I__2908 (
            .O(N__13277),
            .I(N__13234));
    Span4Mux_h I__2907 (
            .O(N__13270),
            .I(N__13229));
    Span4Mux_h I__2906 (
            .O(N__13265),
            .I(N__13229));
    InMux I__2905 (
            .O(N__13264),
            .I(N__13226));
    LocalMux I__2904 (
            .O(N__13261),
            .I(N__13223));
    LocalMux I__2903 (
            .O(N__13256),
            .I(N__13218));
    LocalMux I__2902 (
            .O(N__13253),
            .I(N__13218));
    InMux I__2901 (
            .O(N__13252),
            .I(N__13215));
    Odrv4 I__2900 (
            .O(N__13247),
            .I(bZ0Z_3));
    LocalMux I__2899 (
            .O(N__13244),
            .I(bZ0Z_3));
    LocalMux I__2898 (
            .O(N__13239),
            .I(bZ0Z_3));
    Odrv12 I__2897 (
            .O(N__13234),
            .I(bZ0Z_3));
    Odrv4 I__2896 (
            .O(N__13229),
            .I(bZ0Z_3));
    LocalMux I__2895 (
            .O(N__13226),
            .I(bZ0Z_3));
    Odrv4 I__2894 (
            .O(N__13223),
            .I(bZ0Z_3));
    Odrv12 I__2893 (
            .O(N__13218),
            .I(bZ0Z_3));
    LocalMux I__2892 (
            .O(N__13215),
            .I(bZ0Z_3));
    CascadeMux I__2891 (
            .O(N__13196),
            .I(N__13193));
    InMux I__2890 (
            .O(N__13193),
            .I(N__13190));
    LocalMux I__2889 (
            .O(N__13190),
            .I(N__13187));
    Odrv12 I__2888 (
            .O(N__13187),
            .I(\ALU.addsub_axb_3_l_ofxZ0 ));
    CascadeMux I__2887 (
            .O(N__13184),
            .I(N__13179));
    InMux I__2886 (
            .O(N__13183),
            .I(N__13175));
    InMux I__2885 (
            .O(N__13182),
            .I(N__13172));
    InMux I__2884 (
            .O(N__13179),
            .I(N__13168));
    InMux I__2883 (
            .O(N__13178),
            .I(N__13165));
    LocalMux I__2882 (
            .O(N__13175),
            .I(N__13160));
    LocalMux I__2881 (
            .O(N__13172),
            .I(N__13160));
    InMux I__2880 (
            .O(N__13171),
            .I(N__13157));
    LocalMux I__2879 (
            .O(N__13168),
            .I(N__13145));
    LocalMux I__2878 (
            .O(N__13165),
            .I(N__13142));
    Span4Mux_v I__2877 (
            .O(N__13160),
            .I(N__13137));
    LocalMux I__2876 (
            .O(N__13157),
            .I(N__13137));
    InMux I__2875 (
            .O(N__13156),
            .I(N__13132));
    InMux I__2874 (
            .O(N__13155),
            .I(N__13132));
    InMux I__2873 (
            .O(N__13154),
            .I(N__13129));
    InMux I__2872 (
            .O(N__13153),
            .I(N__13126));
    InMux I__2871 (
            .O(N__13152),
            .I(N__13115));
    InMux I__2870 (
            .O(N__13151),
            .I(N__13115));
    InMux I__2869 (
            .O(N__13150),
            .I(N__13115));
    InMux I__2868 (
            .O(N__13149),
            .I(N__13115));
    InMux I__2867 (
            .O(N__13148),
            .I(N__13115));
    Span4Mux_v I__2866 (
            .O(N__13145),
            .I(N__13108));
    Span4Mux_h I__2865 (
            .O(N__13142),
            .I(N__13108));
    Span4Mux_h I__2864 (
            .O(N__13137),
            .I(N__13108));
    LocalMux I__2863 (
            .O(N__13132),
            .I(bZ0Z_8));
    LocalMux I__2862 (
            .O(N__13129),
            .I(bZ0Z_8));
    LocalMux I__2861 (
            .O(N__13126),
            .I(bZ0Z_8));
    LocalMux I__2860 (
            .O(N__13115),
            .I(bZ0Z_8));
    Odrv4 I__2859 (
            .O(N__13108),
            .I(bZ0Z_8));
    InMux I__2858 (
            .O(N__13097),
            .I(N__13094));
    LocalMux I__2857 (
            .O(N__13094),
            .I(\ALU.regsA_result_cry_9_ma_2 ));
    CascadeMux I__2856 (
            .O(N__13091),
            .I(N__13086));
    CascadeMux I__2855 (
            .O(N__13090),
            .I(N__13082));
    InMux I__2854 (
            .O(N__13089),
            .I(N__13076));
    InMux I__2853 (
            .O(N__13086),
            .I(N__13073));
    InMux I__2852 (
            .O(N__13085),
            .I(N__13070));
    InMux I__2851 (
            .O(N__13082),
            .I(N__13064));
    InMux I__2850 (
            .O(N__13081),
            .I(N__13061));
    InMux I__2849 (
            .O(N__13080),
            .I(N__13056));
    InMux I__2848 (
            .O(N__13079),
            .I(N__13056));
    LocalMux I__2847 (
            .O(N__13076),
            .I(N__13049));
    LocalMux I__2846 (
            .O(N__13073),
            .I(N__13049));
    LocalMux I__2845 (
            .O(N__13070),
            .I(N__13046));
    CascadeMux I__2844 (
            .O(N__13069),
            .I(N__13040));
    CascadeMux I__2843 (
            .O(N__13068),
            .I(N__13036));
    CascadeMux I__2842 (
            .O(N__13067),
            .I(N__13033));
    LocalMux I__2841 (
            .O(N__13064),
            .I(N__13027));
    LocalMux I__2840 (
            .O(N__13061),
            .I(N__13027));
    LocalMux I__2839 (
            .O(N__13056),
            .I(N__13024));
    InMux I__2838 (
            .O(N__13055),
            .I(N__13019));
    InMux I__2837 (
            .O(N__13054),
            .I(N__13019));
    Span4Mux_v I__2836 (
            .O(N__13049),
            .I(N__13016));
    Span4Mux_h I__2835 (
            .O(N__13046),
            .I(N__13013));
    InMux I__2834 (
            .O(N__13045),
            .I(N__13010));
    InMux I__2833 (
            .O(N__13044),
            .I(N__13007));
    InMux I__2832 (
            .O(N__13043),
            .I(N__12994));
    InMux I__2831 (
            .O(N__13040),
            .I(N__12994));
    InMux I__2830 (
            .O(N__13039),
            .I(N__12994));
    InMux I__2829 (
            .O(N__13036),
            .I(N__12994));
    InMux I__2828 (
            .O(N__13033),
            .I(N__12994));
    InMux I__2827 (
            .O(N__13032),
            .I(N__12994));
    Span4Mux_h I__2826 (
            .O(N__13027),
            .I(N__12989));
    Span4Mux_h I__2825 (
            .O(N__13024),
            .I(N__12989));
    LocalMux I__2824 (
            .O(N__13019),
            .I(bZ0Z_6));
    Odrv4 I__2823 (
            .O(N__13016),
            .I(bZ0Z_6));
    Odrv4 I__2822 (
            .O(N__13013),
            .I(bZ0Z_6));
    LocalMux I__2821 (
            .O(N__13010),
            .I(bZ0Z_6));
    LocalMux I__2820 (
            .O(N__13007),
            .I(bZ0Z_6));
    LocalMux I__2819 (
            .O(N__12994),
            .I(bZ0Z_6));
    Odrv4 I__2818 (
            .O(N__12989),
            .I(bZ0Z_6));
    InMux I__2817 (
            .O(N__12974),
            .I(N__12971));
    LocalMux I__2816 (
            .O(N__12971),
            .I(\ALU.regsA_result_cry_7_ma_3 ));
    CascadeMux I__2815 (
            .O(N__12968),
            .I(N__12963));
    InMux I__2814 (
            .O(N__12967),
            .I(N__12958));
    InMux I__2813 (
            .O(N__12966),
            .I(N__12955));
    InMux I__2812 (
            .O(N__12963),
            .I(N__12952));
    CascadeMux I__2811 (
            .O(N__12962),
            .I(N__12942));
    CascadeMux I__2810 (
            .O(N__12961),
            .I(N__12935));
    LocalMux I__2809 (
            .O(N__12958),
            .I(N__12931));
    LocalMux I__2808 (
            .O(N__12955),
            .I(N__12921));
    LocalMux I__2807 (
            .O(N__12952),
            .I(N__12921));
    InMux I__2806 (
            .O(N__12951),
            .I(N__12914));
    InMux I__2805 (
            .O(N__12950),
            .I(N__12914));
    InMux I__2804 (
            .O(N__12949),
            .I(N__12914));
    InMux I__2803 (
            .O(N__12948),
            .I(N__12899));
    InMux I__2802 (
            .O(N__12947),
            .I(N__12899));
    InMux I__2801 (
            .O(N__12946),
            .I(N__12899));
    InMux I__2800 (
            .O(N__12945),
            .I(N__12899));
    InMux I__2799 (
            .O(N__12942),
            .I(N__12899));
    InMux I__2798 (
            .O(N__12941),
            .I(N__12899));
    InMux I__2797 (
            .O(N__12940),
            .I(N__12899));
    InMux I__2796 (
            .O(N__12939),
            .I(N__12894));
    InMux I__2795 (
            .O(N__12938),
            .I(N__12894));
    InMux I__2794 (
            .O(N__12935),
            .I(N__12889));
    InMux I__2793 (
            .O(N__12934),
            .I(N__12889));
    Span12Mux_v I__2792 (
            .O(N__12931),
            .I(N__12886));
    InMux I__2791 (
            .O(N__12930),
            .I(N__12875));
    InMux I__2790 (
            .O(N__12929),
            .I(N__12875));
    InMux I__2789 (
            .O(N__12928),
            .I(N__12875));
    InMux I__2788 (
            .O(N__12927),
            .I(N__12875));
    InMux I__2787 (
            .O(N__12926),
            .I(N__12875));
    Span4Mux_h I__2786 (
            .O(N__12921),
            .I(N__12866));
    LocalMux I__2785 (
            .O(N__12914),
            .I(N__12866));
    LocalMux I__2784 (
            .O(N__12899),
            .I(N__12866));
    LocalMux I__2783 (
            .O(N__12894),
            .I(N__12866));
    LocalMux I__2782 (
            .O(N__12889),
            .I(aZ0Z_7));
    Odrv12 I__2781 (
            .O(N__12886),
            .I(aZ0Z_7));
    LocalMux I__2780 (
            .O(N__12875),
            .I(aZ0Z_7));
    Odrv4 I__2779 (
            .O(N__12866),
            .I(aZ0Z_7));
    CascadeMux I__2778 (
            .O(N__12857),
            .I(N__12853));
    InMux I__2777 (
            .O(N__12856),
            .I(N__12846));
    InMux I__2776 (
            .O(N__12853),
            .I(N__12846));
    InMux I__2775 (
            .O(N__12852),
            .I(N__12839));
    InMux I__2774 (
            .O(N__12851),
            .I(N__12839));
    LocalMux I__2773 (
            .O(N__12846),
            .I(N__12836));
    InMux I__2772 (
            .O(N__12845),
            .I(N__12833));
    InMux I__2771 (
            .O(N__12844),
            .I(N__12827));
    LocalMux I__2770 (
            .O(N__12839),
            .I(N__12824));
    Span4Mux_v I__2769 (
            .O(N__12836),
            .I(N__12821));
    LocalMux I__2768 (
            .O(N__12833),
            .I(N__12818));
    InMux I__2767 (
            .O(N__12832),
            .I(N__12813));
    InMux I__2766 (
            .O(N__12831),
            .I(N__12813));
    InMux I__2765 (
            .O(N__12830),
            .I(N__12810));
    LocalMux I__2764 (
            .O(N__12827),
            .I(N__12807));
    Span4Mux_h I__2763 (
            .O(N__12824),
            .I(N__12798));
    Span4Mux_v I__2762 (
            .O(N__12821),
            .I(N__12789));
    Span4Mux_h I__2761 (
            .O(N__12818),
            .I(N__12789));
    LocalMux I__2760 (
            .O(N__12813),
            .I(N__12789));
    LocalMux I__2759 (
            .O(N__12810),
            .I(N__12789));
    Span4Mux_h I__2758 (
            .O(N__12807),
            .I(N__12786));
    InMux I__2757 (
            .O(N__12806),
            .I(N__12781));
    InMux I__2756 (
            .O(N__12805),
            .I(N__12781));
    InMux I__2755 (
            .O(N__12804),
            .I(N__12772));
    InMux I__2754 (
            .O(N__12803),
            .I(N__12772));
    InMux I__2753 (
            .O(N__12802),
            .I(N__12772));
    InMux I__2752 (
            .O(N__12801),
            .I(N__12772));
    Odrv4 I__2751 (
            .O(N__12798),
            .I(bZ0Z_7));
    Odrv4 I__2750 (
            .O(N__12789),
            .I(bZ0Z_7));
    Odrv4 I__2749 (
            .O(N__12786),
            .I(bZ0Z_7));
    LocalMux I__2748 (
            .O(N__12781),
            .I(bZ0Z_7));
    LocalMux I__2747 (
            .O(N__12772),
            .I(bZ0Z_7));
    CascadeMux I__2746 (
            .O(N__12761),
            .I(N__12758));
    InMux I__2745 (
            .O(N__12758),
            .I(N__12755));
    LocalMux I__2744 (
            .O(N__12755),
            .I(\ALU.regsA_result_cry_8_ma_2 ));
    InMux I__2743 (
            .O(N__12752),
            .I(N__12749));
    LocalMux I__2742 (
            .O(N__12749),
            .I(N__12746));
    Span4Mux_h I__2741 (
            .O(N__12746),
            .I(N__12738));
    InMux I__2740 (
            .O(N__12745),
            .I(N__12733));
    InMux I__2739 (
            .O(N__12744),
            .I(N__12733));
    InMux I__2738 (
            .O(N__12743),
            .I(N__12728));
    InMux I__2737 (
            .O(N__12742),
            .I(N__12728));
    InMux I__2736 (
            .O(N__12741),
            .I(N__12725));
    Span4Mux_h I__2735 (
            .O(N__12738),
            .I(N__12722));
    LocalMux I__2734 (
            .O(N__12733),
            .I(\FTDI.baudAccZ0Z_2 ));
    LocalMux I__2733 (
            .O(N__12728),
            .I(\FTDI.baudAccZ0Z_2 ));
    LocalMux I__2732 (
            .O(N__12725),
            .I(\FTDI.baudAccZ0Z_2 ));
    Odrv4 I__2731 (
            .O(N__12722),
            .I(\FTDI.baudAccZ0Z_2 ));
    CEMux I__2730 (
            .O(N__12713),
            .I(N__12709));
    CEMux I__2729 (
            .O(N__12712),
            .I(N__12706));
    LocalMux I__2728 (
            .O(N__12709),
            .I(N__12703));
    LocalMux I__2727 (
            .O(N__12706),
            .I(N__12700));
    Span4Mux_v I__2726 (
            .O(N__12703),
            .I(N__12697));
    Span4Mux_h I__2725 (
            .O(N__12700),
            .I(N__12694));
    Odrv4 I__2724 (
            .O(N__12697),
            .I(\FTDI.un1_TXstate_0_sqmuxa_0_i ));
    Odrv4 I__2723 (
            .O(N__12694),
            .I(\FTDI.un1_TXstate_0_sqmuxa_0_i ));
    InMux I__2722 (
            .O(N__12689),
            .I(N__12686));
    LocalMux I__2721 (
            .O(N__12686),
            .I(N__12683));
    Span4Mux_h I__2720 (
            .O(N__12683),
            .I(N__12679));
    InMux I__2719 (
            .O(N__12682),
            .I(N__12676));
    Odrv4 I__2718 (
            .O(N__12679),
            .I(TXstartZ0));
    LocalMux I__2717 (
            .O(N__12676),
            .I(TXstartZ0));
    CEMux I__2716 (
            .O(N__12671),
            .I(N__12668));
    LocalMux I__2715 (
            .O(N__12668),
            .I(N__12665));
    Sp12to4 I__2714 (
            .O(N__12665),
            .I(N__12662));
    Odrv12 I__2713 (
            .O(N__12662),
            .I(un1_testState31_0_0));
    InMux I__2712 (
            .O(N__12659),
            .I(N__12656));
    LocalMux I__2711 (
            .O(N__12656),
            .I(\ALU.regsA_result_cry_6_ma_3 ));
    CascadeMux I__2710 (
            .O(N__12653),
            .I(N__12645));
    CascadeMux I__2709 (
            .O(N__12652),
            .I(N__12642));
    InMux I__2708 (
            .O(N__12651),
            .I(N__12633));
    InMux I__2707 (
            .O(N__12650),
            .I(N__12633));
    InMux I__2706 (
            .O(N__12649),
            .I(N__12630));
    InMux I__2705 (
            .O(N__12648),
            .I(N__12627));
    InMux I__2704 (
            .O(N__12645),
            .I(N__12622));
    InMux I__2703 (
            .O(N__12642),
            .I(N__12619));
    CascadeMux I__2702 (
            .O(N__12641),
            .I(N__12616));
    CascadeMux I__2701 (
            .O(N__12640),
            .I(N__12612));
    CascadeMux I__2700 (
            .O(N__12639),
            .I(N__12609));
    InMux I__2699 (
            .O(N__12638),
            .I(N__12604));
    LocalMux I__2698 (
            .O(N__12633),
            .I(N__12597));
    LocalMux I__2697 (
            .O(N__12630),
            .I(N__12594));
    LocalMux I__2696 (
            .O(N__12627),
            .I(N__12591));
    CascadeMux I__2695 (
            .O(N__12626),
            .I(N__12588));
    CascadeMux I__2694 (
            .O(N__12625),
            .I(N__12585));
    LocalMux I__2693 (
            .O(N__12622),
            .I(N__12582));
    LocalMux I__2692 (
            .O(N__12619),
            .I(N__12579));
    InMux I__2691 (
            .O(N__12616),
            .I(N__12568));
    InMux I__2690 (
            .O(N__12615),
            .I(N__12568));
    InMux I__2689 (
            .O(N__12612),
            .I(N__12568));
    InMux I__2688 (
            .O(N__12609),
            .I(N__12568));
    InMux I__2687 (
            .O(N__12608),
            .I(N__12568));
    InMux I__2686 (
            .O(N__12607),
            .I(N__12565));
    LocalMux I__2685 (
            .O(N__12604),
            .I(N__12562));
    InMux I__2684 (
            .O(N__12603),
            .I(N__12559));
    InMux I__2683 (
            .O(N__12602),
            .I(N__12552));
    InMux I__2682 (
            .O(N__12601),
            .I(N__12552));
    InMux I__2681 (
            .O(N__12600),
            .I(N__12552));
    Span4Mux_v I__2680 (
            .O(N__12597),
            .I(N__12547));
    Span4Mux_v I__2679 (
            .O(N__12594),
            .I(N__12547));
    Span4Mux_h I__2678 (
            .O(N__12591),
            .I(N__12544));
    InMux I__2677 (
            .O(N__12588),
            .I(N__12539));
    InMux I__2676 (
            .O(N__12585),
            .I(N__12539));
    Span4Mux_h I__2675 (
            .O(N__12582),
            .I(N__12530));
    Span4Mux_v I__2674 (
            .O(N__12579),
            .I(N__12530));
    LocalMux I__2673 (
            .O(N__12568),
            .I(N__12530));
    LocalMux I__2672 (
            .O(N__12565),
            .I(N__12530));
    Odrv12 I__2671 (
            .O(N__12562),
            .I(aZ0Z_1));
    LocalMux I__2670 (
            .O(N__12559),
            .I(aZ0Z_1));
    LocalMux I__2669 (
            .O(N__12552),
            .I(aZ0Z_1));
    Odrv4 I__2668 (
            .O(N__12547),
            .I(aZ0Z_1));
    Odrv4 I__2667 (
            .O(N__12544),
            .I(aZ0Z_1));
    LocalMux I__2666 (
            .O(N__12539),
            .I(aZ0Z_1));
    Odrv4 I__2665 (
            .O(N__12530),
            .I(aZ0Z_1));
    CascadeMux I__2664 (
            .O(N__12515),
            .I(N__12512));
    InMux I__2663 (
            .O(N__12512),
            .I(N__12509));
    LocalMux I__2662 (
            .O(N__12509),
            .I(N__12506));
    Odrv12 I__2661 (
            .O(N__12506),
            .I(\ALU.regsA_result_axb_8_l_ofx ));
    InMux I__2660 (
            .O(N__12503),
            .I(N__12500));
    LocalMux I__2659 (
            .O(N__12500),
            .I(N__12497));
    Span4Mux_h I__2658 (
            .O(N__12497),
            .I(N__12494));
    Odrv4 I__2657 (
            .O(N__12494),
            .I(\ALU.regsA_result_cry_7_ma ));
    CascadeMux I__2656 (
            .O(N__12491),
            .I(N__12488));
    InMux I__2655 (
            .O(N__12488),
            .I(N__12485));
    LocalMux I__2654 (
            .O(N__12485),
            .I(N__12482));
    Span4Mux_v I__2653 (
            .O(N__12482),
            .I(N__12479));
    Odrv4 I__2652 (
            .O(N__12479),
            .I(\ALU.regsA_result_axb_8_l_ofx_1 ));
    InMux I__2651 (
            .O(N__12476),
            .I(N__12473));
    LocalMux I__2650 (
            .O(N__12473),
            .I(N__12470));
    Span4Mux_h I__2649 (
            .O(N__12470),
            .I(N__12467));
    Odrv4 I__2648 (
            .O(N__12467),
            .I(\ALU.regsA_result_cry_9_ma_1 ));
    CascadeMux I__2647 (
            .O(N__12464),
            .I(N__12461));
    InMux I__2646 (
            .O(N__12461),
            .I(N__12458));
    LocalMux I__2645 (
            .O(N__12458),
            .I(N__12450));
    InMux I__2644 (
            .O(N__12457),
            .I(N__12445));
    InMux I__2643 (
            .O(N__12456),
            .I(N__12445));
    InMux I__2642 (
            .O(N__12455),
            .I(N__12437));
    InMux I__2641 (
            .O(N__12454),
            .I(N__12437));
    InMux I__2640 (
            .O(N__12453),
            .I(N__12434));
    Span4Mux_h I__2639 (
            .O(N__12450),
            .I(N__12429));
    LocalMux I__2638 (
            .O(N__12445),
            .I(N__12429));
    InMux I__2637 (
            .O(N__12444),
            .I(N__12424));
    InMux I__2636 (
            .O(N__12443),
            .I(N__12424));
    InMux I__2635 (
            .O(N__12442),
            .I(N__12421));
    LocalMux I__2634 (
            .O(N__12437),
            .I(N__12418));
    LocalMux I__2633 (
            .O(N__12434),
            .I(N__12413));
    Span4Mux_v I__2632 (
            .O(N__12429),
            .I(N__12413));
    LocalMux I__2631 (
            .O(N__12424),
            .I(aZ0Z_2));
    LocalMux I__2630 (
            .O(N__12421),
            .I(aZ0Z_2));
    Odrv12 I__2629 (
            .O(N__12418),
            .I(aZ0Z_2));
    Odrv4 I__2628 (
            .O(N__12413),
            .I(aZ0Z_2));
    CascadeMux I__2627 (
            .O(N__12404),
            .I(N__12401));
    InMux I__2626 (
            .O(N__12401),
            .I(N__12398));
    LocalMux I__2625 (
            .O(N__12398),
            .I(N__12395));
    Span4Mux_h I__2624 (
            .O(N__12395),
            .I(N__12392));
    Odrv4 I__2623 (
            .O(N__12392),
            .I(\ALU.regsA_result_axb_9_l_ofx_1 ));
    InMux I__2622 (
            .O(N__12389),
            .I(N__12386));
    LocalMux I__2621 (
            .O(N__12386),
            .I(\ALU.regsA_result_axb_8_l_ofx_2 ));
    InMux I__2620 (
            .O(N__12383),
            .I(N__12380));
    LocalMux I__2619 (
            .O(N__12380),
            .I(N__12375));
    InMux I__2618 (
            .O(N__12379),
            .I(N__12372));
    InMux I__2617 (
            .O(N__12378),
            .I(N__12365));
    Span4Mux_v I__2616 (
            .O(N__12375),
            .I(N__12362));
    LocalMux I__2615 (
            .O(N__12372),
            .I(N__12359));
    InMux I__2614 (
            .O(N__12371),
            .I(N__12356));
    InMux I__2613 (
            .O(N__12370),
            .I(N__12348));
    InMux I__2612 (
            .O(N__12369),
            .I(N__12343));
    InMux I__2611 (
            .O(N__12368),
            .I(N__12343));
    LocalMux I__2610 (
            .O(N__12365),
            .I(N__12340));
    Span4Mux_h I__2609 (
            .O(N__12362),
            .I(N__12337));
    Span4Mux_v I__2608 (
            .O(N__12359),
            .I(N__12332));
    LocalMux I__2607 (
            .O(N__12356),
            .I(N__12332));
    InMux I__2606 (
            .O(N__12355),
            .I(N__12327));
    InMux I__2605 (
            .O(N__12354),
            .I(N__12327));
    InMux I__2604 (
            .O(N__12353),
            .I(N__12324));
    InMux I__2603 (
            .O(N__12352),
            .I(N__12319));
    InMux I__2602 (
            .O(N__12351),
            .I(N__12319));
    LocalMux I__2601 (
            .O(N__12348),
            .I(N__12314));
    LocalMux I__2600 (
            .O(N__12343),
            .I(N__12314));
    Span4Mux_h I__2599 (
            .O(N__12340),
            .I(N__12311));
    Odrv4 I__2598 (
            .O(N__12337),
            .I(bZ0Z_9));
    Odrv4 I__2597 (
            .O(N__12332),
            .I(bZ0Z_9));
    LocalMux I__2596 (
            .O(N__12327),
            .I(bZ0Z_9));
    LocalMux I__2595 (
            .O(N__12324),
            .I(bZ0Z_9));
    LocalMux I__2594 (
            .O(N__12319),
            .I(bZ0Z_9));
    Odrv4 I__2593 (
            .O(N__12314),
            .I(bZ0Z_9));
    Odrv4 I__2592 (
            .O(N__12311),
            .I(bZ0Z_9));
    CascadeMux I__2591 (
            .O(N__12296),
            .I(N__12293));
    InMux I__2590 (
            .O(N__12293),
            .I(N__12290));
    LocalMux I__2589 (
            .O(N__12290),
            .I(\ALU.regsA_result_axb_9_l_ofx_2 ));
    InMux I__2588 (
            .O(N__12287),
            .I(N__12283));
    InMux I__2587 (
            .O(N__12286),
            .I(N__12278));
    LocalMux I__2586 (
            .O(N__12283),
            .I(N__12275));
    InMux I__2585 (
            .O(N__12282),
            .I(N__12272));
    InMux I__2584 (
            .O(N__12281),
            .I(N__12268));
    LocalMux I__2583 (
            .O(N__12278),
            .I(N__12261));
    Span4Mux_h I__2582 (
            .O(N__12275),
            .I(N__12261));
    LocalMux I__2581 (
            .O(N__12272),
            .I(N__12261));
    InMux I__2580 (
            .O(N__12271),
            .I(N__12258));
    LocalMux I__2579 (
            .O(N__12268),
            .I(N__12255));
    Span4Mux_v I__2578 (
            .O(N__12261),
            .I(N__12252));
    LocalMux I__2577 (
            .O(N__12258),
            .I(RXbuffer_5));
    Odrv4 I__2576 (
            .O(N__12255),
            .I(RXbuffer_5));
    Odrv4 I__2575 (
            .O(N__12252),
            .I(RXbuffer_5));
    CEMux I__2574 (
            .O(N__12245),
            .I(N__12238));
    CEMux I__2573 (
            .O(N__12244),
            .I(N__12235));
    CEMux I__2572 (
            .O(N__12243),
            .I(N__12232));
    CEMux I__2571 (
            .O(N__12242),
            .I(N__12228));
    CEMux I__2570 (
            .O(N__12241),
            .I(N__12225));
    LocalMux I__2569 (
            .O(N__12238),
            .I(N__12222));
    LocalMux I__2568 (
            .O(N__12235),
            .I(N__12217));
    LocalMux I__2567 (
            .O(N__12232),
            .I(N__12217));
    CEMux I__2566 (
            .O(N__12231),
            .I(N__12214));
    LocalMux I__2565 (
            .O(N__12228),
            .I(N__12210));
    LocalMux I__2564 (
            .O(N__12225),
            .I(N__12207));
    Span4Mux_v I__2563 (
            .O(N__12222),
            .I(N__12200));
    Span4Mux_h I__2562 (
            .O(N__12217),
            .I(N__12200));
    LocalMux I__2561 (
            .O(N__12214),
            .I(N__12200));
    CEMux I__2560 (
            .O(N__12213),
            .I(N__12196));
    Span4Mux_v I__2559 (
            .O(N__12210),
            .I(N__12193));
    Span4Mux_h I__2558 (
            .O(N__12207),
            .I(N__12190));
    Span4Mux_h I__2557 (
            .O(N__12200),
            .I(N__12187));
    CEMux I__2556 (
            .O(N__12199),
            .I(N__12184));
    LocalMux I__2555 (
            .O(N__12196),
            .I(N__12181));
    Span4Mux_h I__2554 (
            .O(N__12193),
            .I(N__12176));
    Span4Mux_v I__2553 (
            .O(N__12190),
            .I(N__12176));
    Span4Mux_h I__2552 (
            .O(N__12187),
            .I(N__12173));
    LocalMux I__2551 (
            .O(N__12184),
            .I(N__12170));
    Span4Mux_h I__2550 (
            .O(N__12181),
            .I(N__12167));
    Odrv4 I__2549 (
            .O(N__12176),
            .I(RXready_RNIICV7_1));
    Odrv4 I__2548 (
            .O(N__12173),
            .I(RXready_RNIICV7_1));
    Odrv12 I__2547 (
            .O(N__12170),
            .I(RXready_RNIICV7_1));
    Odrv4 I__2546 (
            .O(N__12167),
            .I(RXready_RNIICV7_1));
    CascadeMux I__2545 (
            .O(N__12158),
            .I(N__12155));
    InMux I__2544 (
            .O(N__12155),
            .I(N__12152));
    LocalMux I__2543 (
            .O(N__12152),
            .I(N__12149));
    Span4Mux_v I__2542 (
            .O(N__12149),
            .I(N__12146));
    Odrv4 I__2541 (
            .O(N__12146),
            .I(\ALU.regsA_result_cry_1_ma ));
    InMux I__2540 (
            .O(N__12143),
            .I(N__12140));
    LocalMux I__2539 (
            .O(N__12140),
            .I(N__12137));
    Span4Mux_v I__2538 (
            .O(N__12137),
            .I(N__12134));
    Odrv4 I__2537 (
            .O(N__12134),
            .I(\ALU.regsA_result_cry_3_ma_3 ));
    InMux I__2536 (
            .O(N__12131),
            .I(N__12128));
    LocalMux I__2535 (
            .O(N__12128),
            .I(N__12125));
    Span4Mux_h I__2534 (
            .O(N__12125),
            .I(N__12122));
    Odrv4 I__2533 (
            .O(N__12122),
            .I(\ALU.regsA_result_cry_2_ma ));
    InMux I__2532 (
            .O(N__12119),
            .I(N__12116));
    LocalMux I__2531 (
            .O(N__12116),
            .I(N__12111));
    InMux I__2530 (
            .O(N__12115),
            .I(N__12108));
    InMux I__2529 (
            .O(N__12114),
            .I(N__12105));
    Span4Mux_h I__2528 (
            .O(N__12111),
            .I(N__12100));
    LocalMux I__2527 (
            .O(N__12108),
            .I(N__12097));
    LocalMux I__2526 (
            .O(N__12105),
            .I(N__12094));
    InMux I__2525 (
            .O(N__12104),
            .I(N__12091));
    InMux I__2524 (
            .O(N__12103),
            .I(N__12088));
    Span4Mux_h I__2523 (
            .O(N__12100),
            .I(N__12085));
    Sp12to4 I__2522 (
            .O(N__12097),
            .I(N__12082));
    Span4Mux_v I__2521 (
            .O(N__12094),
            .I(N__12077));
    LocalMux I__2520 (
            .O(N__12091),
            .I(N__12077));
    LocalMux I__2519 (
            .O(N__12088),
            .I(RXbuffer_7));
    Odrv4 I__2518 (
            .O(N__12085),
            .I(RXbuffer_7));
    Odrv12 I__2517 (
            .O(N__12082),
            .I(RXbuffer_7));
    Odrv4 I__2516 (
            .O(N__12077),
            .I(RXbuffer_7));
    CascadeMux I__2515 (
            .O(N__12068),
            .I(N__12058));
    CascadeMux I__2514 (
            .O(N__12067),
            .I(N__12054));
    CascadeMux I__2513 (
            .O(N__12066),
            .I(N__12050));
    InMux I__2512 (
            .O(N__12065),
            .I(N__12045));
    InMux I__2511 (
            .O(N__12064),
            .I(N__12040));
    InMux I__2510 (
            .O(N__12063),
            .I(N__12040));
    InMux I__2509 (
            .O(N__12062),
            .I(N__12037));
    CascadeMux I__2508 (
            .O(N__12061),
            .I(N__12030));
    InMux I__2507 (
            .O(N__12058),
            .I(N__12027));
    InMux I__2506 (
            .O(N__12057),
            .I(N__12022));
    InMux I__2505 (
            .O(N__12054),
            .I(N__12019));
    InMux I__2504 (
            .O(N__12053),
            .I(N__12014));
    InMux I__2503 (
            .O(N__12050),
            .I(N__12014));
    InMux I__2502 (
            .O(N__12049),
            .I(N__12010));
    InMux I__2501 (
            .O(N__12048),
            .I(N__12007));
    LocalMux I__2500 (
            .O(N__12045),
            .I(N__12000));
    LocalMux I__2499 (
            .O(N__12040),
            .I(N__12000));
    LocalMux I__2498 (
            .O(N__12037),
            .I(N__12000));
    InMux I__2497 (
            .O(N__12036),
            .I(N__11995));
    InMux I__2496 (
            .O(N__12035),
            .I(N__11995));
    InMux I__2495 (
            .O(N__12034),
            .I(N__11990));
    InMux I__2494 (
            .O(N__12033),
            .I(N__11987));
    InMux I__2493 (
            .O(N__12030),
            .I(N__11984));
    LocalMux I__2492 (
            .O(N__12027),
            .I(N__11981));
    InMux I__2491 (
            .O(N__12026),
            .I(N__11976));
    InMux I__2490 (
            .O(N__12025),
            .I(N__11976));
    LocalMux I__2489 (
            .O(N__12022),
            .I(N__11971));
    LocalMux I__2488 (
            .O(N__12019),
            .I(N__11971));
    LocalMux I__2487 (
            .O(N__12014),
            .I(N__11964));
    InMux I__2486 (
            .O(N__12013),
            .I(N__11961));
    LocalMux I__2485 (
            .O(N__12010),
            .I(N__11952));
    LocalMux I__2484 (
            .O(N__12007),
            .I(N__11952));
    Span4Mux_v I__2483 (
            .O(N__12000),
            .I(N__11952));
    LocalMux I__2482 (
            .O(N__11995),
            .I(N__11952));
    CascadeMux I__2481 (
            .O(N__11994),
            .I(N__11949));
    CascadeMux I__2480 (
            .O(N__11993),
            .I(N__11941));
    LocalMux I__2479 (
            .O(N__11990),
            .I(N__11933));
    LocalMux I__2478 (
            .O(N__11987),
            .I(N__11933));
    LocalMux I__2477 (
            .O(N__11984),
            .I(N__11933));
    Span4Mux_v I__2476 (
            .O(N__11981),
            .I(N__11926));
    LocalMux I__2475 (
            .O(N__11976),
            .I(N__11926));
    Span4Mux_v I__2474 (
            .O(N__11971),
            .I(N__11926));
    InMux I__2473 (
            .O(N__11970),
            .I(N__11923));
    InMux I__2472 (
            .O(N__11969),
            .I(N__11920));
    InMux I__2471 (
            .O(N__11968),
            .I(N__11915));
    InMux I__2470 (
            .O(N__11967),
            .I(N__11915));
    Span4Mux_v I__2469 (
            .O(N__11964),
            .I(N__11908));
    LocalMux I__2468 (
            .O(N__11961),
            .I(N__11908));
    Span4Mux_v I__2467 (
            .O(N__11952),
            .I(N__11908));
    InMux I__2466 (
            .O(N__11949),
            .I(N__11905));
    CascadeMux I__2465 (
            .O(N__11948),
            .I(N__11901));
    CascadeMux I__2464 (
            .O(N__11947),
            .I(N__11898));
    InMux I__2463 (
            .O(N__11946),
            .I(N__11895));
    InMux I__2462 (
            .O(N__11945),
            .I(N__11892));
    InMux I__2461 (
            .O(N__11944),
            .I(N__11887));
    InMux I__2460 (
            .O(N__11941),
            .I(N__11887));
    InMux I__2459 (
            .O(N__11940),
            .I(N__11884));
    Span4Mux_h I__2458 (
            .O(N__11933),
            .I(N__11879));
    Span4Mux_h I__2457 (
            .O(N__11926),
            .I(N__11879));
    LocalMux I__2456 (
            .O(N__11923),
            .I(N__11876));
    LocalMux I__2455 (
            .O(N__11920),
            .I(N__11873));
    LocalMux I__2454 (
            .O(N__11915),
            .I(N__11866));
    Span4Mux_h I__2453 (
            .O(N__11908),
            .I(N__11866));
    LocalMux I__2452 (
            .O(N__11905),
            .I(N__11866));
    InMux I__2451 (
            .O(N__11904),
            .I(N__11859));
    InMux I__2450 (
            .O(N__11901),
            .I(N__11859));
    InMux I__2449 (
            .O(N__11898),
            .I(N__11859));
    LocalMux I__2448 (
            .O(N__11895),
            .I(bZ0Z_1));
    LocalMux I__2447 (
            .O(N__11892),
            .I(bZ0Z_1));
    LocalMux I__2446 (
            .O(N__11887),
            .I(bZ0Z_1));
    LocalMux I__2445 (
            .O(N__11884),
            .I(bZ0Z_1));
    Odrv4 I__2444 (
            .O(N__11879),
            .I(bZ0Z_1));
    Odrv12 I__2443 (
            .O(N__11876),
            .I(bZ0Z_1));
    Odrv4 I__2442 (
            .O(N__11873),
            .I(bZ0Z_1));
    Odrv4 I__2441 (
            .O(N__11866),
            .I(bZ0Z_1));
    LocalMux I__2440 (
            .O(N__11859),
            .I(bZ0Z_1));
    InMux I__2439 (
            .O(N__11840),
            .I(N__11837));
    LocalMux I__2438 (
            .O(N__11837),
            .I(\ALU.regsA_result_cry_2_ma_5 ));
    CascadeMux I__2437 (
            .O(N__11834),
            .I(N__11828));
    InMux I__2436 (
            .O(N__11833),
            .I(N__11821));
    InMux I__2435 (
            .O(N__11832),
            .I(N__11818));
    InMux I__2434 (
            .O(N__11831),
            .I(N__11815));
    InMux I__2433 (
            .O(N__11828),
            .I(N__11811));
    InMux I__2432 (
            .O(N__11827),
            .I(N__11808));
    InMux I__2431 (
            .O(N__11826),
            .I(N__11803));
    InMux I__2430 (
            .O(N__11825),
            .I(N__11803));
    InMux I__2429 (
            .O(N__11824),
            .I(N__11800));
    LocalMux I__2428 (
            .O(N__11821),
            .I(N__11794));
    LocalMux I__2427 (
            .O(N__11818),
            .I(N__11789));
    LocalMux I__2426 (
            .O(N__11815),
            .I(N__11789));
    CascadeMux I__2425 (
            .O(N__11814),
            .I(N__11786));
    LocalMux I__2424 (
            .O(N__11811),
            .I(N__11776));
    LocalMux I__2423 (
            .O(N__11808),
            .I(N__11776));
    LocalMux I__2422 (
            .O(N__11803),
            .I(N__11771));
    LocalMux I__2421 (
            .O(N__11800),
            .I(N__11771));
    InMux I__2420 (
            .O(N__11799),
            .I(N__11766));
    InMux I__2419 (
            .O(N__11798),
            .I(N__11766));
    InMux I__2418 (
            .O(N__11797),
            .I(N__11763));
    Span4Mux_h I__2417 (
            .O(N__11794),
            .I(N__11758));
    Span4Mux_v I__2416 (
            .O(N__11789),
            .I(N__11758));
    InMux I__2415 (
            .O(N__11786),
            .I(N__11753));
    InMux I__2414 (
            .O(N__11785),
            .I(N__11753));
    InMux I__2413 (
            .O(N__11784),
            .I(N__11750));
    InMux I__2412 (
            .O(N__11783),
            .I(N__11743));
    InMux I__2411 (
            .O(N__11782),
            .I(N__11738));
    InMux I__2410 (
            .O(N__11781),
            .I(N__11738));
    Span4Mux_v I__2409 (
            .O(N__11776),
            .I(N__11731));
    Span4Mux_v I__2408 (
            .O(N__11771),
            .I(N__11731));
    LocalMux I__2407 (
            .O(N__11766),
            .I(N__11731));
    LocalMux I__2406 (
            .O(N__11763),
            .I(N__11724));
    Span4Mux_h I__2405 (
            .O(N__11758),
            .I(N__11724));
    LocalMux I__2404 (
            .O(N__11753),
            .I(N__11719));
    LocalMux I__2403 (
            .O(N__11750),
            .I(N__11719));
    InMux I__2402 (
            .O(N__11749),
            .I(N__11716));
    InMux I__2401 (
            .O(N__11748),
            .I(N__11711));
    InMux I__2400 (
            .O(N__11747),
            .I(N__11711));
    InMux I__2399 (
            .O(N__11746),
            .I(N__11708));
    LocalMux I__2398 (
            .O(N__11743),
            .I(N__11705));
    LocalMux I__2397 (
            .O(N__11738),
            .I(N__11700));
    Span4Mux_h I__2396 (
            .O(N__11731),
            .I(N__11700));
    InMux I__2395 (
            .O(N__11730),
            .I(N__11695));
    InMux I__2394 (
            .O(N__11729),
            .I(N__11695));
    Odrv4 I__2393 (
            .O(N__11724),
            .I(bZ0Z_2));
    Odrv12 I__2392 (
            .O(N__11719),
            .I(bZ0Z_2));
    LocalMux I__2391 (
            .O(N__11716),
            .I(bZ0Z_2));
    LocalMux I__2390 (
            .O(N__11711),
            .I(bZ0Z_2));
    LocalMux I__2389 (
            .O(N__11708),
            .I(bZ0Z_2));
    Odrv4 I__2388 (
            .O(N__11705),
            .I(bZ0Z_2));
    Odrv4 I__2387 (
            .O(N__11700),
            .I(bZ0Z_2));
    LocalMux I__2386 (
            .O(N__11695),
            .I(bZ0Z_2));
    InMux I__2385 (
            .O(N__11678),
            .I(N__11675));
    LocalMux I__2384 (
            .O(N__11675),
            .I(\ALU.regsA_result_cry_3_ma_5 ));
    CascadeMux I__2383 (
            .O(N__11672),
            .I(N__11669));
    InMux I__2382 (
            .O(N__11669),
            .I(N__11666));
    LocalMux I__2381 (
            .O(N__11666),
            .I(\ALU.regsA_result_cry_4_ma_4 ));
    CascadeMux I__2380 (
            .O(N__11663),
            .I(N__11654));
    CascadeMux I__2379 (
            .O(N__11662),
            .I(N__11647));
    InMux I__2378 (
            .O(N__11661),
            .I(N__11641));
    InMux I__2377 (
            .O(N__11660),
            .I(N__11638));
    InMux I__2376 (
            .O(N__11659),
            .I(N__11635));
    InMux I__2375 (
            .O(N__11658),
            .I(N__11630));
    InMux I__2374 (
            .O(N__11657),
            .I(N__11630));
    InMux I__2373 (
            .O(N__11654),
            .I(N__11627));
    InMux I__2372 (
            .O(N__11653),
            .I(N__11620));
    InMux I__2371 (
            .O(N__11652),
            .I(N__11620));
    InMux I__2370 (
            .O(N__11651),
            .I(N__11620));
    InMux I__2369 (
            .O(N__11650),
            .I(N__11617));
    InMux I__2368 (
            .O(N__11647),
            .I(N__11612));
    InMux I__2367 (
            .O(N__11646),
            .I(N__11612));
    InMux I__2366 (
            .O(N__11645),
            .I(N__11607));
    InMux I__2365 (
            .O(N__11644),
            .I(N__11603));
    LocalMux I__2364 (
            .O(N__11641),
            .I(N__11595));
    LocalMux I__2363 (
            .O(N__11638),
            .I(N__11595));
    LocalMux I__2362 (
            .O(N__11635),
            .I(N__11595));
    LocalMux I__2361 (
            .O(N__11630),
            .I(N__11592));
    LocalMux I__2360 (
            .O(N__11627),
            .I(N__11587));
    LocalMux I__2359 (
            .O(N__11620),
            .I(N__11587));
    LocalMux I__2358 (
            .O(N__11617),
            .I(N__11580));
    LocalMux I__2357 (
            .O(N__11612),
            .I(N__11580));
    InMux I__2356 (
            .O(N__11611),
            .I(N__11577));
    InMux I__2355 (
            .O(N__11610),
            .I(N__11574));
    LocalMux I__2354 (
            .O(N__11607),
            .I(N__11571));
    InMux I__2353 (
            .O(N__11606),
            .I(N__11568));
    LocalMux I__2352 (
            .O(N__11603),
            .I(N__11565));
    InMux I__2351 (
            .O(N__11602),
            .I(N__11562));
    Span4Mux_v I__2350 (
            .O(N__11595),
            .I(N__11555));
    Span4Mux_v I__2349 (
            .O(N__11592),
            .I(N__11555));
    Span4Mux_v I__2348 (
            .O(N__11587),
            .I(N__11555));
    InMux I__2347 (
            .O(N__11586),
            .I(N__11550));
    InMux I__2346 (
            .O(N__11585),
            .I(N__11550));
    Span4Mux_h I__2345 (
            .O(N__11580),
            .I(N__11547));
    LocalMux I__2344 (
            .O(N__11577),
            .I(N__11542));
    LocalMux I__2343 (
            .O(N__11574),
            .I(N__11542));
    Span4Mux_h I__2342 (
            .O(N__11571),
            .I(N__11535));
    LocalMux I__2341 (
            .O(N__11568),
            .I(N__11535));
    Span4Mux_h I__2340 (
            .O(N__11565),
            .I(N__11535));
    LocalMux I__2339 (
            .O(N__11562),
            .I(bZ0Z_4));
    Odrv4 I__2338 (
            .O(N__11555),
            .I(bZ0Z_4));
    LocalMux I__2337 (
            .O(N__11550),
            .I(bZ0Z_4));
    Odrv4 I__2336 (
            .O(N__11547),
            .I(bZ0Z_4));
    Odrv4 I__2335 (
            .O(N__11542),
            .I(bZ0Z_4));
    Odrv4 I__2334 (
            .O(N__11535),
            .I(bZ0Z_4));
    InMux I__2333 (
            .O(N__11522),
            .I(N__11519));
    LocalMux I__2332 (
            .O(N__11519),
            .I(\ALU.regsA_result_cry_5_ma_4 ));
    CascadeMux I__2331 (
            .O(N__11516),
            .I(\FTDI.N_23_cascade_ ));
    InMux I__2330 (
            .O(N__11513),
            .I(N__11498));
    InMux I__2329 (
            .O(N__11512),
            .I(N__11498));
    InMux I__2328 (
            .O(N__11511),
            .I(N__11498));
    InMux I__2327 (
            .O(N__11510),
            .I(N__11498));
    InMux I__2326 (
            .O(N__11509),
            .I(N__11498));
    LocalMux I__2325 (
            .O(N__11498),
            .I(\FTDI.RXstateZ0Z_0 ));
    CascadeMux I__2324 (
            .O(N__11495),
            .I(N__11485));
    CascadeMux I__2323 (
            .O(N__11494),
            .I(N__11481));
    InMux I__2322 (
            .O(N__11493),
            .I(N__11476));
    InMux I__2321 (
            .O(N__11492),
            .I(N__11476));
    InMux I__2320 (
            .O(N__11491),
            .I(N__11461));
    InMux I__2319 (
            .O(N__11490),
            .I(N__11461));
    InMux I__2318 (
            .O(N__11489),
            .I(N__11461));
    InMux I__2317 (
            .O(N__11488),
            .I(N__11461));
    InMux I__2316 (
            .O(N__11485),
            .I(N__11461));
    InMux I__2315 (
            .O(N__11484),
            .I(N__11461));
    InMux I__2314 (
            .O(N__11481),
            .I(N__11461));
    LocalMux I__2313 (
            .O(N__11476),
            .I(\FTDI.RXstateZ0Z_3 ));
    LocalMux I__2312 (
            .O(N__11461),
            .I(\FTDI.RXstateZ0Z_3 ));
    CascadeMux I__2311 (
            .O(N__11456),
            .I(N__11453));
    InMux I__2310 (
            .O(N__11453),
            .I(N__11444));
    InMux I__2309 (
            .O(N__11452),
            .I(N__11444));
    InMux I__2308 (
            .O(N__11451),
            .I(N__11437));
    InMux I__2307 (
            .O(N__11450),
            .I(N__11437));
    InMux I__2306 (
            .O(N__11449),
            .I(N__11437));
    LocalMux I__2305 (
            .O(N__11444),
            .I(\FTDI.RXstateZ0Z_2 ));
    LocalMux I__2304 (
            .O(N__11437),
            .I(\FTDI.RXstateZ0Z_2 ));
    CascadeMux I__2303 (
            .O(N__11432),
            .I(N__11428));
    InMux I__2302 (
            .O(N__11431),
            .I(N__11423));
    InMux I__2301 (
            .O(N__11428),
            .I(N__11423));
    LocalMux I__2300 (
            .O(N__11423),
            .I(\FTDI.N_28 ));
    InMux I__2299 (
            .O(N__11420),
            .I(N__11410));
    InMux I__2298 (
            .O(N__11419),
            .I(N__11410));
    InMux I__2297 (
            .O(N__11418),
            .I(N__11401));
    InMux I__2296 (
            .O(N__11417),
            .I(N__11401));
    InMux I__2295 (
            .O(N__11416),
            .I(N__11401));
    InMux I__2294 (
            .O(N__11415),
            .I(N__11401));
    LocalMux I__2293 (
            .O(N__11410),
            .I(\FTDI.RXstateZ0Z_1 ));
    LocalMux I__2292 (
            .O(N__11401),
            .I(\FTDI.RXstateZ0Z_1 ));
    CEMux I__2291 (
            .O(N__11396),
            .I(N__11391));
    CEMux I__2290 (
            .O(N__11395),
            .I(N__11388));
    CEMux I__2289 (
            .O(N__11394),
            .I(N__11384));
    LocalMux I__2288 (
            .O(N__11391),
            .I(N__11381));
    LocalMux I__2287 (
            .O(N__11388),
            .I(N__11378));
    CEMux I__2286 (
            .O(N__11387),
            .I(N__11375));
    LocalMux I__2285 (
            .O(N__11384),
            .I(N__11371));
    Span4Mux_v I__2284 (
            .O(N__11381),
            .I(N__11368));
    Span4Mux_h I__2283 (
            .O(N__11378),
            .I(N__11363));
    LocalMux I__2282 (
            .O(N__11375),
            .I(N__11363));
    CEMux I__2281 (
            .O(N__11374),
            .I(N__11360));
    Span4Mux_h I__2280 (
            .O(N__11371),
            .I(N__11357));
    Span4Mux_h I__2279 (
            .O(N__11368),
            .I(N__11354));
    Span4Mux_v I__2278 (
            .O(N__11363),
            .I(N__11349));
    LocalMux I__2277 (
            .O(N__11360),
            .I(N__11349));
    Span4Mux_h I__2276 (
            .O(N__11357),
            .I(N__11346));
    Span4Mux_h I__2275 (
            .O(N__11354),
            .I(N__11341));
    Span4Mux_v I__2274 (
            .O(N__11349),
            .I(N__11341));
    Odrv4 I__2273 (
            .O(N__11346),
            .I(RXready_RNIICV7_0));
    Odrv4 I__2272 (
            .O(N__11341),
            .I(RXready_RNIICV7_0));
    InMux I__2271 (
            .O(N__11336),
            .I(N__11333));
    LocalMux I__2270 (
            .O(N__11333),
            .I(N__11328));
    InMux I__2269 (
            .O(N__11332),
            .I(N__11325));
    InMux I__2268 (
            .O(N__11331),
            .I(N__11322));
    Span4Mux_v I__2267 (
            .O(N__11328),
            .I(N__11315));
    LocalMux I__2266 (
            .O(N__11325),
            .I(N__11315));
    LocalMux I__2265 (
            .O(N__11322),
            .I(N__11311));
    InMux I__2264 (
            .O(N__11321),
            .I(N__11308));
    InMux I__2263 (
            .O(N__11320),
            .I(N__11305));
    Span4Mux_h I__2262 (
            .O(N__11315),
            .I(N__11302));
    InMux I__2261 (
            .O(N__11314),
            .I(N__11299));
    Span4Mux_v I__2260 (
            .O(N__11311),
            .I(N__11294));
    LocalMux I__2259 (
            .O(N__11308),
            .I(N__11294));
    LocalMux I__2258 (
            .O(N__11305),
            .I(RXbuffer_1));
    Odrv4 I__2257 (
            .O(N__11302),
            .I(RXbuffer_1));
    LocalMux I__2256 (
            .O(N__11299),
            .I(RXbuffer_1));
    Odrv4 I__2255 (
            .O(N__11294),
            .I(RXbuffer_1));
    CascadeMux I__2254 (
            .O(N__11285),
            .I(N__11273));
    InMux I__2253 (
            .O(N__11284),
            .I(N__11266));
    InMux I__2252 (
            .O(N__11283),
            .I(N__11266));
    InMux I__2251 (
            .O(N__11282),
            .I(N__11257));
    InMux I__2250 (
            .O(N__11281),
            .I(N__11257));
    InMux I__2249 (
            .O(N__11280),
            .I(N__11257));
    InMux I__2248 (
            .O(N__11279),
            .I(N__11254));
    InMux I__2247 (
            .O(N__11278),
            .I(N__11241));
    InMux I__2246 (
            .O(N__11277),
            .I(N__11241));
    InMux I__2245 (
            .O(N__11276),
            .I(N__11241));
    InMux I__2244 (
            .O(N__11273),
            .I(N__11241));
    InMux I__2243 (
            .O(N__11272),
            .I(N__11241));
    InMux I__2242 (
            .O(N__11271),
            .I(N__11241));
    LocalMux I__2241 (
            .O(N__11266),
            .I(N__11238));
    InMux I__2240 (
            .O(N__11265),
            .I(N__11235));
    InMux I__2239 (
            .O(N__11264),
            .I(N__11232));
    LocalMux I__2238 (
            .O(N__11257),
            .I(N__11223));
    LocalMux I__2237 (
            .O(N__11254),
            .I(N__11223));
    LocalMux I__2236 (
            .O(N__11241),
            .I(N__11223));
    Span4Mux_h I__2235 (
            .O(N__11238),
            .I(N__11216));
    LocalMux I__2234 (
            .O(N__11235),
            .I(N__11216));
    LocalMux I__2233 (
            .O(N__11232),
            .I(N__11216));
    InMux I__2232 (
            .O(N__11231),
            .I(N__11213));
    InMux I__2231 (
            .O(N__11230),
            .I(N__11210));
    Span4Mux_v I__2230 (
            .O(N__11223),
            .I(N__11207));
    Span4Mux_v I__2229 (
            .O(N__11216),
            .I(N__11204));
    LocalMux I__2228 (
            .O(N__11213),
            .I(N__11197));
    LocalMux I__2227 (
            .O(N__11210),
            .I(N__11197));
    Span4Mux_h I__2226 (
            .O(N__11207),
            .I(N__11194));
    Span4Mux_h I__2225 (
            .O(N__11204),
            .I(N__11191));
    InMux I__2224 (
            .O(N__11203),
            .I(N__11186));
    InMux I__2223 (
            .O(N__11202),
            .I(N__11186));
    Span4Mux_h I__2222 (
            .O(N__11197),
            .I(N__11181));
    Span4Mux_h I__2221 (
            .O(N__11194),
            .I(N__11181));
    Odrv4 I__2220 (
            .O(N__11191),
            .I(opZ0Z_1));
    LocalMux I__2219 (
            .O(N__11186),
            .I(opZ0Z_1));
    Odrv4 I__2218 (
            .O(N__11181),
            .I(opZ0Z_1));
    InMux I__2217 (
            .O(N__11174),
            .I(N__11171));
    LocalMux I__2216 (
            .O(N__11171),
            .I(N__11168));
    Span4Mux_h I__2215 (
            .O(N__11168),
            .I(N__11165));
    Span4Mux_h I__2214 (
            .O(N__11165),
            .I(N__11162));
    Odrv4 I__2213 (
            .O(N__11162),
            .I(\ALU.addsub_4 ));
    InMux I__2212 (
            .O(N__11159),
            .I(N__11156));
    LocalMux I__2211 (
            .O(N__11156),
            .I(\ALU.mult_4 ));
    InMux I__2210 (
            .O(N__11153),
            .I(N__11150));
    LocalMux I__2209 (
            .O(N__11150),
            .I(N__11147));
    Sp12to4 I__2208 (
            .O(N__11147),
            .I(N__11144));
    Span12Mux_v I__2207 (
            .O(N__11144),
            .I(N__11141));
    Odrv12 I__2206 (
            .O(N__11141),
            .I(res_4));
    InMux I__2205 (
            .O(N__11138),
            .I(N__11135));
    LocalMux I__2204 (
            .O(N__11135),
            .I(N__11132));
    Span12Mux_v I__2203 (
            .O(N__11132),
            .I(N__11129));
    Odrv12 I__2202 (
            .O(N__11129),
            .I(\ALU.regsA_result_cry_2_ma_0 ));
    CascadeMux I__2201 (
            .O(N__11126),
            .I(N__11123));
    InMux I__2200 (
            .O(N__11123),
            .I(N__11120));
    LocalMux I__2199 (
            .O(N__11120),
            .I(N__11117));
    Span4Mux_h I__2198 (
            .O(N__11117),
            .I(N__11114));
    Span4Mux_v I__2197 (
            .O(N__11114),
            .I(N__11111));
    Odrv4 I__2196 (
            .O(N__11111),
            .I(\ALU.regsA_result_cry_10_ma_1 ));
    InMux I__2195 (
            .O(N__11108),
            .I(N__11100));
    InMux I__2194 (
            .O(N__11107),
            .I(N__11100));
    InMux I__2193 (
            .O(N__11106),
            .I(N__11096));
    InMux I__2192 (
            .O(N__11105),
            .I(N__11091));
    LocalMux I__2191 (
            .O(N__11100),
            .I(N__11088));
    InMux I__2190 (
            .O(N__11099),
            .I(N__11085));
    LocalMux I__2189 (
            .O(N__11096),
            .I(N__11081));
    InMux I__2188 (
            .O(N__11095),
            .I(N__11078));
    InMux I__2187 (
            .O(N__11094),
            .I(N__11075));
    LocalMux I__2186 (
            .O(N__11091),
            .I(N__11072));
    Span12Mux_h I__2185 (
            .O(N__11088),
            .I(N__11067));
    LocalMux I__2184 (
            .O(N__11085),
            .I(N__11067));
    InMux I__2183 (
            .O(N__11084),
            .I(N__11064));
    Span4Mux_h I__2182 (
            .O(N__11081),
            .I(N__11061));
    LocalMux I__2181 (
            .O(N__11078),
            .I(N__11058));
    LocalMux I__2180 (
            .O(N__11075),
            .I(N__11053));
    Span4Mux_h I__2179 (
            .O(N__11072),
            .I(N__11053));
    Span12Mux_v I__2178 (
            .O(N__11067),
            .I(N__11050));
    LocalMux I__2177 (
            .O(N__11064),
            .I(RXbuffer_2));
    Odrv4 I__2176 (
            .O(N__11061),
            .I(RXbuffer_2));
    Odrv12 I__2175 (
            .O(N__11058),
            .I(RXbuffer_2));
    Odrv4 I__2174 (
            .O(N__11053),
            .I(RXbuffer_2));
    Odrv12 I__2173 (
            .O(N__11050),
            .I(RXbuffer_2));
    InMux I__2172 (
            .O(N__11039),
            .I(N__11036));
    LocalMux I__2171 (
            .O(N__11036),
            .I(N__11033));
    Odrv12 I__2170 (
            .O(N__11033),
            .I(TXbufferZ0Z_7));
    InMux I__2169 (
            .O(N__11030),
            .I(N__11027));
    LocalMux I__2168 (
            .O(N__11027),
            .I(\FTDI.TXshiftZ0Z_7 ));
    InMux I__2167 (
            .O(N__11024),
            .I(N__11020));
    InMux I__2166 (
            .O(N__11023),
            .I(N__11017));
    LocalMux I__2165 (
            .O(N__11020),
            .I(N__11012));
    LocalMux I__2164 (
            .O(N__11017),
            .I(N__11012));
    Span4Mux_h I__2163 (
            .O(N__11012),
            .I(N__11009));
    Span4Mux_h I__2162 (
            .O(N__11009),
            .I(N__11006));
    Span4Mux_v I__2161 (
            .O(N__11006),
            .I(N__11003));
    Odrv4 I__2160 (
            .O(N__11003),
            .I(RX_c));
    CascadeMux I__2159 (
            .O(N__11000),
            .I(\FTDI.m13_ns_1_cascade_ ));
    CEMux I__2158 (
            .O(N__10997),
            .I(N__10994));
    LocalMux I__2157 (
            .O(N__10994),
            .I(N__10990));
    CEMux I__2156 (
            .O(N__10993),
            .I(N__10987));
    Span4Mux_v I__2155 (
            .O(N__10990),
            .I(N__10984));
    LocalMux I__2154 (
            .O(N__10987),
            .I(N__10981));
    Span4Mux_h I__2153 (
            .O(N__10984),
            .I(N__10978));
    Span4Mux_h I__2152 (
            .O(N__10981),
            .I(N__10975));
    Odrv4 I__2151 (
            .O(N__10978),
            .I(\FTDI.N_201_2 ));
    Odrv4 I__2150 (
            .O(N__10975),
            .I(\FTDI.N_201_2 ));
    InMux I__2149 (
            .O(N__10970),
            .I(N__10967));
    LocalMux I__2148 (
            .O(N__10967),
            .I(N__10964));
    Span4Mux_v I__2147 (
            .O(N__10964),
            .I(N__10960));
    InMux I__2146 (
            .O(N__10963),
            .I(N__10957));
    Span4Mux_h I__2145 (
            .O(N__10960),
            .I(N__10950));
    LocalMux I__2144 (
            .O(N__10957),
            .I(N__10950));
    InMux I__2143 (
            .O(N__10956),
            .I(N__10947));
    InMux I__2142 (
            .O(N__10955),
            .I(N__10944));
    Span4Mux_v I__2141 (
            .O(N__10950),
            .I(N__10939));
    LocalMux I__2140 (
            .O(N__10947),
            .I(N__10936));
    LocalMux I__2139 (
            .O(N__10944),
            .I(N__10933));
    InMux I__2138 (
            .O(N__10943),
            .I(N__10930));
    InMux I__2137 (
            .O(N__10942),
            .I(N__10927));
    Span4Mux_h I__2136 (
            .O(N__10939),
            .I(N__10924));
    Span4Mux_v I__2135 (
            .O(N__10936),
            .I(N__10917));
    Span4Mux_h I__2134 (
            .O(N__10933),
            .I(N__10917));
    LocalMux I__2133 (
            .O(N__10930),
            .I(N__10917));
    LocalMux I__2132 (
            .O(N__10927),
            .I(RXbuffer_4));
    Odrv4 I__2131 (
            .O(N__10924),
            .I(RXbuffer_4));
    Odrv4 I__2130 (
            .O(N__10917),
            .I(RXbuffer_4));
    CascadeMux I__2129 (
            .O(N__10910),
            .I(N__10907));
    InMux I__2128 (
            .O(N__10907),
            .I(N__10904));
    LocalMux I__2127 (
            .O(N__10904),
            .I(\ALU.regsA_result_axb_5_l_ofx_2 ));
    InMux I__2126 (
            .O(N__10901),
            .I(N__10898));
    LocalMux I__2125 (
            .O(N__10898),
            .I(N__10895));
    Span4Mux_h I__2124 (
            .O(N__10895),
            .I(N__10892));
    Odrv4 I__2123 (
            .O(N__10892),
            .I(\ALU.addsub_axb_4_l_ofxZ0 ));
    InMux I__2122 (
            .O(N__10889),
            .I(N__10886));
    LocalMux I__2121 (
            .O(N__10886),
            .I(\ALU.regsA_result_cry_4_ma_2 ));
    InMux I__2120 (
            .O(N__10883),
            .I(N__10880));
    LocalMux I__2119 (
            .O(N__10880),
            .I(\ALU.regsA_result_cry_5_ma_2 ));
    InMux I__2118 (
            .O(N__10877),
            .I(N__10874));
    LocalMux I__2117 (
            .O(N__10874),
            .I(\ALU.regsA_result_cry_6_ma_1 ));
    CascadeMux I__2116 (
            .O(N__10871),
            .I(N__10868));
    InMux I__2115 (
            .O(N__10868),
            .I(N__10865));
    LocalMux I__2114 (
            .O(N__10865),
            .I(N__10862));
    Span4Mux_h I__2113 (
            .O(N__10862),
            .I(N__10859));
    Odrv4 I__2112 (
            .O(N__10859),
            .I(\ALU.regsA_result_axb_9_l_ofx ));
    CascadeMux I__2111 (
            .O(N__10856),
            .I(N__10853));
    InMux I__2110 (
            .O(N__10853),
            .I(N__10849));
    InMux I__2109 (
            .O(N__10852),
            .I(N__10844));
    LocalMux I__2108 (
            .O(N__10849),
            .I(N__10840));
    CascadeMux I__2107 (
            .O(N__10848),
            .I(N__10837));
    CascadeMux I__2106 (
            .O(N__10847),
            .I(N__10834));
    LocalMux I__2105 (
            .O(N__10844),
            .I(N__10830));
    CascadeMux I__2104 (
            .O(N__10843),
            .I(N__10824));
    Span4Mux_v I__2103 (
            .O(N__10840),
            .I(N__10819));
    InMux I__2102 (
            .O(N__10837),
            .I(N__10814));
    InMux I__2101 (
            .O(N__10834),
            .I(N__10814));
    InMux I__2100 (
            .O(N__10833),
            .I(N__10811));
    Span4Mux_v I__2099 (
            .O(N__10830),
            .I(N__10808));
    InMux I__2098 (
            .O(N__10829),
            .I(N__10803));
    InMux I__2097 (
            .O(N__10828),
            .I(N__10803));
    InMux I__2096 (
            .O(N__10827),
            .I(N__10800));
    InMux I__2095 (
            .O(N__10824),
            .I(N__10793));
    InMux I__2094 (
            .O(N__10823),
            .I(N__10793));
    InMux I__2093 (
            .O(N__10822),
            .I(N__10793));
    Span4Mux_h I__2092 (
            .O(N__10819),
            .I(N__10786));
    LocalMux I__2091 (
            .O(N__10814),
            .I(N__10786));
    LocalMux I__2090 (
            .O(N__10811),
            .I(N__10786));
    Odrv4 I__2089 (
            .O(N__10808),
            .I(aZ0Z_4));
    LocalMux I__2088 (
            .O(N__10803),
            .I(aZ0Z_4));
    LocalMux I__2087 (
            .O(N__10800),
            .I(aZ0Z_4));
    LocalMux I__2086 (
            .O(N__10793),
            .I(aZ0Z_4));
    Odrv4 I__2085 (
            .O(N__10786),
            .I(aZ0Z_4));
    CascadeMux I__2084 (
            .O(N__10775),
            .I(N__10772));
    InMux I__2083 (
            .O(N__10772),
            .I(N__10769));
    LocalMux I__2082 (
            .O(N__10769),
            .I(\ALU.regsA_result_axb_9_l_ofx_0 ));
    CascadeMux I__2081 (
            .O(N__10766),
            .I(N__10763));
    InMux I__2080 (
            .O(N__10763),
            .I(N__10760));
    LocalMux I__2079 (
            .O(N__10760),
            .I(N__10757));
    Span4Mux_h I__2078 (
            .O(N__10757),
            .I(N__10754));
    Odrv4 I__2077 (
            .O(N__10754),
            .I(\ALU.mult_AdderTree2_bigtree_642 ));
    InMux I__2076 (
            .O(N__10751),
            .I(bfn_15_14_0_));
    InMux I__2075 (
            .O(N__10748),
            .I(\ALU.regsA_result_cry_9 ));
    InMux I__2074 (
            .O(N__10745),
            .I(N__10742));
    LocalMux I__2073 (
            .O(N__10742),
            .I(N__10739));
    Odrv4 I__2072 (
            .O(N__10739),
            .I(\ALU.regsA_result_cry_9_THRU_CO ));
    InMux I__2071 (
            .O(N__10736),
            .I(N__10733));
    LocalMux I__2070 (
            .O(N__10733),
            .I(N__10730));
    Span4Mux_v I__2069 (
            .O(N__10730),
            .I(N__10727));
    Odrv4 I__2068 (
            .O(N__10727),
            .I(\ALU.regsA_result_cry_9_ma_0 ));
    CascadeMux I__2067 (
            .O(N__10724),
            .I(N__10721));
    InMux I__2066 (
            .O(N__10721),
            .I(N__10718));
    LocalMux I__2065 (
            .O(N__10718),
            .I(\ALU.regsA_result_cry_2_ma_3 ));
    InMux I__2064 (
            .O(N__10715),
            .I(N__10712));
    LocalMux I__2063 (
            .O(N__10712),
            .I(\ALU.regsA_result_cry_7_ma_1 ));
    InMux I__2062 (
            .O(N__10709),
            .I(N__10706));
    LocalMux I__2061 (
            .O(N__10706),
            .I(N__10703));
    Odrv4 I__2060 (
            .O(N__10703),
            .I(\ALU.regsA_result_axb_10 ));
    CascadeMux I__2059 (
            .O(N__10700),
            .I(N__10697));
    InMux I__2058 (
            .O(N__10697),
            .I(N__10694));
    LocalMux I__2057 (
            .O(N__10694),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_4 ));
    InMux I__2056 (
            .O(N__10691),
            .I(N__10688));
    LocalMux I__2055 (
            .O(N__10688),
            .I(N__10685));
    Odrv4 I__2054 (
            .O(N__10685),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_6 ));
    CascadeMux I__2053 (
            .O(N__10682),
            .I(N__10679));
    InMux I__2052 (
            .O(N__10679),
            .I(N__10676));
    LocalMux I__2051 (
            .O(N__10676),
            .I(\ALU.regsA_result_axb_4_l_ofx_2 ));
    CascadeMux I__2050 (
            .O(N__10673),
            .I(N__10670));
    InMux I__2049 (
            .O(N__10670),
            .I(N__10667));
    LocalMux I__2048 (
            .O(N__10667),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_5 ));
    CascadeMux I__2047 (
            .O(N__10664),
            .I(N__10661));
    InMux I__2046 (
            .O(N__10661),
            .I(N__10658));
    LocalMux I__2045 (
            .O(N__10658),
            .I(\ALU.regsA_result_axb_2_l_ofx_5 ));
    InMux I__2044 (
            .O(N__10655),
            .I(N__10652));
    LocalMux I__2043 (
            .O(N__10652),
            .I(N__10649));
    Span4Mux_h I__2042 (
            .O(N__10649),
            .I(N__10646));
    Odrv4 I__2041 (
            .O(N__10646),
            .I(\ALU.mult_AdderTree2_bigtree_635 ));
    InMux I__2040 (
            .O(N__10643),
            .I(\ALU.regsA_result_cry_1_9 ));
    CascadeMux I__2039 (
            .O(N__10640),
            .I(N__10637));
    InMux I__2038 (
            .O(N__10637),
            .I(N__10634));
    LocalMux I__2037 (
            .O(N__10634),
            .I(\ALU.regsA_result_axb_3_l_ofx_5 ));
    InMux I__2036 (
            .O(N__10631),
            .I(N__10628));
    LocalMux I__2035 (
            .O(N__10628),
            .I(N__10625));
    Span4Mux_v I__2034 (
            .O(N__10625),
            .I(N__10622));
    Odrv4 I__2033 (
            .O(N__10622),
            .I(\ALU.mult_AdderTree2_bigtree_636 ));
    InMux I__2032 (
            .O(N__10619),
            .I(\ALU.regsA_result_cry_2_11 ));
    InMux I__2031 (
            .O(N__10616),
            .I(N__10613));
    LocalMux I__2030 (
            .O(N__10613),
            .I(\ALU.regsA_result_axb_4_l_ofx_4 ));
    InMux I__2029 (
            .O(N__10610),
            .I(N__10607));
    LocalMux I__2028 (
            .O(N__10607),
            .I(N__10604));
    Span4Mux_v I__2027 (
            .O(N__10604),
            .I(N__10601));
    Odrv4 I__2026 (
            .O(N__10601),
            .I(\ALU.mult_AdderTree2_bigtree_637 ));
    InMux I__2025 (
            .O(N__10598),
            .I(\ALU.regsA_result_cry_3_11 ));
    CascadeMux I__2024 (
            .O(N__10595),
            .I(N__10592));
    InMux I__2023 (
            .O(N__10592),
            .I(N__10589));
    LocalMux I__2022 (
            .O(N__10589),
            .I(\ALU.regsA_result_axb_5_l_ofx_4 ));
    InMux I__2021 (
            .O(N__10586),
            .I(N__10583));
    LocalMux I__2020 (
            .O(N__10583),
            .I(N__10580));
    Span4Mux_h I__2019 (
            .O(N__10580),
            .I(N__10577));
    Odrv4 I__2018 (
            .O(N__10577),
            .I(\ALU.mult_AdderTree2_bigtree_638 ));
    InMux I__2017 (
            .O(N__10574),
            .I(\ALU.regsA_result_cry_4_10 ));
    CascadeMux I__2016 (
            .O(N__10571),
            .I(N__10568));
    InMux I__2015 (
            .O(N__10568),
            .I(N__10565));
    LocalMux I__2014 (
            .O(N__10565),
            .I(\ALU.regsA_result_axb_6_l_ofx_3 ));
    InMux I__2013 (
            .O(N__10562),
            .I(N__10559));
    LocalMux I__2012 (
            .O(N__10559),
            .I(N__10556));
    Span4Mux_h I__2011 (
            .O(N__10556),
            .I(N__10553));
    Odrv4 I__2010 (
            .O(N__10553),
            .I(\ALU.mult_AdderTree2_bigtree_639 ));
    InMux I__2009 (
            .O(N__10550),
            .I(\ALU.regsA_result_cry_5_10 ));
    CascadeMux I__2008 (
            .O(N__10547),
            .I(N__10544));
    InMux I__2007 (
            .O(N__10544),
            .I(N__10541));
    LocalMux I__2006 (
            .O(N__10541),
            .I(\ALU.regsA_result_axb_7_l_ofx_3 ));
    InMux I__2005 (
            .O(N__10538),
            .I(N__10535));
    LocalMux I__2004 (
            .O(N__10535),
            .I(N__10532));
    Span4Mux_h I__2003 (
            .O(N__10532),
            .I(N__10529));
    Odrv4 I__2002 (
            .O(N__10529),
            .I(\ALU.mult_AdderTree2_bigtree_640 ));
    InMux I__2001 (
            .O(N__10526),
            .I(\ALU.regsA_result_cry_6_9 ));
    CascadeMux I__2000 (
            .O(N__10523),
            .I(N__10520));
    InMux I__1999 (
            .O(N__10520),
            .I(N__10517));
    LocalMux I__1998 (
            .O(N__10517),
            .I(N__10514));
    Span4Mux_h I__1997 (
            .O(N__10514),
            .I(N__10511));
    Odrv4 I__1996 (
            .O(N__10511),
            .I(\ALU.mult_AdderTree2_bigtree_641 ));
    InMux I__1995 (
            .O(N__10508),
            .I(\ALU.regsA_result_cry_7_8 ));
    InMux I__1994 (
            .O(N__10505),
            .I(N__10500));
    CascadeMux I__1993 (
            .O(N__10504),
            .I(N__10496));
    CascadeMux I__1992 (
            .O(N__10503),
            .I(N__10492));
    LocalMux I__1991 (
            .O(N__10500),
            .I(N__10488));
    InMux I__1990 (
            .O(N__10499),
            .I(N__10477));
    InMux I__1989 (
            .O(N__10496),
            .I(N__10477));
    InMux I__1988 (
            .O(N__10495),
            .I(N__10477));
    InMux I__1987 (
            .O(N__10492),
            .I(N__10477));
    InMux I__1986 (
            .O(N__10491),
            .I(N__10477));
    Odrv4 I__1985 (
            .O(N__10488),
            .I(a_fastZ0Z_4));
    LocalMux I__1984 (
            .O(N__10477),
            .I(a_fastZ0Z_4));
    CascadeMux I__1983 (
            .O(N__10472),
            .I(N__10467));
    InMux I__1982 (
            .O(N__10471),
            .I(N__10462));
    InMux I__1981 (
            .O(N__10470),
            .I(N__10462));
    InMux I__1980 (
            .O(N__10467),
            .I(N__10459));
    LocalMux I__1979 (
            .O(N__10462),
            .I(N__10456));
    LocalMux I__1978 (
            .O(N__10459),
            .I(N__10453));
    Span4Mux_v I__1977 (
            .O(N__10456),
            .I(N__10448));
    Span4Mux_v I__1976 (
            .O(N__10453),
            .I(N__10448));
    Odrv4 I__1975 (
            .O(N__10448),
            .I(\ALU.mult_AdderTree2_bigtree_796 ));
    InMux I__1974 (
            .O(N__10445),
            .I(N__10442));
    LocalMux I__1973 (
            .O(N__10442),
            .I(N__10439));
    Span4Mux_v I__1972 (
            .O(N__10439),
            .I(N__10436));
    Span4Mux_h I__1971 (
            .O(N__10436),
            .I(N__10433));
    Span4Mux_h I__1970 (
            .O(N__10433),
            .I(N__10430));
    Odrv4 I__1969 (
            .O(N__10430),
            .I(\ALU.mult_AdderTree2_bigtree_634 ));
    InMux I__1968 (
            .O(N__10427),
            .I(N__10424));
    LocalMux I__1967 (
            .O(N__10424),
            .I(N__10421));
    Span4Mux_v I__1966 (
            .O(N__10421),
            .I(N__10414));
    InMux I__1965 (
            .O(N__10420),
            .I(N__10411));
    InMux I__1964 (
            .O(N__10419),
            .I(N__10408));
    InMux I__1963 (
            .O(N__10418),
            .I(N__10405));
    InMux I__1962 (
            .O(N__10417),
            .I(N__10402));
    Span4Mux_h I__1961 (
            .O(N__10414),
            .I(N__10395));
    LocalMux I__1960 (
            .O(N__10411),
            .I(N__10395));
    LocalMux I__1959 (
            .O(N__10408),
            .I(N__10395));
    LocalMux I__1958 (
            .O(N__10405),
            .I(RXbuffer_3));
    LocalMux I__1957 (
            .O(N__10402),
            .I(RXbuffer_3));
    Odrv4 I__1956 (
            .O(N__10395),
            .I(RXbuffer_3));
    CascadeMux I__1955 (
            .O(N__10388),
            .I(N__10385));
    InMux I__1954 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__1953 (
            .O(N__10382),
            .I(N__10379));
    Span4Mux_v I__1952 (
            .O(N__10379),
            .I(N__10376));
    Span4Mux_h I__1951 (
            .O(N__10376),
            .I(N__10373));
    Odrv4 I__1950 (
            .O(N__10373),
            .I(\ALU.mult_AdderTree2_bigtree_599 ));
    InMux I__1949 (
            .O(N__10370),
            .I(N__10367));
    LocalMux I__1948 (
            .O(N__10367),
            .I(N__10364));
    Span4Mux_v I__1947 (
            .O(N__10364),
            .I(N__10361));
    Odrv4 I__1946 (
            .O(N__10361),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_3 ));
    InMux I__1945 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__1944 (
            .O(N__10355),
            .I(N__10352));
    Span4Mux_v I__1943 (
            .O(N__10352),
            .I(N__10349));
    Odrv4 I__1942 (
            .O(N__10349),
            .I(\ALU.regsA_result_axb_2_l_ofx_3 ));
    CascadeMux I__1941 (
            .O(N__10346),
            .I(N__10343));
    InMux I__1940 (
            .O(N__10343),
            .I(N__10340));
    LocalMux I__1939 (
            .O(N__10340),
            .I(N__10337));
    Span4Mux_v I__1938 (
            .O(N__10337),
            .I(N__10334));
    Odrv4 I__1937 (
            .O(N__10334),
            .I(\ALU.regsA_result_axb_3_l_ofx_3 ));
    InMux I__1936 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__1935 (
            .O(N__10328),
            .I(N__10325));
    Span4Mux_v I__1934 (
            .O(N__10325),
            .I(N__10322));
    Odrv4 I__1933 (
            .O(N__10322),
            .I(\ALU.regsA_result_cry_0_c_RNO ));
    InMux I__1932 (
            .O(N__10319),
            .I(N__10316));
    LocalMux I__1931 (
            .O(N__10316),
            .I(\FTDI.TXshiftZ0Z_6 ));
    InMux I__1930 (
            .O(N__10313),
            .I(N__10310));
    LocalMux I__1929 (
            .O(N__10310),
            .I(N__10307));
    Odrv4 I__1928 (
            .O(N__10307),
            .I(TXbufferZ0Z_5));
    InMux I__1927 (
            .O(N__10304),
            .I(N__10301));
    LocalMux I__1926 (
            .O(N__10301),
            .I(\FTDI.TXshiftZ0Z_5 ));
    InMux I__1925 (
            .O(N__10298),
            .I(N__10295));
    LocalMux I__1924 (
            .O(N__10295),
            .I(\ALU.regsA_result_cry_11_ma_0 ));
    InMux I__1923 (
            .O(N__10292),
            .I(N__10288));
    CascadeMux I__1922 (
            .O(N__10291),
            .I(N__10283));
    LocalMux I__1921 (
            .O(N__10288),
            .I(N__10280));
    InMux I__1920 (
            .O(N__10287),
            .I(N__10277));
    CascadeMux I__1919 (
            .O(N__10286),
            .I(N__10272));
    InMux I__1918 (
            .O(N__10283),
            .I(N__10268));
    Span4Mux_v I__1917 (
            .O(N__10280),
            .I(N__10263));
    LocalMux I__1916 (
            .O(N__10277),
            .I(N__10263));
    CascadeMux I__1915 (
            .O(N__10276),
            .I(N__10259));
    InMux I__1914 (
            .O(N__10275),
            .I(N__10255));
    InMux I__1913 (
            .O(N__10272),
            .I(N__10250));
    InMux I__1912 (
            .O(N__10271),
            .I(N__10250));
    LocalMux I__1911 (
            .O(N__10268),
            .I(N__10247));
    Span4Mux_v I__1910 (
            .O(N__10263),
            .I(N__10244));
    InMux I__1909 (
            .O(N__10262),
            .I(N__10237));
    InMux I__1908 (
            .O(N__10259),
            .I(N__10237));
    InMux I__1907 (
            .O(N__10258),
            .I(N__10237));
    LocalMux I__1906 (
            .O(N__10255),
            .I(bZ0Z_11));
    LocalMux I__1905 (
            .O(N__10250),
            .I(bZ0Z_11));
    Odrv12 I__1904 (
            .O(N__10247),
            .I(bZ0Z_11));
    Odrv4 I__1903 (
            .O(N__10244),
            .I(bZ0Z_11));
    LocalMux I__1902 (
            .O(N__10237),
            .I(bZ0Z_11));
    CascadeMux I__1901 (
            .O(N__10226),
            .I(N__10223));
    InMux I__1900 (
            .O(N__10223),
            .I(N__10220));
    LocalMux I__1899 (
            .O(N__10220),
            .I(\ALU.regsA_result_axb_11_l_ofx_0 ));
    InMux I__1898 (
            .O(N__10217),
            .I(N__10214));
    LocalMux I__1897 (
            .O(N__10214),
            .I(\ALU.regsA_result_cry_10_ma_0 ));
    InMux I__1896 (
            .O(N__10211),
            .I(N__10208));
    LocalMux I__1895 (
            .O(N__10208),
            .I(TXbufferZ0Z_1));
    InMux I__1894 (
            .O(N__10205),
            .I(N__10202));
    LocalMux I__1893 (
            .O(N__10202),
            .I(N__10199));
    Odrv4 I__1892 (
            .O(N__10199),
            .I(TXbufferZ0Z_2));
    InMux I__1891 (
            .O(N__10196),
            .I(N__10193));
    LocalMux I__1890 (
            .O(N__10193),
            .I(\FTDI.TXshiftZ0Z_2 ));
    InMux I__1889 (
            .O(N__10190),
            .I(N__10187));
    LocalMux I__1888 (
            .O(N__10187),
            .I(N__10184));
    Odrv4 I__1887 (
            .O(N__10184),
            .I(TXbufferZ0Z_6));
    InMux I__1886 (
            .O(N__10181),
            .I(N__10178));
    LocalMux I__1885 (
            .O(N__10178),
            .I(TXbufferZ0Z_4));
    InMux I__1884 (
            .O(N__10175),
            .I(N__10172));
    LocalMux I__1883 (
            .O(N__10172),
            .I(\FTDI.TXshiftZ0Z_1 ));
    InMux I__1882 (
            .O(N__10169),
            .I(N__10166));
    LocalMux I__1881 (
            .O(N__10166),
            .I(N__10163));
    Odrv4 I__1880 (
            .O(N__10163),
            .I(TXbufferZ0Z_0));
    InMux I__1879 (
            .O(N__10160),
            .I(N__10157));
    LocalMux I__1878 (
            .O(N__10157),
            .I(\FTDI.TXshiftZ0Z_4 ));
    InMux I__1877 (
            .O(N__10154),
            .I(N__10151));
    LocalMux I__1876 (
            .O(N__10151),
            .I(TXbufferZ0Z_3));
    InMux I__1875 (
            .O(N__10148),
            .I(N__10145));
    LocalMux I__1874 (
            .O(N__10145),
            .I(\FTDI.TXshiftZ0Z_3 ));
    CascadeMux I__1873 (
            .O(N__10142),
            .I(N__10139));
    InMux I__1872 (
            .O(N__10139),
            .I(N__10136));
    LocalMux I__1871 (
            .O(N__10136),
            .I(N__10133));
    Odrv4 I__1870 (
            .O(N__10133),
            .I(\ALU.regsA_result_axb_6_l_ofx_1 ));
    CascadeMux I__1869 (
            .O(N__10130),
            .I(N__10127));
    InMux I__1868 (
            .O(N__10127),
            .I(N__10124));
    LocalMux I__1867 (
            .O(N__10124),
            .I(\ALU.mult_AdderTree2_bigtree_604 ));
    InMux I__1866 (
            .O(N__10121),
            .I(\ALU.regsA_result_cry_5_8 ));
    CascadeMux I__1865 (
            .O(N__10118),
            .I(N__10115));
    InMux I__1864 (
            .O(N__10115),
            .I(N__10112));
    LocalMux I__1863 (
            .O(N__10112),
            .I(\ALU.regsA_result_axb_7_l_ofx_1 ));
    CascadeMux I__1862 (
            .O(N__10109),
            .I(N__10106));
    InMux I__1861 (
            .O(N__10106),
            .I(N__10103));
    LocalMux I__1860 (
            .O(N__10103),
            .I(\ALU.mult_AdderTree2_bigtree_605 ));
    InMux I__1859 (
            .O(N__10100),
            .I(\ALU.regsA_result_cry_6_7 ));
    InMux I__1858 (
            .O(N__10097),
            .I(N__10094));
    LocalMux I__1857 (
            .O(N__10094),
            .I(N__10091));
    Odrv4 I__1856 (
            .O(N__10091),
            .I(\ALU.regsA_result_axb_8_l_ofx_0 ));
    CascadeMux I__1855 (
            .O(N__10088),
            .I(N__10085));
    InMux I__1854 (
            .O(N__10085),
            .I(N__10082));
    LocalMux I__1853 (
            .O(N__10082),
            .I(N__10079));
    Odrv4 I__1852 (
            .O(N__10079),
            .I(\ALU.regsA_result_cry_8_ma_0 ));
    CascadeMux I__1851 (
            .O(N__10076),
            .I(N__10073));
    InMux I__1850 (
            .O(N__10073),
            .I(N__10070));
    LocalMux I__1849 (
            .O(N__10070),
            .I(\ALU.mult_AdderTree2_bigtree_606 ));
    InMux I__1848 (
            .O(N__10067),
            .I(\ALU.regsA_result_cry_7_6 ));
    CascadeMux I__1847 (
            .O(N__10064),
            .I(N__10061));
    InMux I__1846 (
            .O(N__10061),
            .I(N__10058));
    LocalMux I__1845 (
            .O(N__10058),
            .I(\ALU.mult_AdderTree2_bigtree_607 ));
    InMux I__1844 (
            .O(N__10055),
            .I(bfn_14_16_0_));
    InMux I__1843 (
            .O(N__10052),
            .I(N__10049));
    LocalMux I__1842 (
            .O(N__10049),
            .I(\ALU.mult_AdderTree2_bigtree_608 ));
    InMux I__1841 (
            .O(N__10046),
            .I(\ALU.regsA_result_cry_9_4 ));
    InMux I__1840 (
            .O(N__10043),
            .I(N__10040));
    LocalMux I__1839 (
            .O(N__10040),
            .I(\ALU.mult_AdderTree2_bigtree_609 ));
    InMux I__1838 (
            .O(N__10037),
            .I(\ALU.regsA_result_cry_10_3 ));
    CascadeMux I__1837 (
            .O(N__10034),
            .I(N__10031));
    InMux I__1836 (
            .O(N__10031),
            .I(N__10028));
    LocalMux I__1835 (
            .O(N__10028),
            .I(N__10025));
    Span4Mux_v I__1834 (
            .O(N__10025),
            .I(N__10022));
    Odrv4 I__1833 (
            .O(N__10022),
            .I(\ALU.regsA_result_axb_12_1 ));
    InMux I__1832 (
            .O(N__10019),
            .I(\ALU.regsA_result_cry_11_1 ));
    CascadeMux I__1831 (
            .O(N__10016),
            .I(N__10013));
    InMux I__1830 (
            .O(N__10013),
            .I(N__10010));
    LocalMux I__1829 (
            .O(N__10010),
            .I(N__10007));
    Span4Mux_v I__1828 (
            .O(N__10007),
            .I(N__10004));
    Odrv4 I__1827 (
            .O(N__10004),
            .I(\ALU.regsA_result_axb_12 ));
    CascadeMux I__1826 (
            .O(N__10001),
            .I(N__9998));
    InMux I__1825 (
            .O(N__9998),
            .I(N__9995));
    LocalMux I__1824 (
            .O(N__9995),
            .I(\ALU.regsA_result_axb_10_l_ofx_0 ));
    InMux I__1823 (
            .O(N__9992),
            .I(N__9989));
    LocalMux I__1822 (
            .O(N__9989),
            .I(N__9986));
    Odrv4 I__1821 (
            .O(N__9986),
            .I(\ALU.regsA_result_cry_8_ma_1 ));
    InMux I__1820 (
            .O(N__9983),
            .I(\ALU.regsA_result_cry_1_7 ));
    CascadeMux I__1819 (
            .O(N__9980),
            .I(N__9977));
    InMux I__1818 (
            .O(N__9977),
            .I(N__9974));
    LocalMux I__1817 (
            .O(N__9974),
            .I(\ALU.mult_AdderTree2_bigtree_601 ));
    InMux I__1816 (
            .O(N__9971),
            .I(\ALU.regsA_result_cry_2_9 ));
    CascadeMux I__1815 (
            .O(N__9968),
            .I(N__9965));
    InMux I__1814 (
            .O(N__9965),
            .I(N__9962));
    LocalMux I__1813 (
            .O(N__9962),
            .I(\ALU.mult_AdderTree2_bigtree_602 ));
    InMux I__1812 (
            .O(N__9959),
            .I(\ALU.regsA_result_cry_3_9 ));
    CascadeMux I__1811 (
            .O(N__9956),
            .I(N__9953));
    InMux I__1810 (
            .O(N__9953),
            .I(N__9950));
    LocalMux I__1809 (
            .O(N__9950),
            .I(\ALU.mult_AdderTree2_bigtree_603 ));
    InMux I__1808 (
            .O(N__9947),
            .I(\ALU.regsA_result_cry_4_8 ));
    CascadeMux I__1807 (
            .O(N__9944),
            .I(N__9941));
    InMux I__1806 (
            .O(N__9941),
            .I(N__9938));
    LocalMux I__1805 (
            .O(N__9938),
            .I(N__9935));
    Span4Mux_v I__1804 (
            .O(N__9935),
            .I(N__9932));
    Odrv4 I__1803 (
            .O(N__9932),
            .I(\ALU.regsA_result_axb_6_l_ofx ));
    CascadeMux I__1802 (
            .O(N__9929),
            .I(N__9926));
    InMux I__1801 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__1800 (
            .O(N__9923),
            .I(N__9920));
    Span4Mux_h I__1799 (
            .O(N__9920),
            .I(N__9917));
    Odrv4 I__1798 (
            .O(N__9917),
            .I(\ALU.regsA_result_cry_5_ma ));
    InMux I__1797 (
            .O(N__9914),
            .I(N__9911));
    LocalMux I__1796 (
            .O(N__9911),
            .I(N__9908));
    Span4Mux_h I__1795 (
            .O(N__9908),
            .I(N__9905));
    Odrv4 I__1794 (
            .O(N__9905),
            .I(\ALU.regsA_result_axb_6_l_ofx_2 ));
    CascadeMux I__1793 (
            .O(N__9902),
            .I(N__9899));
    InMux I__1792 (
            .O(N__9899),
            .I(N__9896));
    LocalMux I__1791 (
            .O(N__9896),
            .I(N__9893));
    Odrv4 I__1790 (
            .O(N__9893),
            .I(\ALU.regsA_result_cry_7_ma_2 ));
    InMux I__1789 (
            .O(N__9890),
            .I(N__9887));
    LocalMux I__1788 (
            .O(N__9887),
            .I(N__9884));
    Span4Mux_h I__1787 (
            .O(N__9884),
            .I(N__9881));
    Odrv4 I__1786 (
            .O(N__9881),
            .I(\ALU.regsA_result_axb_7_l_ofx_2 ));
    InMux I__1785 (
            .O(N__9878),
            .I(N__9875));
    LocalMux I__1784 (
            .O(N__9875),
            .I(N__9872));
    Span4Mux_v I__1783 (
            .O(N__9872),
            .I(N__9869));
    Odrv4 I__1782 (
            .O(N__9869),
            .I(\ALU.regsA_result_cry_6_ma ));
    InMux I__1781 (
            .O(N__9866),
            .I(N__9863));
    LocalMux I__1780 (
            .O(N__9863),
            .I(\ALU.regsA_result_cry_2_ma_4 ));
    InMux I__1779 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1778 (
            .O(N__9857),
            .I(\ALU.regsA_result_cry_3_ma_4 ));
    CascadeMux I__1777 (
            .O(N__9854),
            .I(N__9851));
    InMux I__1776 (
            .O(N__9851),
            .I(N__9848));
    LocalMux I__1775 (
            .O(N__9848),
            .I(\ALU.regsA_result_cry_4_ma_3 ));
    CascadeMux I__1774 (
            .O(N__9845),
            .I(N__9842));
    InMux I__1773 (
            .O(N__9842),
            .I(N__9839));
    LocalMux I__1772 (
            .O(N__9839),
            .I(N__9836));
    Span4Mux_v I__1771 (
            .O(N__9836),
            .I(N__9833));
    Odrv4 I__1770 (
            .O(N__9833),
            .I(\ALU.mult_AdderTree2_bigtree_831 ));
    InMux I__1769 (
            .O(N__9830),
            .I(N__9825));
    InMux I__1768 (
            .O(N__9829),
            .I(N__9822));
    CascadeMux I__1767 (
            .O(N__9828),
            .I(N__9819));
    LocalMux I__1766 (
            .O(N__9825),
            .I(N__9816));
    LocalMux I__1765 (
            .O(N__9822),
            .I(N__9813));
    InMux I__1764 (
            .O(N__9819),
            .I(N__9810));
    Odrv4 I__1763 (
            .O(N__9816),
            .I(\ALU.mult_AdderTree2_bigtree_530 ));
    Odrv4 I__1762 (
            .O(N__9813),
            .I(\ALU.mult_AdderTree2_bigtree_530 ));
    LocalMux I__1761 (
            .O(N__9810),
            .I(\ALU.mult_AdderTree2_bigtree_530 ));
    InMux I__1760 (
            .O(N__9803),
            .I(N__9798));
    InMux I__1759 (
            .O(N__9802),
            .I(N__9795));
    InMux I__1758 (
            .O(N__9801),
            .I(N__9792));
    LocalMux I__1757 (
            .O(N__9798),
            .I(N__9786));
    LocalMux I__1756 (
            .O(N__9795),
            .I(N__9783));
    LocalMux I__1755 (
            .O(N__9792),
            .I(N__9780));
    InMux I__1754 (
            .O(N__9791),
            .I(N__9777));
    CascadeMux I__1753 (
            .O(N__9790),
            .I(N__9774));
    CascadeMux I__1752 (
            .O(N__9789),
            .I(N__9770));
    Span4Mux_v I__1751 (
            .O(N__9786),
            .I(N__9764));
    Span4Mux_v I__1750 (
            .O(N__9783),
            .I(N__9764));
    Span4Mux_h I__1749 (
            .O(N__9780),
            .I(N__9759));
    LocalMux I__1748 (
            .O(N__9777),
            .I(N__9759));
    InMux I__1747 (
            .O(N__9774),
            .I(N__9750));
    InMux I__1746 (
            .O(N__9773),
            .I(N__9750));
    InMux I__1745 (
            .O(N__9770),
            .I(N__9750));
    InMux I__1744 (
            .O(N__9769),
            .I(N__9750));
    Odrv4 I__1743 (
            .O(N__9764),
            .I(a_2_repZ0Z1));
    Odrv4 I__1742 (
            .O(N__9759),
            .I(a_2_repZ0Z1));
    LocalMux I__1741 (
            .O(N__9750),
            .I(a_2_repZ0Z1));
    InMux I__1740 (
            .O(N__9743),
            .I(N__9740));
    LocalMux I__1739 (
            .O(N__9740),
            .I(\ALU.regsA_result_cry_0_c_RNO_0 ));
    InMux I__1738 (
            .O(N__9737),
            .I(N__9734));
    LocalMux I__1737 (
            .O(N__9734),
            .I(N__9731));
    Odrv12 I__1736 (
            .O(N__9731),
            .I(\ALU.regsA_result_cry_4_ma ));
    CascadeMux I__1735 (
            .O(N__9728),
            .I(N__9725));
    InMux I__1734 (
            .O(N__9725),
            .I(N__9722));
    LocalMux I__1733 (
            .O(N__9722),
            .I(N__9719));
    Span4Mux_h I__1732 (
            .O(N__9719),
            .I(N__9716));
    Odrv4 I__1731 (
            .O(N__9716),
            .I(\ALU.regsA_result_cry_6_ma_2 ));
    CascadeMux I__1730 (
            .O(N__9713),
            .I(N__9710));
    InMux I__1729 (
            .O(N__9710),
            .I(N__9707));
    LocalMux I__1728 (
            .O(N__9707),
            .I(\ALU.regsA_result_axb_2_l_ofx_4 ));
    CascadeMux I__1727 (
            .O(N__9704),
            .I(N__9701));
    InMux I__1726 (
            .O(N__9701),
            .I(N__9698));
    LocalMux I__1725 (
            .O(N__9698),
            .I(\ALU.regsA_result_axb_3_l_ofx_4 ));
    InMux I__1724 (
            .O(N__9695),
            .I(N__9692));
    LocalMux I__1723 (
            .O(N__9692),
            .I(\ALU.regsA_result_axb_4_l_ofx_3 ));
    CascadeMux I__1722 (
            .O(N__9689),
            .I(N__9686));
    InMux I__1721 (
            .O(N__9686),
            .I(N__9683));
    LocalMux I__1720 (
            .O(N__9683),
            .I(\ALU.regsA_result_axb_5_l_ofx_3 ));
    InMux I__1719 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__1718 (
            .O(N__9677),
            .I(N__9674));
    Odrv4 I__1717 (
            .O(N__9674),
            .I(\ALU.mult_AdderTree2_bigtree_564 ));
    CascadeMux I__1716 (
            .O(N__9671),
            .I(N__9668));
    InMux I__1715 (
            .O(N__9668),
            .I(N__9664));
    InMux I__1714 (
            .O(N__9667),
            .I(N__9661));
    LocalMux I__1713 (
            .O(N__9664),
            .I(a_fastZ0Z_2));
    LocalMux I__1712 (
            .O(N__9661),
            .I(a_fastZ0Z_2));
    CascadeMux I__1711 (
            .O(N__9656),
            .I(N__9653));
    InMux I__1710 (
            .O(N__9653),
            .I(N__9650));
    LocalMux I__1709 (
            .O(N__9650),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_4 ));
    InMux I__1708 (
            .O(N__9647),
            .I(N__9644));
    LocalMux I__1707 (
            .O(N__9644),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_5 ));
    CascadeMux I__1706 (
            .O(N__9641),
            .I(N__9638));
    InMux I__1705 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__1704 (
            .O(N__9635),
            .I(N__9632));
    Span4Mux_v I__1703 (
            .O(N__9632),
            .I(N__9629));
    Odrv4 I__1702 (
            .O(N__9629),
            .I(\ALU.regsA_result_axb_11_l_ofx ));
    InMux I__1701 (
            .O(N__9626),
            .I(N__9623));
    LocalMux I__1700 (
            .O(N__9623),
            .I(N__9620));
    Span4Mux_h I__1699 (
            .O(N__9620),
            .I(N__9617));
    Span4Mux_v I__1698 (
            .O(N__9617),
            .I(N__9614));
    Odrv4 I__1697 (
            .O(N__9614),
            .I(\ALU.regsA_result_cry_10_ma ));
    CascadeMux I__1696 (
            .O(N__9611),
            .I(N__9608));
    InMux I__1695 (
            .O(N__9608),
            .I(N__9605));
    LocalMux I__1694 (
            .O(N__9605),
            .I(N__9602));
    Odrv4 I__1693 (
            .O(N__9602),
            .I(\ALU.regsA_result_axb_11_l_ofx_1 ));
    InMux I__1692 (
            .O(N__9599),
            .I(N__9596));
    LocalMux I__1691 (
            .O(N__9596),
            .I(N__9590));
    CascadeMux I__1690 (
            .O(N__9595),
            .I(N__9587));
    CascadeMux I__1689 (
            .O(N__9594),
            .I(N__9584));
    CascadeMux I__1688 (
            .O(N__9593),
            .I(N__9578));
    Span4Mux_h I__1687 (
            .O(N__9590),
            .I(N__9574));
    InMux I__1686 (
            .O(N__9587),
            .I(N__9565));
    InMux I__1685 (
            .O(N__9584),
            .I(N__9565));
    InMux I__1684 (
            .O(N__9583),
            .I(N__9565));
    InMux I__1683 (
            .O(N__9582),
            .I(N__9565));
    InMux I__1682 (
            .O(N__9581),
            .I(N__9558));
    InMux I__1681 (
            .O(N__9578),
            .I(N__9558));
    InMux I__1680 (
            .O(N__9577),
            .I(N__9558));
    Odrv4 I__1679 (
            .O(N__9574),
            .I(bZ0Z_12));
    LocalMux I__1678 (
            .O(N__9565),
            .I(bZ0Z_12));
    LocalMux I__1677 (
            .O(N__9558),
            .I(bZ0Z_12));
    CascadeMux I__1676 (
            .O(N__9551),
            .I(N__9548));
    InMux I__1675 (
            .O(N__9548),
            .I(N__9545));
    LocalMux I__1674 (
            .O(N__9545),
            .I(N__9542));
    Span4Mux_v I__1673 (
            .O(N__9542),
            .I(N__9539));
    Odrv4 I__1672 (
            .O(N__9539),
            .I(\ALU.regsA_result_axb_12_l_ofx_0 ));
    InMux I__1671 (
            .O(N__9536),
            .I(N__9533));
    LocalMux I__1670 (
            .O(N__9533),
            .I(N__9530));
    Odrv4 I__1669 (
            .O(N__9530),
            .I(\ALU.regsA_result_axb_10_l_ofx_1 ));
    InMux I__1668 (
            .O(N__9527),
            .I(N__9524));
    LocalMux I__1667 (
            .O(N__9524),
            .I(N__9521));
    Span4Mux_v I__1666 (
            .O(N__9521),
            .I(N__9518));
    Odrv4 I__1665 (
            .O(N__9518),
            .I(\ALU.regsA_result_cry_11_ma_1 ));
    InMux I__1664 (
            .O(N__9515),
            .I(N__9512));
    LocalMux I__1663 (
            .O(N__9512),
            .I(\ALU.mult_AdderTree2_bigtree_840 ));
    InMux I__1662 (
            .O(N__9509),
            .I(\ALU.regsA_result_cry_10_1 ));
    InMux I__1661 (
            .O(N__9506),
            .I(\ALU.regsA_result_cry_11 ));
    InMux I__1660 (
            .O(N__9503),
            .I(N__9500));
    LocalMux I__1659 (
            .O(N__9500),
            .I(N__9497));
    Odrv4 I__1658 (
            .O(N__9497),
            .I(\ALU.regsA_result_cry_11_THRU_CO ));
    CascadeMux I__1657 (
            .O(N__9494),
            .I(N__9491));
    InMux I__1656 (
            .O(N__9491),
            .I(N__9488));
    LocalMux I__1655 (
            .O(N__9488),
            .I(N__9485));
    Odrv4 I__1654 (
            .O(N__9485),
            .I(\ALU.regsA_result_axb_10_l_ofx ));
    InMux I__1653 (
            .O(N__9482),
            .I(N__9479));
    LocalMux I__1652 (
            .O(N__9479),
            .I(N__9476));
    Span4Mux_v I__1651 (
            .O(N__9476),
            .I(N__9473));
    Odrv4 I__1650 (
            .O(N__9473),
            .I(\ALU.addsub_3 ));
    InMux I__1649 (
            .O(N__9470),
            .I(N__9467));
    LocalMux I__1648 (
            .O(N__9467),
            .I(N__9464));
    Odrv12 I__1647 (
            .O(N__9464),
            .I(\ALU.mult_3 ));
    CascadeMux I__1646 (
            .O(N__9461),
            .I(N__9458));
    InMux I__1645 (
            .O(N__9458),
            .I(N__9455));
    LocalMux I__1644 (
            .O(N__9455),
            .I(N__9452));
    Span4Mux_v I__1643 (
            .O(N__9452),
            .I(N__9449));
    Odrv4 I__1642 (
            .O(N__9449),
            .I(res_11));
    InMux I__1641 (
            .O(N__9446),
            .I(N__9443));
    LocalMux I__1640 (
            .O(N__9443),
            .I(res_3));
    IoInMux I__1639 (
            .O(N__9440),
            .I(N__9437));
    LocalMux I__1638 (
            .O(N__9437),
            .I(N__9434));
    IoSpan4Mux I__1637 (
            .O(N__9434),
            .I(N__9431));
    Span4Mux_s3_h I__1636 (
            .O(N__9431),
            .I(N__9428));
    Sp12to4 I__1635 (
            .O(N__9428),
            .I(N__9424));
    InMux I__1634 (
            .O(N__9427),
            .I(N__9421));
    Span12Mux_s10_h I__1633 (
            .O(N__9424),
            .I(N__9418));
    LocalMux I__1632 (
            .O(N__9421),
            .I(N__9415));
    Odrv12 I__1631 (
            .O(N__9418),
            .I(GPIO1_c));
    Odrv4 I__1630 (
            .O(N__9415),
            .I(GPIO1_c));
    CascadeMux I__1629 (
            .O(N__9410),
            .I(N__9407));
    InMux I__1628 (
            .O(N__9407),
            .I(N__9404));
    LocalMux I__1627 (
            .O(N__9404),
            .I(N__9401));
    Odrv4 I__1626 (
            .O(N__9401),
            .I(res_9));
    CascadeMux I__1625 (
            .O(N__9398),
            .I(N__9395));
    InMux I__1624 (
            .O(N__9395),
            .I(N__9392));
    LocalMux I__1623 (
            .O(N__9392),
            .I(N__9389));
    Odrv4 I__1622 (
            .O(N__9389),
            .I(res_12));
    CEMux I__1621 (
            .O(N__9386),
            .I(N__9382));
    CEMux I__1620 (
            .O(N__9385),
            .I(N__9379));
    LocalMux I__1619 (
            .O(N__9382),
            .I(TXstate_fast_RNIP6NA1_3));
    LocalMux I__1618 (
            .O(N__9379),
            .I(TXstate_fast_RNIP6NA1_3));
    CascadeMux I__1617 (
            .O(N__9374),
            .I(N__9371));
    InMux I__1616 (
            .O(N__9371),
            .I(N__9368));
    LocalMux I__1615 (
            .O(N__9368),
            .I(\ALU.mult_AdderTree2_bigtree_832 ));
    InMux I__1614 (
            .O(N__9365),
            .I(\ALU.regsA_result_cry_2_4 ));
    CascadeMux I__1613 (
            .O(N__9362),
            .I(N__9359));
    InMux I__1612 (
            .O(N__9359),
            .I(N__9356));
    LocalMux I__1611 (
            .O(N__9356),
            .I(\ALU.mult_AdderTree2_bigtree_833 ));
    InMux I__1610 (
            .O(N__9353),
            .I(\ALU.regsA_result_cry_3_5 ));
    CascadeMux I__1609 (
            .O(N__9350),
            .I(N__9347));
    InMux I__1608 (
            .O(N__9347),
            .I(N__9344));
    LocalMux I__1607 (
            .O(N__9344),
            .I(\ALU.mult_AdderTree2_bigtree_834 ));
    InMux I__1606 (
            .O(N__9341),
            .I(\ALU.regsA_result_cry_4_4 ));
    CascadeMux I__1605 (
            .O(N__9338),
            .I(N__9335));
    InMux I__1604 (
            .O(N__9335),
            .I(N__9332));
    LocalMux I__1603 (
            .O(N__9332),
            .I(\ALU.mult_AdderTree2_bigtree_835 ));
    InMux I__1602 (
            .O(N__9329),
            .I(\ALU.regsA_result_cry_5_5 ));
    CascadeMux I__1601 (
            .O(N__9326),
            .I(N__9323));
    InMux I__1600 (
            .O(N__9323),
            .I(N__9320));
    LocalMux I__1599 (
            .O(N__9320),
            .I(\ALU.mult_AdderTree2_bigtree_836 ));
    InMux I__1598 (
            .O(N__9317),
            .I(\ALU.regsA_result_cry_6_4 ));
    CascadeMux I__1597 (
            .O(N__9314),
            .I(N__9311));
    InMux I__1596 (
            .O(N__9311),
            .I(N__9308));
    LocalMux I__1595 (
            .O(N__9308),
            .I(\ALU.mult_AdderTree2_bigtree_837 ));
    InMux I__1594 (
            .O(N__9305),
            .I(\ALU.regsA_result_cry_7_4 ));
    CascadeMux I__1593 (
            .O(N__9302),
            .I(N__9299));
    InMux I__1592 (
            .O(N__9299),
            .I(N__9296));
    LocalMux I__1591 (
            .O(N__9296),
            .I(\ALU.mult_AdderTree2_bigtree_838 ));
    InMux I__1590 (
            .O(N__9293),
            .I(\ALU.regsA_result_cry_8_1 ));
    CascadeMux I__1589 (
            .O(N__9290),
            .I(N__9287));
    InMux I__1588 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__1587 (
            .O(N__9284),
            .I(\ALU.mult_AdderTree2_bigtree_839 ));
    InMux I__1586 (
            .O(N__9281),
            .I(bfn_13_16_0_));
    InMux I__1585 (
            .O(N__9278),
            .I(N__9275));
    LocalMux I__1584 (
            .O(N__9275),
            .I(\ALU.mult_AdderTree2_bigtree_538 ));
    CascadeMux I__1583 (
            .O(N__9272),
            .I(N__9269));
    InMux I__1582 (
            .O(N__9269),
            .I(N__9266));
    LocalMux I__1581 (
            .O(N__9266),
            .I(N__9263));
    Odrv4 I__1580 (
            .O(N__9263),
            .I(\ALU.mult_AdderTree2_bigtree_571 ));
    InMux I__1579 (
            .O(N__9260),
            .I(N__9257));
    LocalMux I__1578 (
            .O(N__9257),
            .I(\ALU.mult_AdderTree2_bigtree_802 ));
    InMux I__1577 (
            .O(N__9254),
            .I(bfn_13_14_0_));
    InMux I__1576 (
            .O(N__9251),
            .I(N__9248));
    LocalMux I__1575 (
            .O(N__9248),
            .I(\ALU.mult_AdderTree2_bigtree_539 ));
    CascadeMux I__1574 (
            .O(N__9245),
            .I(N__9242));
    InMux I__1573 (
            .O(N__9242),
            .I(N__9239));
    LocalMux I__1572 (
            .O(N__9239),
            .I(N__9236));
    Odrv4 I__1571 (
            .O(N__9236),
            .I(\ALU.mult_AdderTree2_bigtree_572 ));
    InMux I__1570 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__1569 (
            .O(N__9230),
            .I(\ALU.mult_AdderTree2_bigtree_803 ));
    InMux I__1568 (
            .O(N__9227),
            .I(\ALU.regsA_result_cry_8_0 ));
    InMux I__1567 (
            .O(N__9224),
            .I(N__9221));
    LocalMux I__1566 (
            .O(N__9221),
            .I(\ALU.mult_AdderTree2_bigtree_540 ));
    CascadeMux I__1565 (
            .O(N__9218),
            .I(N__9215));
    InMux I__1564 (
            .O(N__9215),
            .I(N__9212));
    LocalMux I__1563 (
            .O(N__9212),
            .I(N__9209));
    Odrv4 I__1562 (
            .O(N__9209),
            .I(\ALU.mult_AdderTree2_bigtree_573 ));
    InMux I__1561 (
            .O(N__9206),
            .I(N__9203));
    LocalMux I__1560 (
            .O(N__9203),
            .I(N__9200));
    Span4Mux_v I__1559 (
            .O(N__9200),
            .I(N__9197));
    Odrv4 I__1558 (
            .O(N__9197),
            .I(\ALU.mult_AdderTree2_bigtree_804 ));
    InMux I__1557 (
            .O(N__9194),
            .I(\ALU.regsA_result_cry_9_1 ));
    InMux I__1556 (
            .O(N__9191),
            .I(N__9188));
    LocalMux I__1555 (
            .O(N__9188),
            .I(\ALU.mult_AdderTree2_bigtree_541 ));
    CascadeMux I__1554 (
            .O(N__9185),
            .I(N__9182));
    InMux I__1553 (
            .O(N__9182),
            .I(N__9179));
    LocalMux I__1552 (
            .O(N__9179),
            .I(N__9176));
    Odrv4 I__1551 (
            .O(N__9176),
            .I(\ALU.mult_AdderTree2_bigtree_574 ));
    InMux I__1550 (
            .O(N__9173),
            .I(N__9170));
    LocalMux I__1549 (
            .O(N__9170),
            .I(N__9167));
    Odrv4 I__1548 (
            .O(N__9167),
            .I(\ALU.mult_AdderTree2_bigtree_805 ));
    InMux I__1547 (
            .O(N__9164),
            .I(\ALU.regsA_result_cry_10_0 ));
    InMux I__1546 (
            .O(N__9161),
            .I(N__9158));
    LocalMux I__1545 (
            .O(N__9158),
            .I(\ALU.mult_AdderTree2_bigtree_542 ));
    CascadeMux I__1544 (
            .O(N__9155),
            .I(N__9152));
    InMux I__1543 (
            .O(N__9152),
            .I(N__9149));
    LocalMux I__1542 (
            .O(N__9149),
            .I(N__9146));
    Odrv4 I__1541 (
            .O(N__9146),
            .I(\ALU.mult_AdderTree2_bigtree_575 ));
    InMux I__1540 (
            .O(N__9143),
            .I(N__9140));
    LocalMux I__1539 (
            .O(N__9140),
            .I(N__9137));
    Odrv4 I__1538 (
            .O(N__9137),
            .I(\ALU.mult_AdderTree2_bigtree_806 ));
    InMux I__1537 (
            .O(N__9134),
            .I(\ALU.regsA_result_cry_11_2 ));
    InMux I__1536 (
            .O(N__9131),
            .I(N__9128));
    LocalMux I__1535 (
            .O(N__9128),
            .I(\ALU.mult_AdderTree2_bigtree_543 ));
    CascadeMux I__1534 (
            .O(N__9125),
            .I(N__9122));
    InMux I__1533 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__1532 (
            .O(N__9119),
            .I(N__9116));
    Span4Mux_h I__1531 (
            .O(N__9116),
            .I(N__9113));
    Odrv4 I__1530 (
            .O(N__9113),
            .I(\ALU.mult_AdderTree2_bigtree_576 ));
    CascadeMux I__1529 (
            .O(N__9110),
            .I(N__9107));
    InMux I__1528 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__1527 (
            .O(N__9104),
            .I(N__9101));
    Odrv4 I__1526 (
            .O(N__9101),
            .I(\ALU.mult_AdderTree2_bigtree_807 ));
    InMux I__1525 (
            .O(N__9098),
            .I(\ALU.regsA_result_cry_12 ));
    InMux I__1524 (
            .O(N__9095),
            .I(N__9092));
    LocalMux I__1523 (
            .O(N__9092),
            .I(\ALU.regsA_result_axb_14 ));
    InMux I__1522 (
            .O(N__9089),
            .I(\ALU.regsA_result_cry_13 ));
    InMux I__1521 (
            .O(N__9086),
            .I(N__9083));
    LocalMux I__1520 (
            .O(N__9083),
            .I(N__9080));
    Odrv4 I__1519 (
            .O(N__9080),
            .I(\ALU.regsA_result_axb_12_0 ));
    CascadeMux I__1518 (
            .O(N__9077),
            .I(N__9074));
    InMux I__1517 (
            .O(N__9074),
            .I(N__9071));
    LocalMux I__1516 (
            .O(N__9071),
            .I(\ALU.mult_AdderTree2_bigtree_531 ));
    InMux I__1515 (
            .O(N__9068),
            .I(\ALU.regsA_result_cry_0_1 ));
    InMux I__1514 (
            .O(N__9065),
            .I(N__9062));
    LocalMux I__1513 (
            .O(N__9062),
            .I(\ALU.mult_AdderTree2_bigtree_532 ));
    CascadeMux I__1512 (
            .O(N__9059),
            .I(N__9056));
    InMux I__1511 (
            .O(N__9056),
            .I(N__9053));
    LocalMux I__1510 (
            .O(N__9053),
            .I(N__9050));
    Odrv4 I__1509 (
            .O(N__9050),
            .I(\ALU.mult_AdderTree2_bigtree_565 ));
    InMux I__1508 (
            .O(N__9047),
            .I(\ALU.regsA_result_cry_1_2 ));
    InMux I__1507 (
            .O(N__9044),
            .I(N__9041));
    LocalMux I__1506 (
            .O(N__9041),
            .I(\ALU.mult_AdderTree2_bigtree_533 ));
    CascadeMux I__1505 (
            .O(N__9038),
            .I(N__9035));
    InMux I__1504 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__1503 (
            .O(N__9032),
            .I(N__9029));
    Odrv4 I__1502 (
            .O(N__9029),
            .I(\ALU.mult_AdderTree2_bigtree_566 ));
    InMux I__1501 (
            .O(N__9026),
            .I(N__9023));
    LocalMux I__1500 (
            .O(N__9023),
            .I(N__9020));
    Odrv4 I__1499 (
            .O(N__9020),
            .I(\ALU.mult_AdderTree2_bigtree_797 ));
    InMux I__1498 (
            .O(N__9017),
            .I(\ALU.regsA_result_cry_2_3 ));
    InMux I__1497 (
            .O(N__9014),
            .I(N__9011));
    LocalMux I__1496 (
            .O(N__9011),
            .I(\ALU.mult_AdderTree2_bigtree_534 ));
    CascadeMux I__1495 (
            .O(N__9008),
            .I(N__9005));
    InMux I__1494 (
            .O(N__9005),
            .I(N__9002));
    LocalMux I__1493 (
            .O(N__9002),
            .I(N__8999));
    Odrv4 I__1492 (
            .O(N__8999),
            .I(\ALU.mult_AdderTree2_bigtree_567 ));
    InMux I__1491 (
            .O(N__8996),
            .I(N__8993));
    LocalMux I__1490 (
            .O(N__8993),
            .I(N__8990));
    Odrv4 I__1489 (
            .O(N__8990),
            .I(\ALU.mult_AdderTree2_bigtree_798 ));
    InMux I__1488 (
            .O(N__8987),
            .I(\ALU.regsA_result_cry_3_3 ));
    InMux I__1487 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__1486 (
            .O(N__8981),
            .I(\ALU.mult_AdderTree2_bigtree_535 ));
    CascadeMux I__1485 (
            .O(N__8978),
            .I(N__8975));
    InMux I__1484 (
            .O(N__8975),
            .I(N__8972));
    LocalMux I__1483 (
            .O(N__8972),
            .I(N__8969));
    Odrv4 I__1482 (
            .O(N__8969),
            .I(\ALU.mult_AdderTree2_bigtree_568 ));
    InMux I__1481 (
            .O(N__8966),
            .I(N__8963));
    LocalMux I__1480 (
            .O(N__8963),
            .I(N__8960));
    Span12Mux_v I__1479 (
            .O(N__8960),
            .I(N__8957));
    Odrv12 I__1478 (
            .O(N__8957),
            .I(\ALU.mult_AdderTree2_bigtree_799 ));
    InMux I__1477 (
            .O(N__8954),
            .I(\ALU.regsA_result_cry_4_2 ));
    InMux I__1476 (
            .O(N__8951),
            .I(N__8948));
    LocalMux I__1475 (
            .O(N__8948),
            .I(\ALU.mult_AdderTree2_bigtree_536 ));
    CascadeMux I__1474 (
            .O(N__8945),
            .I(N__8942));
    InMux I__1473 (
            .O(N__8942),
            .I(N__8939));
    LocalMux I__1472 (
            .O(N__8939),
            .I(N__8936));
    Odrv4 I__1471 (
            .O(N__8936),
            .I(\ALU.mult_AdderTree2_bigtree_569 ));
    InMux I__1470 (
            .O(N__8933),
            .I(N__8930));
    LocalMux I__1469 (
            .O(N__8930),
            .I(N__8927));
    Odrv4 I__1468 (
            .O(N__8927),
            .I(\ALU.mult_AdderTree2_bigtree_800 ));
    InMux I__1467 (
            .O(N__8924),
            .I(\ALU.regsA_result_cry_5_3 ));
    InMux I__1466 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__1465 (
            .O(N__8918),
            .I(\ALU.mult_AdderTree2_bigtree_537 ));
    CascadeMux I__1464 (
            .O(N__8915),
            .I(N__8912));
    InMux I__1463 (
            .O(N__8912),
            .I(N__8909));
    LocalMux I__1462 (
            .O(N__8909),
            .I(N__8906));
    Odrv12 I__1461 (
            .O(N__8906),
            .I(\ALU.mult_AdderTree2_bigtree_570 ));
    InMux I__1460 (
            .O(N__8903),
            .I(N__8900));
    LocalMux I__1459 (
            .O(N__8900),
            .I(N__8897));
    Span4Mux_h I__1458 (
            .O(N__8897),
            .I(N__8894));
    Odrv4 I__1457 (
            .O(N__8894),
            .I(\ALU.mult_AdderTree2_bigtree_801 ));
    InMux I__1456 (
            .O(N__8891),
            .I(\ALU.regsA_result_cry_6_2 ));
    InMux I__1455 (
            .O(N__8888),
            .I(\ALU.regsA_result_cry_7_7 ));
    InMux I__1454 (
            .O(N__8885),
            .I(bfn_13_12_0_));
    InMux I__1453 (
            .O(N__8882),
            .I(\ALU.regsA_result_cry_9_5 ));
    InMux I__1452 (
            .O(N__8879),
            .I(\ALU.regsA_result_cry_10_4 ));
    InMux I__1451 (
            .O(N__8876),
            .I(\ALU.regsA_result_cry_11_4 ));
    InMux I__1450 (
            .O(N__8873),
            .I(N__8870));
    LocalMux I__1449 (
            .O(N__8870),
            .I(N__8867));
    Odrv12 I__1448 (
            .O(N__8867),
            .I(\ALU.regsA_result_cry_13_ma_0 ));
    CascadeMux I__1447 (
            .O(N__8864),
            .I(N__8861));
    InMux I__1446 (
            .O(N__8861),
            .I(N__8858));
    LocalMux I__1445 (
            .O(N__8858),
            .I(N__8855));
    Odrv4 I__1444 (
            .O(N__8855),
            .I(\ALU.regsA_result_axb_13_l_ofx_0 ));
    InMux I__1443 (
            .O(N__8852),
            .I(\ALU.regsA_result_cry_12_1 ));
    InMux I__1442 (
            .O(N__8849),
            .I(\ALU.regsA_result_cry_13_0 ));
    CascadeMux I__1441 (
            .O(N__8846),
            .I(N__8843));
    InMux I__1440 (
            .O(N__8843),
            .I(N__8840));
    LocalMux I__1439 (
            .O(N__8840),
            .I(\ALU.regsA_result_cry_13_0_THRU_CO ));
    InMux I__1438 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__1437 (
            .O(N__8834),
            .I(\ALU.regsA_result_cry_12_ma_0 ));
    InMux I__1436 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__1435 (
            .O(N__8828),
            .I(\ALU.regsA_result_cry_0_0_c_RNO_0 ));
    InMux I__1434 (
            .O(N__8825),
            .I(N__8822));
    LocalMux I__1433 (
            .O(N__8822),
            .I(N__8819));
    Odrv4 I__1432 (
            .O(N__8819),
            .I(\ALU.regsA_result_cry_12_ma ));
    CascadeMux I__1431 (
            .O(N__8816),
            .I(N__8813));
    InMux I__1430 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__1429 (
            .O(N__8810),
            .I(N__8807));
    Odrv4 I__1428 (
            .O(N__8807),
            .I(\ALU.regsA_result_axb_13_l_ofx ));
    InMux I__1427 (
            .O(N__8804),
            .I(\ALU.regsA_result_cry_1_8 ));
    InMux I__1426 (
            .O(N__8801),
            .I(\ALU.regsA_result_cry_2_10 ));
    InMux I__1425 (
            .O(N__8798),
            .I(\ALU.regsA_result_cry_3_10 ));
    InMux I__1424 (
            .O(N__8795),
            .I(N__8792));
    LocalMux I__1423 (
            .O(N__8792),
            .I(N__8789));
    Odrv4 I__1422 (
            .O(N__8789),
            .I(\ALU.regsA_result_cry_5_ma_3 ));
    InMux I__1421 (
            .O(N__8786),
            .I(\ALU.regsA_result_cry_4_9 ));
    InMux I__1420 (
            .O(N__8783),
            .I(\ALU.regsA_result_cry_5_9 ));
    InMux I__1419 (
            .O(N__8780),
            .I(\ALU.regsA_result_cry_6_8 ));
    InMux I__1418 (
            .O(N__8777),
            .I(N__8774));
    LocalMux I__1417 (
            .O(N__8774),
            .I(N__8771));
    Odrv12 I__1416 (
            .O(N__8771),
            .I(res_6));
    InMux I__1415 (
            .O(N__8768),
            .I(N__8765));
    LocalMux I__1414 (
            .O(N__8765),
            .I(res_14));
    InMux I__1413 (
            .O(N__8762),
            .I(N__8759));
    LocalMux I__1412 (
            .O(N__8759),
            .I(N__8756));
    Odrv12 I__1411 (
            .O(N__8756),
            .I(res_15));
    InMux I__1410 (
            .O(N__8753),
            .I(N__8750));
    LocalMux I__1409 (
            .O(N__8750),
            .I(res_7));
    InMux I__1408 (
            .O(N__8747),
            .I(N__8740));
    InMux I__1407 (
            .O(N__8746),
            .I(N__8736));
    CascadeMux I__1406 (
            .O(N__8745),
            .I(N__8733));
    CascadeMux I__1405 (
            .O(N__8744),
            .I(N__8730));
    CascadeMux I__1404 (
            .O(N__8743),
            .I(N__8727));
    LocalMux I__1403 (
            .O(N__8740),
            .I(N__8724));
    InMux I__1402 (
            .O(N__8739),
            .I(N__8720));
    LocalMux I__1401 (
            .O(N__8736),
            .I(N__8716));
    InMux I__1400 (
            .O(N__8733),
            .I(N__8709));
    InMux I__1399 (
            .O(N__8730),
            .I(N__8709));
    InMux I__1398 (
            .O(N__8727),
            .I(N__8709));
    Span4Mux_v I__1397 (
            .O(N__8724),
            .I(N__8706));
    InMux I__1396 (
            .O(N__8723),
            .I(N__8703));
    LocalMux I__1395 (
            .O(N__8720),
            .I(N__8700));
    CascadeMux I__1394 (
            .O(N__8719),
            .I(N__8693));
    Span4Mux_h I__1393 (
            .O(N__8716),
            .I(N__8686));
    LocalMux I__1392 (
            .O(N__8709),
            .I(N__8686));
    Span4Mux_v I__1391 (
            .O(N__8706),
            .I(N__8683));
    LocalMux I__1390 (
            .O(N__8703),
            .I(N__8678));
    Span4Mux_h I__1389 (
            .O(N__8700),
            .I(N__8678));
    InMux I__1388 (
            .O(N__8699),
            .I(N__8675));
    InMux I__1387 (
            .O(N__8698),
            .I(N__8662));
    InMux I__1386 (
            .O(N__8697),
            .I(N__8662));
    InMux I__1385 (
            .O(N__8696),
            .I(N__8662));
    InMux I__1384 (
            .O(N__8693),
            .I(N__8662));
    InMux I__1383 (
            .O(N__8692),
            .I(N__8662));
    InMux I__1382 (
            .O(N__8691),
            .I(N__8662));
    Odrv4 I__1381 (
            .O(N__8686),
            .I(aZ0Z_11));
    Odrv4 I__1380 (
            .O(N__8683),
            .I(aZ0Z_11));
    Odrv4 I__1379 (
            .O(N__8678),
            .I(aZ0Z_11));
    LocalMux I__1378 (
            .O(N__8675),
            .I(aZ0Z_11));
    LocalMux I__1377 (
            .O(N__8662),
            .I(aZ0Z_11));
    CascadeMux I__1376 (
            .O(N__8651),
            .I(N__8648));
    InMux I__1375 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__1374 (
            .O(N__8645),
            .I(N__8642));
    Span4Mux_h I__1373 (
            .O(N__8642),
            .I(N__8639));
    Span4Mux_v I__1372 (
            .O(N__8639),
            .I(N__8636));
    Odrv4 I__1371 (
            .O(N__8636),
            .I(\ALU.addsub_axb_11_l_ofxZ0 ));
    CascadeMux I__1370 (
            .O(N__8633),
            .I(N__8630));
    InMux I__1369 (
            .O(N__8630),
            .I(N__8627));
    LocalMux I__1368 (
            .O(N__8627),
            .I(N__8624));
    Span4Mux_v I__1367 (
            .O(N__8624),
            .I(N__8621));
    Odrv4 I__1366 (
            .O(N__8621),
            .I(\ALU.regsA_result_axb_12_l_ofx ));
    InMux I__1365 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__1364 (
            .O(N__8615),
            .I(N__8612));
    Odrv4 I__1363 (
            .O(N__8612),
            .I(\ALU.regsA_result_cry_11_ma ));
    InMux I__1362 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__1361 (
            .O(N__8606),
            .I(N__8603));
    Span4Mux_h I__1360 (
            .O(N__8603),
            .I(N__8599));
    InMux I__1359 (
            .O(N__8602),
            .I(N__8596));
    Span4Mux_v I__1358 (
            .O(N__8599),
            .I(N__8591));
    LocalMux I__1357 (
            .O(N__8596),
            .I(N__8591));
    Odrv4 I__1356 (
            .O(N__8591),
            .I(\ALU.mult_AdderTree2_bigtree_938 ));
    InMux I__1355 (
            .O(N__8588),
            .I(\ALU.regsA_result_cry_9_0 ));
    InMux I__1354 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__1353 (
            .O(N__8582),
            .I(N__8578));
    InMux I__1352 (
            .O(N__8581),
            .I(N__8575));
    Span4Mux_h I__1351 (
            .O(N__8578),
            .I(N__8572));
    LocalMux I__1350 (
            .O(N__8575),
            .I(N__8569));
    Span4Mux_v I__1349 (
            .O(N__8572),
            .I(N__8564));
    Span4Mux_h I__1348 (
            .O(N__8569),
            .I(N__8564));
    Odrv4 I__1347 (
            .O(N__8564),
            .I(\ALU.mult_AdderTree2_bigtree_939 ));
    InMux I__1346 (
            .O(N__8561),
            .I(\ALU.regsA_result_cry_10 ));
    InMux I__1345 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__1344 (
            .O(N__8555),
            .I(N__8552));
    Span4Mux_h I__1343 (
            .O(N__8552),
            .I(N__8549));
    Span4Mux_v I__1342 (
            .O(N__8549),
            .I(N__8546));
    Odrv4 I__1341 (
            .O(N__8546),
            .I(\ALU.regsA_result_axb_8 ));
    CascadeMux I__1340 (
            .O(N__8543),
            .I(N__8540));
    InMux I__1339 (
            .O(N__8540),
            .I(N__8537));
    LocalMux I__1338 (
            .O(N__8537),
            .I(N__8534));
    Span4Mux_v I__1337 (
            .O(N__8534),
            .I(N__8531));
    Odrv4 I__1336 (
            .O(N__8531),
            .I(\ALU.regsA_result_cry_7_THRU_CO ));
    InMux I__1335 (
            .O(N__8528),
            .I(\ALU.regsA_result_cry_11_0 ));
    InMux I__1334 (
            .O(N__8525),
            .I(N__8522));
    LocalMux I__1333 (
            .O(N__8522),
            .I(N__8519));
    Span4Mux_v I__1332 (
            .O(N__8519),
            .I(N__8516));
    Odrv4 I__1331 (
            .O(N__8516),
            .I(\ALU.regsA_result_axb_8_0 ));
    InMux I__1330 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__1329 (
            .O(N__8510),
            .I(\ALU.mult_5 ));
    InMux I__1328 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__1327 (
            .O(N__8504),
            .I(N__8501));
    Odrv4 I__1326 (
            .O(N__8501),
            .I(\ALU.addsub_5 ));
    InMux I__1325 (
            .O(N__8498),
            .I(N__8495));
    LocalMux I__1324 (
            .O(N__8495),
            .I(N__8492));
    Odrv4 I__1323 (
            .O(N__8492),
            .I(\ALU.addsub_7 ));
    InMux I__1322 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__1321 (
            .O(N__8486),
            .I(\ALU.mult_7 ));
    InMux I__1320 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__1319 (
            .O(N__8480),
            .I(overflow));
    InMux I__1318 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__1317 (
            .O(N__8474),
            .I(N__8471));
    Odrv4 I__1316 (
            .O(N__8471),
            .I(N_91));
    InMux I__1315 (
            .O(N__8468),
            .I(N__8465));
    LocalMux I__1314 (
            .O(N__8465),
            .I(res_13));
    InMux I__1313 (
            .O(N__8462),
            .I(N__8459));
    LocalMux I__1312 (
            .O(N__8459),
            .I(res_5));
    IoInMux I__1311 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__1310 (
            .O(N__8453),
            .I(N__8450));
    IoSpan4Mux I__1309 (
            .O(N__8450),
            .I(N__8447));
    Span4Mux_s3_h I__1308 (
            .O(N__8447),
            .I(N__8444));
    Span4Mux_h I__1307 (
            .O(N__8444),
            .I(N__8441));
    Span4Mux_h I__1306 (
            .O(N__8441),
            .I(N__8438));
    Sp12to4 I__1305 (
            .O(N__8438),
            .I(N__8434));
    InMux I__1304 (
            .O(N__8437),
            .I(N__8431));
    Span12Mux_v I__1303 (
            .O(N__8434),
            .I(N__8426));
    LocalMux I__1302 (
            .O(N__8431),
            .I(N__8426));
    Odrv12 I__1301 (
            .O(N__8426),
            .I(GPIO2_c));
    CascadeMux I__1300 (
            .O(N__8423),
            .I(N__8420));
    InMux I__1299 (
            .O(N__8420),
            .I(N__8417));
    LocalMux I__1298 (
            .O(N__8417),
            .I(res_10));
    InMux I__1297 (
            .O(N__8414),
            .I(\ALU.regsA_result_cry_0 ));
    InMux I__1296 (
            .O(N__8411),
            .I(N__8408));
    LocalMux I__1295 (
            .O(N__8408),
            .I(N__8405));
    Span4Mux_v I__1294 (
            .O(N__8405),
            .I(N__8402));
    Odrv4 I__1293 (
            .O(N__8402),
            .I(\ALU.mult_6 ));
    InMux I__1292 (
            .O(N__8399),
            .I(\ALU.regsA_result_cry_1_0 ));
    InMux I__1291 (
            .O(N__8396),
            .I(\ALU.regsA_result_cry_2_1 ));
    CascadeMux I__1290 (
            .O(N__8393),
            .I(N__8390));
    InMux I__1289 (
            .O(N__8390),
            .I(N__8387));
    LocalMux I__1288 (
            .O(N__8387),
            .I(N__8383));
    InMux I__1287 (
            .O(N__8386),
            .I(N__8380));
    Span4Mux_v I__1286 (
            .O(N__8383),
            .I(N__8377));
    LocalMux I__1285 (
            .O(N__8380),
            .I(\ALU.mult_AdderTree2_bigtree_932 ));
    Odrv4 I__1284 (
            .O(N__8377),
            .I(\ALU.mult_AdderTree2_bigtree_932 ));
    InMux I__1283 (
            .O(N__8372),
            .I(\ALU.regsA_result_cry_3_1 ));
    CascadeMux I__1282 (
            .O(N__8369),
            .I(N__8366));
    InMux I__1281 (
            .O(N__8366),
            .I(N__8363));
    LocalMux I__1280 (
            .O(N__8363),
            .I(N__8360));
    Span4Mux_v I__1279 (
            .O(N__8360),
            .I(N__8357));
    Odrv4 I__1278 (
            .O(N__8357),
            .I(\ALU.mult_AdderTree2_bigtree_933 ));
    InMux I__1277 (
            .O(N__8354),
            .I(\ALU.regsA_result_cry_4_0 ));
    CascadeMux I__1276 (
            .O(N__8351),
            .I(N__8347));
    CascadeMux I__1275 (
            .O(N__8350),
            .I(N__8344));
    InMux I__1274 (
            .O(N__8347),
            .I(N__8341));
    InMux I__1273 (
            .O(N__8344),
            .I(N__8338));
    LocalMux I__1272 (
            .O(N__8341),
            .I(N__8335));
    LocalMux I__1271 (
            .O(N__8338),
            .I(N__8332));
    Span4Mux_h I__1270 (
            .O(N__8335),
            .I(N__8329));
    Span4Mux_h I__1269 (
            .O(N__8332),
            .I(N__8326));
    Odrv4 I__1268 (
            .O(N__8329),
            .I(\ALU.mult_AdderTree2_bigtree_934 ));
    Odrv4 I__1267 (
            .O(N__8326),
            .I(\ALU.mult_AdderTree2_bigtree_934 ));
    InMux I__1266 (
            .O(N__8321),
            .I(\ALU.regsA_result_cry_5_1 ));
    InMux I__1265 (
            .O(N__8318),
            .I(N__8314));
    CascadeMux I__1264 (
            .O(N__8317),
            .I(N__8311));
    LocalMux I__1263 (
            .O(N__8314),
            .I(N__8308));
    InMux I__1262 (
            .O(N__8311),
            .I(N__8305));
    Span4Mux_v I__1261 (
            .O(N__8308),
            .I(N__8302));
    LocalMux I__1260 (
            .O(N__8305),
            .I(N__8299));
    Span4Mux_v I__1259 (
            .O(N__8302),
            .I(N__8296));
    Span4Mux_h I__1258 (
            .O(N__8299),
            .I(N__8293));
    Odrv4 I__1257 (
            .O(N__8296),
            .I(\ALU.mult_AdderTree2_bigtree_935 ));
    Odrv4 I__1256 (
            .O(N__8293),
            .I(\ALU.mult_AdderTree2_bigtree_935 ));
    InMux I__1255 (
            .O(N__8288),
            .I(\ALU.regsA_result_cry_6_0 ));
    CascadeMux I__1254 (
            .O(N__8285),
            .I(N__8282));
    InMux I__1253 (
            .O(N__8282),
            .I(N__8278));
    CascadeMux I__1252 (
            .O(N__8281),
            .I(N__8275));
    LocalMux I__1251 (
            .O(N__8278),
            .I(N__8272));
    InMux I__1250 (
            .O(N__8275),
            .I(N__8269));
    Span4Mux_v I__1249 (
            .O(N__8272),
            .I(N__8266));
    LocalMux I__1248 (
            .O(N__8269),
            .I(N__8263));
    Odrv4 I__1247 (
            .O(N__8266),
            .I(\ALU.mult_AdderTree2_bigtree_936 ));
    Odrv4 I__1246 (
            .O(N__8263),
            .I(\ALU.mult_AdderTree2_bigtree_936 ));
    InMux I__1245 (
            .O(N__8258),
            .I(bfn_12_16_0_));
    InMux I__1244 (
            .O(N__8255),
            .I(N__8251));
    InMux I__1243 (
            .O(N__8254),
            .I(N__8248));
    LocalMux I__1242 (
            .O(N__8251),
            .I(N__8245));
    LocalMux I__1241 (
            .O(N__8248),
            .I(N__8242));
    Span4Mux_h I__1240 (
            .O(N__8245),
            .I(N__8239));
    Span4Mux_h I__1239 (
            .O(N__8242),
            .I(N__8236));
    Odrv4 I__1238 (
            .O(N__8239),
            .I(\ALU.mult_AdderTree2_bigtree_937 ));
    Odrv4 I__1237 (
            .O(N__8236),
            .I(\ALU.mult_AdderTree2_bigtree_937 ));
    InMux I__1236 (
            .O(N__8231),
            .I(\ALU.regsA_result_cry_8 ));
    InMux I__1235 (
            .O(N__8228),
            .I(N__8225));
    LocalMux I__1234 (
            .O(N__8225),
            .I(\ALU.regsA_result_axb_14_l_ofx ));
    CascadeMux I__1233 (
            .O(N__8222),
            .I(N__8219));
    InMux I__1232 (
            .O(N__8219),
            .I(N__8216));
    LocalMux I__1231 (
            .O(N__8216),
            .I(\ALU.addsub_axb_7_l_ofxZ0 ));
    InMux I__1230 (
            .O(N__8213),
            .I(N__8210));
    LocalMux I__1229 (
            .O(N__8210),
            .I(N__8207));
    Odrv12 I__1228 (
            .O(N__8207),
            .I(\ALU.regsA_result_cry_8_ma ));
    InMux I__1227 (
            .O(N__8204),
            .I(N__8201));
    LocalMux I__1226 (
            .O(N__8201),
            .I(\ALU.regsA_result_axb_14_0 ));
    CascadeMux I__1225 (
            .O(N__8198),
            .I(N__8195));
    InMux I__1224 (
            .O(N__8195),
            .I(N__8192));
    LocalMux I__1223 (
            .O(N__8192),
            .I(\ALU.regsA_result_cry_14_ma ));
    CascadeMux I__1222 (
            .O(N__8189),
            .I(N__8186));
    InMux I__1221 (
            .O(N__8186),
            .I(N__8183));
    LocalMux I__1220 (
            .O(N__8183),
            .I(\ALU.addsub_axb_1_l_ofxZ0 ));
    InMux I__1219 (
            .O(N__8180),
            .I(N__8177));
    LocalMux I__1218 (
            .O(N__8177),
            .I(N__8173));
    CascadeMux I__1217 (
            .O(N__8176),
            .I(N__8170));
    Span4Mux_v I__1216 (
            .O(N__8173),
            .I(N__8165));
    InMux I__1215 (
            .O(N__8170),
            .I(N__8158));
    InMux I__1214 (
            .O(N__8169),
            .I(N__8158));
    InMux I__1213 (
            .O(N__8168),
            .I(N__8158));
    Span4Mux_v I__1212 (
            .O(N__8165),
            .I(N__8155));
    LocalMux I__1211 (
            .O(N__8158),
            .I(N__8152));
    Odrv4 I__1210 (
            .O(N__8155),
            .I(bZ0Z_15));
    Odrv12 I__1209 (
            .O(N__8152),
            .I(bZ0Z_15));
    InMux I__1208 (
            .O(N__8147),
            .I(N__8144));
    LocalMux I__1207 (
            .O(N__8144),
            .I(\ALU.overflow_RNOZ0Z_15 ));
    CascadeMux I__1206 (
            .O(N__8141),
            .I(N__8138));
    InMux I__1205 (
            .O(N__8138),
            .I(N__8135));
    LocalMux I__1204 (
            .O(N__8135),
            .I(\ALU.addsub_axb_0_l_ofxZ0 ));
    CascadeMux I__1203 (
            .O(N__8132),
            .I(N__8129));
    InMux I__1202 (
            .O(N__8129),
            .I(N__8126));
    LocalMux I__1201 (
            .O(N__8126),
            .I(\ALU.regsA_result_axb_7_l_ofx ));
    InMux I__1200 (
            .O(N__8123),
            .I(\ALU.regsA_result_cry_6_5 ));
    InMux I__1199 (
            .O(N__8120),
            .I(bfn_12_13_0_));
    InMux I__1198 (
            .O(N__8117),
            .I(\ALU.regsA_result_cry_8_2 ));
    InMux I__1197 (
            .O(N__8114),
            .I(\ALU.regsA_result_cry_9_3 ));
    InMux I__1196 (
            .O(N__8111),
            .I(\ALU.regsA_result_cry_10_2 ));
    InMux I__1195 (
            .O(N__8108),
            .I(\ALU.regsA_result_cry_11_3 ));
    InMux I__1194 (
            .O(N__8105),
            .I(\ALU.regsA_result_cry_12_0 ));
    InMux I__1193 (
            .O(N__8102),
            .I(\ALU.regsA_result_cry_13_1 ));
    InMux I__1192 (
            .O(N__8099),
            .I(\ALU.regsA_result_cry_14 ));
    CascadeMux I__1191 (
            .O(N__8096),
            .I(N__8093));
    InMux I__1190 (
            .O(N__8093),
            .I(N__8090));
    LocalMux I__1189 (
            .O(N__8090),
            .I(\ALU.regsA_result_cry_0_0_c_RNO ));
    InMux I__1188 (
            .O(N__8087),
            .I(N__8084));
    LocalMux I__1187 (
            .O(N__8084),
            .I(\ALU.regsA_result_axb_1_l_ofx ));
    InMux I__1186 (
            .O(N__8081),
            .I(\ALU.regsA_result_cry_0_2 ));
    CascadeMux I__1185 (
            .O(N__8078),
            .I(N__8075));
    InMux I__1184 (
            .O(N__8075),
            .I(N__8072));
    LocalMux I__1183 (
            .O(N__8072),
            .I(\ALU.regsA_result_axb_2_l_ofx ));
    InMux I__1182 (
            .O(N__8069),
            .I(\ALU.regsA_result_cry_1_3 ));
    InMux I__1181 (
            .O(N__8066),
            .I(N__8063));
    LocalMux I__1180 (
            .O(N__8063),
            .I(\ALU.regsA_result_cry_3_ma ));
    CascadeMux I__1179 (
            .O(N__8060),
            .I(N__8057));
    InMux I__1178 (
            .O(N__8057),
            .I(N__8054));
    LocalMux I__1177 (
            .O(N__8054),
            .I(\ALU.regsA_result_axb_3_l_ofx ));
    InMux I__1176 (
            .O(N__8051),
            .I(\ALU.regsA_result_cry_2_5 ));
    CascadeMux I__1175 (
            .O(N__8048),
            .I(N__8045));
    InMux I__1174 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__1173 (
            .O(N__8042),
            .I(\ALU.regsA_result_axb_4_l_ofx ));
    InMux I__1172 (
            .O(N__8039),
            .I(\ALU.regsA_result_cry_3_6 ));
    InMux I__1171 (
            .O(N__8036),
            .I(N__8033));
    LocalMux I__1170 (
            .O(N__8033),
            .I(\ALU.regsA_result_axb_5_l_ofx ));
    InMux I__1169 (
            .O(N__8030),
            .I(\ALU.regsA_result_cry_4_5 ));
    InMux I__1168 (
            .O(N__8027),
            .I(\ALU.regsA_result_cry_5_6 ));
    InMux I__1167 (
            .O(N__8024),
            .I(N__8021));
    LocalMux I__1166 (
            .O(N__8021),
            .I(N__8018));
    Odrv4 I__1165 (
            .O(N__8018),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_2 ));
    InMux I__1164 (
            .O(N__8015),
            .I(N__8012));
    LocalMux I__1163 (
            .O(N__8012),
            .I(N__8009));
    Span4Mux_v I__1162 (
            .O(N__8009),
            .I(N__8006));
    Odrv4 I__1161 (
            .O(N__8006),
            .I(\ALU.regsA_result_cry_2_ma_2 ));
    InMux I__1160 (
            .O(N__8003),
            .I(N__8000));
    LocalMux I__1159 (
            .O(N__8000),
            .I(N__7997));
    Odrv4 I__1158 (
            .O(N__7997),
            .I(\ALU.regsA_result_cry_3_ma_2 ));
    InMux I__1157 (
            .O(N__7994),
            .I(N__7991));
    LocalMux I__1156 (
            .O(N__7991),
            .I(N__7988));
    Odrv4 I__1155 (
            .O(N__7988),
            .I(\ALU.regsA_result_cry_4_ma_1 ));
    InMux I__1154 (
            .O(N__7985),
            .I(N__7981));
    InMux I__1153 (
            .O(N__7984),
            .I(N__7978));
    LocalMux I__1152 (
            .O(N__7981),
            .I(N__7973));
    LocalMux I__1151 (
            .O(N__7978),
            .I(N__7970));
    CascadeMux I__1150 (
            .O(N__7977),
            .I(N__7967));
    CascadeMux I__1149 (
            .O(N__7976),
            .I(N__7964));
    Span4Mux_h I__1148 (
            .O(N__7973),
            .I(N__7957));
    Span4Mux_h I__1147 (
            .O(N__7970),
            .I(N__7957));
    InMux I__1146 (
            .O(N__7967),
            .I(N__7954));
    InMux I__1145 (
            .O(N__7964),
            .I(N__7949));
    InMux I__1144 (
            .O(N__7963),
            .I(N__7949));
    CascadeMux I__1143 (
            .O(N__7962),
            .I(N__7946));
    Span4Mux_v I__1142 (
            .O(N__7957),
            .I(N__7942));
    LocalMux I__1141 (
            .O(N__7954),
            .I(N__7939));
    LocalMux I__1140 (
            .O(N__7949),
            .I(N__7936));
    InMux I__1139 (
            .O(N__7946),
            .I(N__7931));
    InMux I__1138 (
            .O(N__7945),
            .I(N__7931));
    Odrv4 I__1137 (
            .O(N__7942),
            .I(aZ0Z_14));
    Odrv4 I__1136 (
            .O(N__7939),
            .I(aZ0Z_14));
    Odrv12 I__1135 (
            .O(N__7936),
            .I(aZ0Z_14));
    LocalMux I__1134 (
            .O(N__7931),
            .I(aZ0Z_14));
    CascadeMux I__1133 (
            .O(N__7922),
            .I(N__7919));
    InMux I__1132 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__1131 (
            .O(N__7916),
            .I(N__7913));
    Span4Mux_v I__1130 (
            .O(N__7913),
            .I(N__7910));
    Odrv4 I__1129 (
            .O(N__7910),
            .I(\ALU.addsub_axb_14_l_ofxZ0 ));
    CascadeMux I__1128 (
            .O(N__7907),
            .I(N__7903));
    InMux I__1127 (
            .O(N__7906),
            .I(N__7900));
    InMux I__1126 (
            .O(N__7903),
            .I(N__7897));
    LocalMux I__1125 (
            .O(N__7900),
            .I(N__7892));
    LocalMux I__1124 (
            .O(N__7897),
            .I(N__7889));
    InMux I__1123 (
            .O(N__7896),
            .I(N__7886));
    CascadeMux I__1122 (
            .O(N__7895),
            .I(N__7883));
    Span4Mux_v I__1121 (
            .O(N__7892),
            .I(N__7870));
    Span4Mux_h I__1120 (
            .O(N__7889),
            .I(N__7870));
    LocalMux I__1119 (
            .O(N__7886),
            .I(N__7870));
    InMux I__1118 (
            .O(N__7883),
            .I(N__7865));
    InMux I__1117 (
            .O(N__7882),
            .I(N__7865));
    InMux I__1116 (
            .O(N__7881),
            .I(N__7862));
    CascadeMux I__1115 (
            .O(N__7880),
            .I(N__7859));
    CascadeMux I__1114 (
            .O(N__7879),
            .I(N__7856));
    CascadeMux I__1113 (
            .O(N__7878),
            .I(N__7852));
    InMux I__1112 (
            .O(N__7877),
            .I(N__7848));
    Span4Mux_v I__1111 (
            .O(N__7870),
            .I(N__7843));
    LocalMux I__1110 (
            .O(N__7865),
            .I(N__7843));
    LocalMux I__1109 (
            .O(N__7862),
            .I(N__7840));
    InMux I__1108 (
            .O(N__7859),
            .I(N__7829));
    InMux I__1107 (
            .O(N__7856),
            .I(N__7829));
    InMux I__1106 (
            .O(N__7855),
            .I(N__7829));
    InMux I__1105 (
            .O(N__7852),
            .I(N__7829));
    InMux I__1104 (
            .O(N__7851),
            .I(N__7829));
    LocalMux I__1103 (
            .O(N__7848),
            .I(aZ0Z_8));
    Odrv4 I__1102 (
            .O(N__7843),
            .I(aZ0Z_8));
    Odrv4 I__1101 (
            .O(N__7840),
            .I(aZ0Z_8));
    LocalMux I__1100 (
            .O(N__7829),
            .I(aZ0Z_8));
    CascadeMux I__1099 (
            .O(N__7820),
            .I(N__7817));
    InMux I__1098 (
            .O(N__7817),
            .I(N__7814));
    LocalMux I__1097 (
            .O(N__7814),
            .I(N__7811));
    Span4Mux_v I__1096 (
            .O(N__7811),
            .I(N__7808));
    Odrv4 I__1095 (
            .O(N__7808),
            .I(\ALU.addsub_axb_8_l_ofxZ0 ));
    InMux I__1094 (
            .O(N__7805),
            .I(N__7802));
    LocalMux I__1093 (
            .O(N__7802),
            .I(N__7799));
    Span4Mux_v I__1092 (
            .O(N__7799),
            .I(N__7796));
    Odrv4 I__1091 (
            .O(N__7796),
            .I(\ALU.addsub_axb_9_l_ofxZ0 ));
    CascadeMux I__1090 (
            .O(N__7793),
            .I(N__7790));
    InMux I__1089 (
            .O(N__7790),
            .I(N__7785));
    InMux I__1088 (
            .O(N__7789),
            .I(N__7782));
    InMux I__1087 (
            .O(N__7788),
            .I(N__7778));
    LocalMux I__1086 (
            .O(N__7785),
            .I(N__7775));
    LocalMux I__1085 (
            .O(N__7782),
            .I(N__7772));
    InMux I__1084 (
            .O(N__7781),
            .I(N__7769));
    LocalMux I__1083 (
            .O(N__7778),
            .I(N__7764));
    Span4Mux_v I__1082 (
            .O(N__7775),
            .I(N__7751));
    Span4Mux_h I__1081 (
            .O(N__7772),
            .I(N__7751));
    LocalMux I__1080 (
            .O(N__7769),
            .I(N__7751));
    CascadeMux I__1079 (
            .O(N__7768),
            .I(N__7744));
    CascadeMux I__1078 (
            .O(N__7767),
            .I(N__7740));
    Span12Mux_s11_h I__1077 (
            .O(N__7764),
            .I(N__7736));
    InMux I__1076 (
            .O(N__7763),
            .I(N__7725));
    InMux I__1075 (
            .O(N__7762),
            .I(N__7725));
    InMux I__1074 (
            .O(N__7761),
            .I(N__7725));
    InMux I__1073 (
            .O(N__7760),
            .I(N__7725));
    InMux I__1072 (
            .O(N__7759),
            .I(N__7725));
    InMux I__1071 (
            .O(N__7758),
            .I(N__7722));
    Span4Mux_v I__1070 (
            .O(N__7751),
            .I(N__7719));
    InMux I__1069 (
            .O(N__7750),
            .I(N__7714));
    InMux I__1068 (
            .O(N__7749),
            .I(N__7714));
    InMux I__1067 (
            .O(N__7748),
            .I(N__7701));
    InMux I__1066 (
            .O(N__7747),
            .I(N__7701));
    InMux I__1065 (
            .O(N__7744),
            .I(N__7701));
    InMux I__1064 (
            .O(N__7743),
            .I(N__7701));
    InMux I__1063 (
            .O(N__7740),
            .I(N__7701));
    InMux I__1062 (
            .O(N__7739),
            .I(N__7701));
    Odrv12 I__1061 (
            .O(N__7736),
            .I(aZ0Z_9));
    LocalMux I__1060 (
            .O(N__7725),
            .I(aZ0Z_9));
    LocalMux I__1059 (
            .O(N__7722),
            .I(aZ0Z_9));
    Odrv4 I__1058 (
            .O(N__7719),
            .I(aZ0Z_9));
    LocalMux I__1057 (
            .O(N__7714),
            .I(aZ0Z_9));
    LocalMux I__1056 (
            .O(N__7701),
            .I(aZ0Z_9));
    CascadeMux I__1055 (
            .O(N__7688),
            .I(N__7685));
    InMux I__1054 (
            .O(N__7685),
            .I(N__7682));
    LocalMux I__1053 (
            .O(N__7682),
            .I(\ALU.regsA_result_cry_5_ma_1 ));
    InMux I__1052 (
            .O(N__7679),
            .I(N__7676));
    LocalMux I__1051 (
            .O(N__7676),
            .I(\ALU.addsub_15 ));
    InMux I__1050 (
            .O(N__7673),
            .I(N__7670));
    LocalMux I__1049 (
            .O(N__7670),
            .I(\ALU.mult_15 ));
    InMux I__1048 (
            .O(N__7667),
            .I(N__7664));
    LocalMux I__1047 (
            .O(N__7664),
            .I(N__7661));
    Span4Mux_v I__1046 (
            .O(N__7661),
            .I(N__7658));
    Odrv4 I__1045 (
            .O(N__7658),
            .I(\ALU.addsub_6 ));
    CascadeMux I__1044 (
            .O(N__7655),
            .I(\ALU.mult_2_cascade_ ));
    InMux I__1043 (
            .O(N__7652),
            .I(N__7649));
    LocalMux I__1042 (
            .O(N__7649),
            .I(N__7646));
    Span4Mux_v I__1041 (
            .O(N__7646),
            .I(N__7643));
    Odrv4 I__1040 (
            .O(N__7643),
            .I(\ALU.addsub_2 ));
    InMux I__1039 (
            .O(N__7640),
            .I(N__7637));
    LocalMux I__1038 (
            .O(N__7637),
            .I(N__7634));
    Odrv4 I__1037 (
            .O(N__7634),
            .I(\ALU.regsA_result_cry_7_ma_0 ));
    CascadeMux I__1036 (
            .O(N__7631),
            .I(N__7628));
    InMux I__1035 (
            .O(N__7628),
            .I(N__7625));
    LocalMux I__1034 (
            .O(N__7625),
            .I(\ALU.regsA_result_axb_7_l_ofx_0 ));
    CascadeMux I__1033 (
            .O(N__7622),
            .I(N__7619));
    InMux I__1032 (
            .O(N__7619),
            .I(N__7616));
    LocalMux I__1031 (
            .O(N__7616),
            .I(\ALU.regsA_result_axb_8_1 ));
    InMux I__1030 (
            .O(N__7613),
            .I(N__7609));
    InMux I__1029 (
            .O(N__7612),
            .I(N__7606));
    LocalMux I__1028 (
            .O(N__7609),
            .I(N__7603));
    LocalMux I__1027 (
            .O(N__7606),
            .I(N__7600));
    Span4Mux_h I__1026 (
            .O(N__7603),
            .I(N__7597));
    Odrv4 I__1025 (
            .O(N__7600),
            .I(\ALU.mult_ab_128 ));
    Odrv4 I__1024 (
            .O(N__7597),
            .I(\ALU.mult_ab_128 ));
    CascadeMux I__1023 (
            .O(N__7592),
            .I(N__7589));
    InMux I__1022 (
            .O(N__7589),
            .I(N__7586));
    LocalMux I__1021 (
            .O(N__7586),
            .I(\ALU.addsub_8 ));
    InMux I__1020 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__1019 (
            .O(N__7580),
            .I(N__7577));
    Span4Mux_v I__1018 (
            .O(N__7577),
            .I(N__7574));
    Odrv4 I__1017 (
            .O(N__7574),
            .I(res_8));
    InMux I__1016 (
            .O(N__7571),
            .I(N__7568));
    LocalMux I__1015 (
            .O(N__7568),
            .I(\ALU.addsub_11 ));
    InMux I__1014 (
            .O(N__7565),
            .I(N__7562));
    LocalMux I__1013 (
            .O(N__7562),
            .I(\ALU.mult_11 ));
    InMux I__1012 (
            .O(N__7559),
            .I(N__7556));
    LocalMux I__1011 (
            .O(N__7556),
            .I(N__7553));
    Odrv4 I__1010 (
            .O(N__7553),
            .I(\ALU.addsub_0 ));
    IoInMux I__1009 (
            .O(N__7550),
            .I(N__7547));
    LocalMux I__1008 (
            .O(N__7547),
            .I(N__7543));
    InMux I__1007 (
            .O(N__7546),
            .I(N__7540));
    Span12Mux_s4_v I__1006 (
            .O(N__7543),
            .I(N__7537));
    LocalMux I__1005 (
            .O(N__7540),
            .I(N__7534));
    Span12Mux_v I__1004 (
            .O(N__7537),
            .I(N__7531));
    Span4Mux_h I__1003 (
            .O(N__7534),
            .I(N__7528));
    Odrv12 I__1002 (
            .O(N__7531),
            .I(GPIO0_c));
    Odrv4 I__1001 (
            .O(N__7528),
            .I(GPIO0_c));
    InMux I__1000 (
            .O(N__7523),
            .I(N__7520));
    LocalMux I__999 (
            .O(N__7520),
            .I(\ALU.addsub_13 ));
    InMux I__998 (
            .O(N__7517),
            .I(N__7514));
    LocalMux I__997 (
            .O(N__7514),
            .I(\ALU.mult_13 ));
    InMux I__996 (
            .O(N__7511),
            .I(N__7508));
    LocalMux I__995 (
            .O(N__7508),
            .I(N__7505));
    Odrv4 I__994 (
            .O(N__7505),
            .I(\ALU.addsub_12 ));
    InMux I__993 (
            .O(N__7502),
            .I(N__7499));
    LocalMux I__992 (
            .O(N__7499),
            .I(\ALU.mult_12 ));
    InMux I__991 (
            .O(N__7496),
            .I(N__7493));
    LocalMux I__990 (
            .O(N__7493),
            .I(\ALU.mult_1 ));
    InMux I__989 (
            .O(N__7490),
            .I(N__7487));
    LocalMux I__988 (
            .O(N__7487),
            .I(N__7484));
    Odrv4 I__987 (
            .O(N__7484),
            .I(\ALU.addsub_1 ));
    InMux I__986 (
            .O(N__7481),
            .I(N__7478));
    LocalMux I__985 (
            .O(N__7478),
            .I(N__7475));
    Odrv4 I__984 (
            .O(N__7475),
            .I(\ALU.addsub_9 ));
    InMux I__983 (
            .O(N__7472),
            .I(N__7469));
    LocalMux I__982 (
            .O(N__7469),
            .I(\ALU.mult_9 ));
    InMux I__981 (
            .O(N__7466),
            .I(N__7463));
    LocalMux I__980 (
            .O(N__7463),
            .I(N__7460));
    Odrv4 I__979 (
            .O(N__7460),
            .I(\ALU.addsub_10 ));
    InMux I__978 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__977 (
            .O(N__7454),
            .I(\ALU.mult_10 ));
    CascadeMux I__976 (
            .O(N__7451),
            .I(N__7447));
    InMux I__975 (
            .O(N__7450),
            .I(N__7442));
    InMux I__974 (
            .O(N__7447),
            .I(N__7437));
    InMux I__973 (
            .O(N__7446),
            .I(N__7437));
    CascadeMux I__972 (
            .O(N__7445),
            .I(N__7432));
    LocalMux I__971 (
            .O(N__7442),
            .I(N__7427));
    LocalMux I__970 (
            .O(N__7437),
            .I(N__7427));
    InMux I__969 (
            .O(N__7436),
            .I(N__7422));
    InMux I__968 (
            .O(N__7435),
            .I(N__7422));
    InMux I__967 (
            .O(N__7432),
            .I(N__7416));
    Sp12to4 I__966 (
            .O(N__7427),
            .I(N__7411));
    LocalMux I__965 (
            .O(N__7422),
            .I(N__7411));
    InMux I__964 (
            .O(N__7421),
            .I(N__7404));
    InMux I__963 (
            .O(N__7420),
            .I(N__7404));
    InMux I__962 (
            .O(N__7419),
            .I(N__7404));
    LocalMux I__961 (
            .O(N__7416),
            .I(aZ0Z_10));
    Odrv12 I__960 (
            .O(N__7411),
            .I(aZ0Z_10));
    LocalMux I__959 (
            .O(N__7404),
            .I(aZ0Z_10));
    CascadeMux I__958 (
            .O(N__7397),
            .I(N__7394));
    InMux I__957 (
            .O(N__7394),
            .I(N__7391));
    LocalMux I__956 (
            .O(N__7391),
            .I(\ALU.addsub_axb_10_l_ofxZ0 ));
    InMux I__955 (
            .O(N__7388),
            .I(\ALU.addsub_cry_9 ));
    InMux I__954 (
            .O(N__7385),
            .I(\ALU.addsub_cry_10 ));
    InMux I__953 (
            .O(N__7382),
            .I(N__7378));
    InMux I__952 (
            .O(N__7381),
            .I(N__7375));
    LocalMux I__951 (
            .O(N__7378),
            .I(N__7369));
    LocalMux I__950 (
            .O(N__7375),
            .I(N__7366));
    InMux I__949 (
            .O(N__7374),
            .I(N__7363));
    CascadeMux I__948 (
            .O(N__7373),
            .I(N__7358));
    CascadeMux I__947 (
            .O(N__7372),
            .I(N__7354));
    Span4Mux_v I__946 (
            .O(N__7369),
            .I(N__7350));
    Span4Mux_h I__945 (
            .O(N__7366),
            .I(N__7345));
    LocalMux I__944 (
            .O(N__7363),
            .I(N__7345));
    InMux I__943 (
            .O(N__7362),
            .I(N__7342));
    InMux I__942 (
            .O(N__7361),
            .I(N__7339));
    InMux I__941 (
            .O(N__7358),
            .I(N__7334));
    InMux I__940 (
            .O(N__7357),
            .I(N__7334));
    InMux I__939 (
            .O(N__7354),
            .I(N__7329));
    InMux I__938 (
            .O(N__7353),
            .I(N__7329));
    Odrv4 I__937 (
            .O(N__7350),
            .I(aZ0Z_12));
    Odrv4 I__936 (
            .O(N__7345),
            .I(aZ0Z_12));
    LocalMux I__935 (
            .O(N__7342),
            .I(aZ0Z_12));
    LocalMux I__934 (
            .O(N__7339),
            .I(aZ0Z_12));
    LocalMux I__933 (
            .O(N__7334),
            .I(aZ0Z_12));
    LocalMux I__932 (
            .O(N__7329),
            .I(aZ0Z_12));
    CascadeMux I__931 (
            .O(N__7316),
            .I(N__7313));
    InMux I__930 (
            .O(N__7313),
            .I(N__7310));
    LocalMux I__929 (
            .O(N__7310),
            .I(N__7307));
    Odrv12 I__928 (
            .O(N__7307),
            .I(\ALU.addsub_axb_12_l_ofxZ0 ));
    InMux I__927 (
            .O(N__7304),
            .I(\ALU.addsub_cry_11 ));
    InMux I__926 (
            .O(N__7301),
            .I(\ALU.addsub_cry_12 ));
    InMux I__925 (
            .O(N__7298),
            .I(\ALU.addsub_cry_13 ));
    InMux I__924 (
            .O(N__7295),
            .I(N__7291));
    InMux I__923 (
            .O(N__7294),
            .I(N__7286));
    LocalMux I__922 (
            .O(N__7291),
            .I(N__7283));
    InMux I__921 (
            .O(N__7290),
            .I(N__7276));
    InMux I__920 (
            .O(N__7289),
            .I(N__7276));
    LocalMux I__919 (
            .O(N__7286),
            .I(N__7273));
    Span12Mux_v I__918 (
            .O(N__7283),
            .I(N__7270));
    InMux I__917 (
            .O(N__7282),
            .I(N__7265));
    InMux I__916 (
            .O(N__7281),
            .I(N__7265));
    LocalMux I__915 (
            .O(N__7276),
            .I(N__7262));
    Odrv12 I__914 (
            .O(N__7273),
            .I(aZ0Z_15));
    Odrv12 I__913 (
            .O(N__7270),
            .I(aZ0Z_15));
    LocalMux I__912 (
            .O(N__7265),
            .I(aZ0Z_15));
    Odrv4 I__911 (
            .O(N__7262),
            .I(aZ0Z_15));
    CascadeMux I__910 (
            .O(N__7253),
            .I(N__7250));
    InMux I__909 (
            .O(N__7250),
            .I(N__7247));
    LocalMux I__908 (
            .O(N__7247),
            .I(N__7244));
    Odrv4 I__907 (
            .O(N__7244),
            .I(\ALU.addsub_axb_15_l_ofxZ0 ));
    InMux I__906 (
            .O(N__7241),
            .I(bfn_11_16_0_));
    InMux I__905 (
            .O(N__7238),
            .I(N__7235));
    LocalMux I__904 (
            .O(N__7235),
            .I(\ALU.mult_16 ));
    InMux I__903 (
            .O(N__7232),
            .I(\ALU.addsub_cry_15 ));
    InMux I__902 (
            .O(N__7229),
            .I(N__7226));
    LocalMux I__901 (
            .O(N__7226),
            .I(\ALU.addsub_14 ));
    InMux I__900 (
            .O(N__7223),
            .I(N__7220));
    LocalMux I__899 (
            .O(N__7220),
            .I(\ALU.mult_14 ));
    InMux I__898 (
            .O(N__7217),
            .I(\ALU.addsub_cry_0 ));
    CascadeMux I__897 (
            .O(N__7214),
            .I(N__7211));
    InMux I__896 (
            .O(N__7211),
            .I(N__7208));
    LocalMux I__895 (
            .O(N__7208),
            .I(\ALU.addsub_axb_2_l_ofxZ0 ));
    InMux I__894 (
            .O(N__7205),
            .I(\ALU.addsub_cry_1 ));
    InMux I__893 (
            .O(N__7202),
            .I(\ALU.addsub_cry_2 ));
    InMux I__892 (
            .O(N__7199),
            .I(\ALU.addsub_cry_3 ));
    InMux I__891 (
            .O(N__7196),
            .I(\ALU.addsub_cry_4 ));
    InMux I__890 (
            .O(N__7193),
            .I(\ALU.addsub_cry_5 ));
    InMux I__889 (
            .O(N__7190),
            .I(bfn_11_15_0_));
    InMux I__888 (
            .O(N__7187),
            .I(\ALU.addsub_cry_7 ));
    InMux I__887 (
            .O(N__7184),
            .I(\ALU.addsub_cry_8 ));
    InMux I__886 (
            .O(N__7181),
            .I(N__7178));
    LocalMux I__885 (
            .O(N__7178),
            .I(\ALU.regsA_result_axb_6 ));
    InMux I__884 (
            .O(N__7175),
            .I(N__7172));
    LocalMux I__883 (
            .O(N__7172),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_0 ));
    InMux I__882 (
            .O(N__7169),
            .I(\ALU.addsub_cry_0_c_THRU_CO ));
    CascadeMux I__881 (
            .O(N__7166),
            .I(N__7163));
    InMux I__880 (
            .O(N__7163),
            .I(N__7160));
    LocalMux I__879 (
            .O(N__7160),
            .I(\ALU.regsA_result_axb_6_l_ofx_0 ));
    CascadeMux I__878 (
            .O(N__7157),
            .I(N__7154));
    InMux I__877 (
            .O(N__7154),
            .I(N__7151));
    LocalMux I__876 (
            .O(N__7151),
            .I(\ALU.mult_AdderTree2_bigtree_674 ));
    InMux I__875 (
            .O(N__7148),
            .I(\ALU.regsA_result_cry_5_7 ));
    InMux I__874 (
            .O(N__7145),
            .I(N__7142));
    LocalMux I__873 (
            .O(N__7142),
            .I(\ALU.mult_AdderTree2_bigtree_675 ));
    InMux I__872 (
            .O(N__7139),
            .I(\ALU.regsA_result_cry_6_6 ));
    InMux I__871 (
            .O(N__7136),
            .I(N__7133));
    LocalMux I__870 (
            .O(N__7133),
            .I(\ALU.regsA_result_cry_5_0_THRU_CO ));
    InMux I__869 (
            .O(N__7130),
            .I(\ALU.regsA_result_cry_7_0 ));
    CascadeMux I__868 (
            .O(N__7127),
            .I(N__7124));
    InMux I__867 (
            .O(N__7124),
            .I(N__7121));
    LocalMux I__866 (
            .O(N__7121),
            .I(\ALU.regsA_result_axb_8_2 ));
    InMux I__865 (
            .O(N__7118),
            .I(N__7115));
    LocalMux I__864 (
            .O(N__7115),
            .I(N__7112));
    Odrv4 I__863 (
            .O(N__7112),
            .I(\ALU.regsA_result_cry_6_ma_0 ));
    InMux I__862 (
            .O(N__7109),
            .I(N__7106));
    LocalMux I__861 (
            .O(N__7106),
            .I(N__7101));
    CascadeMux I__860 (
            .O(N__7105),
            .I(N__7098));
    InMux I__859 (
            .O(N__7104),
            .I(N__7095));
    Span4Mux_v I__858 (
            .O(N__7101),
            .I(N__7092));
    InMux I__857 (
            .O(N__7098),
            .I(N__7089));
    LocalMux I__856 (
            .O(N__7095),
            .I(\ALU.mult_AdderTree2_bigtree_670 ));
    Odrv4 I__855 (
            .O(N__7092),
            .I(\ALU.mult_AdderTree2_bigtree_670 ));
    LocalMux I__854 (
            .O(N__7089),
            .I(\ALU.mult_AdderTree2_bigtree_670 ));
    InMux I__853 (
            .O(N__7082),
            .I(N__7079));
    LocalMux I__852 (
            .O(N__7079),
            .I(N__7076));
    Odrv4 I__851 (
            .O(N__7076),
            .I(\ALU.regsA_result_cry_2_c_RNO_0 ));
    InMux I__850 (
            .O(N__7073),
            .I(N__7070));
    LocalMux I__849 (
            .O(N__7070),
            .I(\ALU.regsA_result_cry_3_ma_0 ));
    CascadeMux I__848 (
            .O(N__7067),
            .I(N__7064));
    InMux I__847 (
            .O(N__7064),
            .I(N__7061));
    LocalMux I__846 (
            .O(N__7061),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_1 ));
    CascadeMux I__845 (
            .O(N__7058),
            .I(N__7055));
    InMux I__844 (
            .O(N__7055),
            .I(N__7052));
    LocalMux I__843 (
            .O(N__7052),
            .I(\ALU.regsA_result_axb_2_l_ofx_2 ));
    InMux I__842 (
            .O(N__7049),
            .I(\ALU.regsA_result_cry_1_6 ));
    CascadeMux I__841 (
            .O(N__7046),
            .I(N__7043));
    InMux I__840 (
            .O(N__7043),
            .I(N__7040));
    LocalMux I__839 (
            .O(N__7040),
            .I(\ALU.regsA_result_axb_3_l_ofx_2 ));
    CascadeMux I__838 (
            .O(N__7037),
            .I(N__7034));
    InMux I__837 (
            .O(N__7034),
            .I(N__7031));
    LocalMux I__836 (
            .O(N__7031),
            .I(\ALU.mult_AdderTree2_bigtree_671 ));
    InMux I__835 (
            .O(N__7028),
            .I(\ALU.regsA_result_cry_2_8 ));
    CascadeMux I__834 (
            .O(N__7025),
            .I(N__7022));
    InMux I__833 (
            .O(N__7022),
            .I(N__7019));
    LocalMux I__832 (
            .O(N__7019),
            .I(\ALU.regsA_result_axb_4_l_ofx_1 ));
    CascadeMux I__831 (
            .O(N__7016),
            .I(N__7013));
    InMux I__830 (
            .O(N__7013),
            .I(N__7010));
    LocalMux I__829 (
            .O(N__7010),
            .I(\ALU.mult_AdderTree2_bigtree_672 ));
    InMux I__828 (
            .O(N__7007),
            .I(\ALU.regsA_result_cry_3_8 ));
    InMux I__827 (
            .O(N__7004),
            .I(N__7001));
    LocalMux I__826 (
            .O(N__7001),
            .I(N__6998));
    Odrv4 I__825 (
            .O(N__6998),
            .I(\ALU.regsA_result_axb_5_l_ofx_1 ));
    CascadeMux I__824 (
            .O(N__6995),
            .I(N__6992));
    InMux I__823 (
            .O(N__6992),
            .I(N__6989));
    LocalMux I__822 (
            .O(N__6989),
            .I(\ALU.mult_AdderTree2_bigtree_673 ));
    InMux I__821 (
            .O(N__6986),
            .I(\ALU.regsA_result_cry_4_7 ));
    InMux I__820 (
            .O(N__6983),
            .I(bfn_10_17_0_));
    CascadeMux I__819 (
            .O(N__6980),
            .I(N__6977));
    InMux I__818 (
            .O(N__6977),
            .I(N__6973));
    InMux I__817 (
            .O(N__6976),
            .I(N__6970));
    LocalMux I__816 (
            .O(N__6973),
            .I(a_fastZ0Z_10));
    LocalMux I__815 (
            .O(N__6970),
            .I(a_fastZ0Z_10));
    CascadeMux I__814 (
            .O(N__6965),
            .I(N__6962));
    InMux I__813 (
            .O(N__6962),
            .I(N__6959));
    LocalMux I__812 (
            .O(N__6959),
            .I(\ALU.regsA_result_axb_2_l_ofx_1 ));
    CascadeMux I__811 (
            .O(N__6956),
            .I(N__6953));
    InMux I__810 (
            .O(N__6953),
            .I(N__6950));
    LocalMux I__809 (
            .O(N__6950),
            .I(\ALU.regsA_result_axb_3_l_ofx_1 ));
    CascadeMux I__808 (
            .O(N__6947),
            .I(N__6944));
    InMux I__807 (
            .O(N__6944),
            .I(N__6941));
    LocalMux I__806 (
            .O(N__6941),
            .I(N__6938));
    Odrv4 I__805 (
            .O(N__6938),
            .I(\ALU.regsA_result_axb_5_l_ofx_0 ));
    InMux I__804 (
            .O(N__6935),
            .I(N__6932));
    LocalMux I__803 (
            .O(N__6932),
            .I(N__6929));
    Odrv4 I__802 (
            .O(N__6929),
            .I(\ALU.mult_AdderTree2_bigtree_669 ));
    InMux I__801 (
            .O(N__6926),
            .I(\ALU.regsA_result_cry_0_0 ));
    InMux I__800 (
            .O(N__6923),
            .I(N__6920));
    LocalMux I__799 (
            .O(N__6920),
            .I(N__6917));
    Span4Mux_h I__798 (
            .O(N__6917),
            .I(N__6914));
    Odrv4 I__797 (
            .O(N__6914),
            .I(\ALU.regsA_result_cry_5_c_RNI073QE ));
    InMux I__796 (
            .O(N__6911),
            .I(\ALU.regsA_result_cry_1_1 ));
    InMux I__795 (
            .O(N__6908),
            .I(N__6905));
    LocalMux I__794 (
            .O(N__6905),
            .I(N__6902));
    Odrv12 I__793 (
            .O(N__6902),
            .I(\ALU.regsA_result_cry_2_c_RNIHNOEF ));
    InMux I__792 (
            .O(N__6899),
            .I(\ALU.regsA_result_cry_2_2 ));
    InMux I__791 (
            .O(N__6896),
            .I(N__6893));
    LocalMux I__790 (
            .O(N__6893),
            .I(\ALU.regsA_result_cry_7_c_RNI8EG3H ));
    InMux I__789 (
            .O(N__6890),
            .I(\ALU.regsA_result_cry_3_2 ));
    CascadeMux I__788 (
            .O(N__6887),
            .I(N__6884));
    InMux I__787 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__786 (
            .O(N__6881),
            .I(N__6878));
    Span4Mux_v I__785 (
            .O(N__6878),
            .I(N__6875));
    Odrv4 I__784 (
            .O(N__6875),
            .I(\ALU.regsA_result_cry_4_c_RNIA939H ));
    InMux I__783 (
            .O(N__6872),
            .I(\ALU.regsA_result_cry_4_1 ));
    CascadeMux I__782 (
            .O(N__6869),
            .I(N__6866));
    InMux I__781 (
            .O(N__6866),
            .I(N__6863));
    LocalMux I__780 (
            .O(N__6863),
            .I(N__6860));
    Span4Mux_v I__779 (
            .O(N__6860),
            .I(N__6857));
    Odrv4 I__778 (
            .O(N__6857),
            .I(\ALU.regsA_result_cry_5_c_RNIKCNNP ));
    InMux I__777 (
            .O(N__6854),
            .I(\ALU.regsA_result_cry_5_2 ));
    CascadeMux I__776 (
            .O(N__6851),
            .I(N__6848));
    InMux I__775 (
            .O(N__6848),
            .I(N__6845));
    LocalMux I__774 (
            .O(N__6845),
            .I(N__6842));
    Span4Mux_v I__773 (
            .O(N__6842),
            .I(N__6839));
    Odrv4 I__772 (
            .O(N__6839),
            .I(\ALU.regsA_result_cry_6_c_RNICICNO ));
    InMux I__771 (
            .O(N__6836),
            .I(\ALU.regsA_result_cry_6_1 ));
    CascadeMux I__770 (
            .O(N__6833),
            .I(N__6829));
    CascadeMux I__769 (
            .O(N__6832),
            .I(N__6826));
    InMux I__768 (
            .O(N__6829),
            .I(N__6818));
    InMux I__767 (
            .O(N__6826),
            .I(N__6818));
    InMux I__766 (
            .O(N__6825),
            .I(N__6818));
    LocalMux I__765 (
            .O(N__6818),
            .I(\FTDI.baudAccZ0Z_0 ));
    InMux I__764 (
            .O(N__6815),
            .I(N__6809));
    InMux I__763 (
            .O(N__6814),
            .I(N__6809));
    LocalMux I__762 (
            .O(N__6809),
            .I(N__6806));
    Odrv4 I__761 (
            .O(N__6806),
            .I(\FTDI.baudAccZ0Z_1 ));
    CascadeMux I__760 (
            .O(N__6803),
            .I(\FTDI.N_170_0_cascade_ ));
    CascadeMux I__759 (
            .O(N__6800),
            .I(\FTDI.TXstate_cnst_0_0_2_cascade_ ));
    InMux I__758 (
            .O(N__6797),
            .I(N__6793));
    CascadeMux I__757 (
            .O(N__6796),
            .I(N__6789));
    LocalMux I__756 (
            .O(N__6793),
            .I(N__6786));
    InMux I__755 (
            .O(N__6792),
            .I(N__6781));
    InMux I__754 (
            .O(N__6789),
            .I(N__6781));
    Odrv12 I__753 (
            .O(N__6786),
            .I(\ALU.mult_AdderTree2_bigtree_870 ));
    LocalMux I__752 (
            .O(N__6781),
            .I(\ALU.mult_AdderTree2_bigtree_870 ));
    CascadeMux I__751 (
            .O(N__6776),
            .I(N__6772));
    InMux I__750 (
            .O(N__6775),
            .I(N__6765));
    InMux I__749 (
            .O(N__6772),
            .I(N__6758));
    InMux I__748 (
            .O(N__6771),
            .I(N__6758));
    InMux I__747 (
            .O(N__6770),
            .I(N__6758));
    InMux I__746 (
            .O(N__6769),
            .I(N__6753));
    InMux I__745 (
            .O(N__6768),
            .I(N__6753));
    LocalMux I__744 (
            .O(N__6765),
            .I(\FTDI.TXstateZ0Z_1 ));
    LocalMux I__743 (
            .O(N__6758),
            .I(\FTDI.TXstateZ0Z_1 ));
    LocalMux I__742 (
            .O(N__6753),
            .I(\FTDI.TXstateZ0Z_1 ));
    CascadeMux I__741 (
            .O(N__6746),
            .I(N__6742));
    InMux I__740 (
            .O(N__6745),
            .I(N__6739));
    InMux I__739 (
            .O(N__6742),
            .I(N__6736));
    LocalMux I__738 (
            .O(N__6739),
            .I(\FTDI.TXstate_fastZ0Z_3 ));
    LocalMux I__737 (
            .O(N__6736),
            .I(\FTDI.TXstate_fastZ0Z_3 ));
    InMux I__736 (
            .O(N__6731),
            .I(N__6714));
    InMux I__735 (
            .O(N__6730),
            .I(N__6714));
    InMux I__734 (
            .O(N__6729),
            .I(N__6714));
    InMux I__733 (
            .O(N__6728),
            .I(N__6714));
    InMux I__732 (
            .O(N__6727),
            .I(N__6714));
    InMux I__731 (
            .O(N__6726),
            .I(N__6709));
    InMux I__730 (
            .O(N__6725),
            .I(N__6709));
    LocalMux I__729 (
            .O(N__6714),
            .I(\FTDI.TXstateZ0Z_0 ));
    LocalMux I__728 (
            .O(N__6709),
            .I(\FTDI.TXstateZ0Z_0 ));
    CascadeMux I__727 (
            .O(N__6704),
            .I(FTDI_TXready_cascade_));
    CascadeMux I__726 (
            .O(N__6701),
            .I(un1_testState31_0_cascade_));
    InMux I__725 (
            .O(N__6698),
            .I(N__6695));
    LocalMux I__724 (
            .O(N__6695),
            .I(\ALU.mult_AdderTree2_bigtree_741 ));
    InMux I__723 (
            .O(N__6692),
            .I(\ALU.regsA_result_cry_2_6 ));
    InMux I__722 (
            .O(N__6689),
            .I(N__6686));
    LocalMux I__721 (
            .O(N__6686),
            .I(N__6683));
    Span4Mux_h I__720 (
            .O(N__6683),
            .I(N__6680));
    Odrv4 I__719 (
            .O(N__6680),
            .I(\ALU.regsA_result_axb_2 ));
    InMux I__718 (
            .O(N__6677),
            .I(N__6674));
    LocalMux I__717 (
            .O(N__6674),
            .I(N__6671));
    Odrv4 I__716 (
            .O(N__6671),
            .I(\ALU.regsA_result_cry_1_THRU_CO ));
    InMux I__715 (
            .O(N__6668),
            .I(\ALU.regsA_result_cry_3 ));
    InMux I__714 (
            .O(N__6665),
            .I(N__6662));
    LocalMux I__713 (
            .O(N__6662),
            .I(N__6659));
    Odrv4 I__712 (
            .O(N__6659),
            .I(\ALU.regsA_result_axb_4_0 ));
    CascadeMux I__711 (
            .O(N__6656),
            .I(N__6653));
    InMux I__710 (
            .O(N__6653),
            .I(N__6650));
    LocalMux I__709 (
            .O(N__6650),
            .I(\ALU.regsA_result_axb_3_l_ofx_0 ));
    CascadeMux I__708 (
            .O(N__6647),
            .I(N__6644));
    InMux I__707 (
            .O(N__6644),
            .I(N__6641));
    LocalMux I__706 (
            .O(N__6641),
            .I(\ALU.regsA_result_axb_4 ));
    InMux I__705 (
            .O(N__6638),
            .I(N__6634));
    InMux I__704 (
            .O(N__6637),
            .I(N__6631));
    LocalMux I__703 (
            .O(N__6634),
            .I(\ALU.mult_AdderTree2_bigtree_873 ));
    LocalMux I__702 (
            .O(N__6631),
            .I(\ALU.mult_AdderTree2_bigtree_873 ));
    CascadeMux I__701 (
            .O(N__6626),
            .I(N__6623));
    InMux I__700 (
            .O(N__6623),
            .I(N__6620));
    LocalMux I__699 (
            .O(N__6620),
            .I(\ALU.regsA_result_cry_2_c_RNIC59KA ));
    InMux I__698 (
            .O(N__6617),
            .I(\ALU.regsA_result_cry_2 ));
    InMux I__697 (
            .O(N__6614),
            .I(\ALU.regsA_result_cry_3_0 ));
    InMux I__696 (
            .O(N__6611),
            .I(N__6608));
    LocalMux I__695 (
            .O(N__6608),
            .I(\ALU.regsA_result_cry_3_0_THRU_CO ));
    InMux I__694 (
            .O(N__6605),
            .I(N__6602));
    LocalMux I__693 (
            .O(N__6602),
            .I(\ALU.mult_AdderTree2_bigtree_739 ));
    CascadeMux I__692 (
            .O(N__6599),
            .I(N__6596));
    InMux I__691 (
            .O(N__6596),
            .I(N__6593));
    LocalMux I__690 (
            .O(N__6593),
            .I(\ALU.mult_AdderTree2_bigtree_774 ));
    InMux I__689 (
            .O(N__6590),
            .I(N__6587));
    LocalMux I__688 (
            .O(N__6587),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_3 ));
    CascadeMux I__687 (
            .O(N__6584),
            .I(N__6581));
    InMux I__686 (
            .O(N__6581),
            .I(N__6578));
    LocalMux I__685 (
            .O(N__6578),
            .I(\ALU.regsA_result_cry_1_0_c_RNO ));
    CascadeMux I__684 (
            .O(N__6575),
            .I(N__6572));
    InMux I__683 (
            .O(N__6572),
            .I(N__6569));
    LocalMux I__682 (
            .O(N__6569),
            .I(\ALU.regsA_result_axb_2_l_ofx_0 ));
    InMux I__681 (
            .O(N__6566),
            .I(N__6559));
    InMux I__680 (
            .O(N__6565),
            .I(N__6559));
    CascadeMux I__679 (
            .O(N__6564),
            .I(N__6556));
    LocalMux I__678 (
            .O(N__6559),
            .I(N__6553));
    InMux I__677 (
            .O(N__6556),
            .I(N__6550));
    Odrv4 I__676 (
            .O(N__6553),
            .I(\ALU.mult_AdderTree2_bigtree_740 ));
    LocalMux I__675 (
            .O(N__6550),
            .I(\ALU.mult_AdderTree2_bigtree_740 ));
    InMux I__674 (
            .O(N__6545),
            .I(\ALU.regsA_result_cry_1_4 ));
    InMux I__673 (
            .O(N__6542),
            .I(N__6539));
    LocalMux I__672 (
            .O(N__6539),
            .I(\ALU.regsA_result_cry_5_ma_0 ));
    InMux I__671 (
            .O(N__6536),
            .I(N__6533));
    LocalMux I__670 (
            .O(N__6533),
            .I(N__6530));
    Odrv4 I__669 (
            .O(N__6530),
            .I(\ALU.mult_AdderTree2_bigtree_704 ));
    InMux I__668 (
            .O(N__6527),
            .I(\ALU.regsA_result_cry_2_0 ));
    InMux I__667 (
            .O(N__6524),
            .I(N__6521));
    LocalMux I__666 (
            .O(N__6521),
            .I(\ALU.mult_AdderTree2_bigtree_705 ));
    InMux I__665 (
            .O(N__6518),
            .I(\ALU.regsA_result_cry_3_4 ));
    InMux I__664 (
            .O(N__6515),
            .I(N__6512));
    LocalMux I__663 (
            .O(N__6512),
            .I(N__6509));
    Odrv4 I__662 (
            .O(N__6509),
            .I(\ALU.mult_AdderTree2_bigtree_706 ));
    CascadeMux I__661 (
            .O(N__6506),
            .I(N__6503));
    InMux I__660 (
            .O(N__6503),
            .I(N__6500));
    LocalMux I__659 (
            .O(N__6500),
            .I(\ALU.mult_AdderTree2_bigtree_871 ));
    InMux I__658 (
            .O(N__6497),
            .I(\ALU.regsA_result_cry_4_3 ));
    InMux I__657 (
            .O(N__6494),
            .I(N__6491));
    LocalMux I__656 (
            .O(N__6491),
            .I(\ALU.mult_AdderTree2_bigtree_707 ));
    CascadeMux I__655 (
            .O(N__6488),
            .I(N__6484));
    InMux I__654 (
            .O(N__6487),
            .I(N__6481));
    InMux I__653 (
            .O(N__6484),
            .I(N__6478));
    LocalMux I__652 (
            .O(N__6481),
            .I(\ALU.mult_AdderTree2_bigtree_872 ));
    LocalMux I__651 (
            .O(N__6478),
            .I(\ALU.mult_AdderTree2_bigtree_872 ));
    InMux I__650 (
            .O(N__6473),
            .I(\ALU.regsA_result_cry_5_4 ));
    CascadeMux I__649 (
            .O(N__6470),
            .I(N__6467));
    InMux I__648 (
            .O(N__6467),
            .I(N__6464));
    LocalMux I__647 (
            .O(N__6464),
            .I(\ALU.mult_AdderTree2_bigtree_708 ));
    InMux I__646 (
            .O(N__6461),
            .I(\ALU.regsA_result_cry_6_3 ));
    InMux I__645 (
            .O(N__6458),
            .I(\ALU.regsA_result_cry_7_1 ));
    InMux I__644 (
            .O(N__6455),
            .I(N__6452));
    LocalMux I__643 (
            .O(N__6452),
            .I(\ALU.regsA_result_cry_2_c_RNO ));
    InMux I__642 (
            .O(N__6449),
            .I(N__6446));
    LocalMux I__641 (
            .O(N__6446),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0 ));
    CascadeMux I__640 (
            .O(N__6443),
            .I(N__6440));
    InMux I__639 (
            .O(N__6440),
            .I(N__6437));
    LocalMux I__638 (
            .O(N__6437),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_0_1 ));
    InMux I__637 (
            .O(N__6434),
            .I(N__6431));
    LocalMux I__636 (
            .O(N__6431),
            .I(N__6428));
    Odrv4 I__635 (
            .O(N__6428),
            .I(\ALU.regsA_result_cry_2_ma_1 ));
    InMux I__634 (
            .O(N__6425),
            .I(\ALU.regsA_result_cry_1_5 ));
    InMux I__633 (
            .O(N__6422),
            .I(N__6419));
    LocalMux I__632 (
            .O(N__6419),
            .I(N__6416));
    Odrv4 I__631 (
            .O(N__6416),
            .I(\ALU.regsA_result_cry_3_ma_1 ));
    InMux I__630 (
            .O(N__6413),
            .I(\ALU.regsA_result_cry_2_7 ));
    InMux I__629 (
            .O(N__6410),
            .I(N__6407));
    LocalMux I__628 (
            .O(N__6407),
            .I(\ALU.regsA_result_cry_4_ma_0 ));
    InMux I__627 (
            .O(N__6404),
            .I(\ALU.regsA_result_cry_3_7 ));
    InMux I__626 (
            .O(N__6401),
            .I(\ALU.regsA_result_cry_4_6 ));
    InMux I__625 (
            .O(N__6398),
            .I(\ALU.regsA_result_cry_5_0 ));
    CascadeMux I__624 (
            .O(N__6395),
            .I(N__6392));
    InMux I__623 (
            .O(N__6392),
            .I(N__6389));
    LocalMux I__622 (
            .O(N__6389),
            .I(\ALU.regsA_result_axb_4_l_ofx_0 ));
    InMux I__621 (
            .O(N__6386),
            .I(N__6383));
    LocalMux I__620 (
            .O(N__6383),
            .I(\FTDI.TXstate_RNIE1MMZ0Z_2 ));
    CascadeMux I__619 (
            .O(N__6380),
            .I(\FTDI.TXstate_RNIE1MMZ0Z_2_cascade_ ));
    InMux I__618 (
            .O(N__6377),
            .I(N__6374));
    LocalMux I__617 (
            .O(N__6374),
            .I(\ALU.regsA_result_cry_4_c_RNO ));
    InMux I__616 (
            .O(N__6371),
            .I(N__6368));
    LocalMux I__615 (
            .O(N__6368),
            .I(\ALU.regsA_result_cry_1_0_c_RNIKGQO9 ));
    CascadeMux I__614 (
            .O(N__6365),
            .I(\FTDI.i2_mux_cascade_ ));
    CascadeMux I__613 (
            .O(N__6362),
            .I(N__6359));
    InMux I__612 (
            .O(N__6359),
            .I(N__6356));
    LocalMux I__611 (
            .O(N__6356),
            .I(\ALU.regsA_result_cry_1_0_c_RNO_2 ));
    InMux I__610 (
            .O(N__6353),
            .I(\ALU.regsA_result_cry_1 ));
    InMux I__609 (
            .O(N__6350),
            .I(\ALU.regsA_result_cry_4 ));
    InMux I__608 (
            .O(N__6347),
            .I(\ALU.regsA_result_cry_5 ));
    InMux I__607 (
            .O(N__6344),
            .I(\ALU.regsA_result_cry_6 ));
    InMux I__606 (
            .O(N__6341),
            .I(\ALU.regsA_result_cry_7 ));
    InMux I__605 (
            .O(N__6338),
            .I(N__6335));
    LocalMux I__604 (
            .O(N__6335),
            .I(clkdivZ0Z_17));
    InMux I__603 (
            .O(N__6332),
            .I(clkdiv_cry_16));
    InMux I__602 (
            .O(N__6329),
            .I(N__6326));
    LocalMux I__601 (
            .O(N__6326),
            .I(clkdivZ0Z_18));
    InMux I__600 (
            .O(N__6323),
            .I(clkdiv_cry_17));
    InMux I__599 (
            .O(N__6320),
            .I(N__6317));
    LocalMux I__598 (
            .O(N__6317),
            .I(clkdivZ0Z_19));
    InMux I__597 (
            .O(N__6314),
            .I(clkdiv_cry_18));
    InMux I__596 (
            .O(N__6311),
            .I(N__6308));
    LocalMux I__595 (
            .O(N__6308),
            .I(clkdivZ0Z_20));
    InMux I__594 (
            .O(N__6305),
            .I(clkdiv_cry_19));
    InMux I__593 (
            .O(N__6302),
            .I(N__6299));
    LocalMux I__592 (
            .O(N__6299),
            .I(clkdivZ0Z_21));
    InMux I__591 (
            .O(N__6296),
            .I(clkdiv_cry_20));
    InMux I__590 (
            .O(N__6293),
            .I(N__6290));
    LocalMux I__589 (
            .O(N__6290),
            .I(clkdivZ0Z_22));
    InMux I__588 (
            .O(N__6287),
            .I(clkdiv_cry_21));
    InMux I__587 (
            .O(N__6284),
            .I(clkdiv_cry_22));
    IoInMux I__586 (
            .O(N__6281),
            .I(N__6278));
    LocalMux I__585 (
            .O(N__6278),
            .I(N__6275));
    Span12Mux_s10_v I__584 (
            .O(N__6275),
            .I(N__6271));
    InMux I__583 (
            .O(N__6274),
            .I(N__6268));
    Odrv12 I__582 (
            .O(N__6271),
            .I(GPIO3_c));
    LocalMux I__581 (
            .O(N__6268),
            .I(GPIO3_c));
    InMux I__580 (
            .O(N__6263),
            .I(N__6260));
    LocalMux I__579 (
            .O(N__6260),
            .I(clkdivZ0Z_8));
    InMux I__578 (
            .O(N__6257),
            .I(bfn_1_14_0_));
    InMux I__577 (
            .O(N__6254),
            .I(N__6251));
    LocalMux I__576 (
            .O(N__6251),
            .I(clkdivZ0Z_9));
    InMux I__575 (
            .O(N__6248),
            .I(clkdiv_cry_8));
    InMux I__574 (
            .O(N__6245),
            .I(N__6242));
    LocalMux I__573 (
            .O(N__6242),
            .I(clkdivZ0Z_10));
    InMux I__572 (
            .O(N__6239),
            .I(clkdiv_cry_9));
    InMux I__571 (
            .O(N__6236),
            .I(N__6233));
    LocalMux I__570 (
            .O(N__6233),
            .I(clkdivZ0Z_11));
    InMux I__569 (
            .O(N__6230),
            .I(clkdiv_cry_10));
    InMux I__568 (
            .O(N__6227),
            .I(N__6224));
    LocalMux I__567 (
            .O(N__6224),
            .I(clkdivZ0Z_12));
    InMux I__566 (
            .O(N__6221),
            .I(clkdiv_cry_11));
    InMux I__565 (
            .O(N__6218),
            .I(N__6215));
    LocalMux I__564 (
            .O(N__6215),
            .I(clkdivZ0Z_13));
    InMux I__563 (
            .O(N__6212),
            .I(clkdiv_cry_12));
    InMux I__562 (
            .O(N__6209),
            .I(N__6206));
    LocalMux I__561 (
            .O(N__6206),
            .I(clkdivZ0Z_14));
    InMux I__560 (
            .O(N__6203),
            .I(clkdiv_cry_13));
    InMux I__559 (
            .O(N__6200),
            .I(N__6197));
    LocalMux I__558 (
            .O(N__6197),
            .I(clkdivZ0Z_15));
    InMux I__557 (
            .O(N__6194),
            .I(clkdiv_cry_14));
    InMux I__556 (
            .O(N__6191),
            .I(N__6188));
    LocalMux I__555 (
            .O(N__6188),
            .I(clkdivZ0Z_16));
    InMux I__554 (
            .O(N__6185),
            .I(bfn_1_15_0_));
    InMux I__553 (
            .O(N__6182),
            .I(N__6179));
    LocalMux I__552 (
            .O(N__6179),
            .I(clkdivZ0Z_0));
    InMux I__551 (
            .O(N__6176),
            .I(bfn_1_13_0_));
    InMux I__550 (
            .O(N__6173),
            .I(N__6170));
    LocalMux I__549 (
            .O(N__6170),
            .I(clkdivZ0Z_1));
    InMux I__548 (
            .O(N__6167),
            .I(clkdiv_cry_0));
    InMux I__547 (
            .O(N__6164),
            .I(N__6161));
    LocalMux I__546 (
            .O(N__6161),
            .I(clkdivZ0Z_2));
    InMux I__545 (
            .O(N__6158),
            .I(clkdiv_cry_1));
    InMux I__544 (
            .O(N__6155),
            .I(N__6152));
    LocalMux I__543 (
            .O(N__6152),
            .I(clkdivZ0Z_3));
    InMux I__542 (
            .O(N__6149),
            .I(clkdiv_cry_2));
    InMux I__541 (
            .O(N__6146),
            .I(N__6143));
    LocalMux I__540 (
            .O(N__6143),
            .I(clkdivZ0Z_4));
    InMux I__539 (
            .O(N__6140),
            .I(clkdiv_cry_3));
    InMux I__538 (
            .O(N__6137),
            .I(N__6134));
    LocalMux I__537 (
            .O(N__6134),
            .I(clkdivZ0Z_5));
    InMux I__536 (
            .O(N__6131),
            .I(clkdiv_cry_4));
    InMux I__535 (
            .O(N__6128),
            .I(N__6125));
    LocalMux I__534 (
            .O(N__6125),
            .I(clkdivZ0Z_6));
    InMux I__533 (
            .O(N__6122),
            .I(clkdiv_cry_5));
    InMux I__532 (
            .O(N__6119),
            .I(N__6116));
    LocalMux I__531 (
            .O(N__6116),
            .I(clkdivZ0Z_7));
    InMux I__530 (
            .O(N__6113),
            .I(clkdiv_cry_6));
    INV \INVFTDI.gap_1C  (
            .O(\INVFTDI.gap_1C_net ),
            .I(N__16076));
    INV \INVFTDI.RXstate_2C  (
            .O(\INVFTDI.RXstate_2C_net ),
            .I(N__16074));
    INV \INVFTDI.RXstate_3C  (
            .O(\INVFTDI.RXstate_3C_net ),
            .I(N__16073));
    INV \INVFTDI.TXshift_7C  (
            .O(\INVFTDI.TXshift_7C_net ),
            .I(N__16110));
    INV \INVFTDI.RXbuffer_5C  (
            .O(\INVFTDI.RXbuffer_5C_net ),
            .I(N__16078));
    INV \INVFTDI.RXbuffer_2C  (
            .O(\INVFTDI.RXbuffer_2C_net ),
            .I(N__16075));
    INV \INVFTDI.TXshift_1C  (
            .O(\INVFTDI.TXshift_1C_net ),
            .I(N__16112));
    INV \INVFTDI.TXstate_2C  (
            .O(\INVFTDI.TXstate_2C_net ),
            .I(N__16117));
    INV \INVFTDI.baudAcc_0C  (
            .O(\INVFTDI.baudAcc_0C_net ),
            .I(N__16113));
    INV \INVFTDI.TXstate_0C  (
            .O(\INVFTDI.TXstate_0C_net ),
            .I(N__16121));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\ALU.addsub_cry_6 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\ALU.addsub_cry_14 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\ALU.regsA_result_cry_7_9 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\ALU.regsA_result_cry_7_2 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(\ALU.regsA_result_cry_9_2 ),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\ALU.regsA_result_cry_7_3 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\ALU.regsA_result_cry_8_5 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\ALU.regsA_result_cry_8_3 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\ALU.regsA_result_cry_8_4 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\ALU.regsA_result_cry_7_5 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(clkdiv_cry_7),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(clkdiv_cry_15),
            .carryinitout(bfn_1_15_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam clkdiv_0_LC_1_13_0.C_ON=1'b1;
    defparam clkdiv_0_LC_1_13_0.SEQ_MODE=4'b1000;
    defparam clkdiv_0_LC_1_13_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_0_LC_1_13_0 (
            .in0(_gnd_net_),
            .in1(N__6182),
            .in2(_gnd_net_),
            .in3(N__6176),
            .lcout(clkdivZ0Z_0),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(clkdiv_cry_0),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_1_LC_1_13_1.C_ON=1'b1;
    defparam clkdiv_1_LC_1_13_1.SEQ_MODE=4'b1000;
    defparam clkdiv_1_LC_1_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_1_LC_1_13_1 (
            .in0(_gnd_net_),
            .in1(N__6173),
            .in2(_gnd_net_),
            .in3(N__6167),
            .lcout(clkdivZ0Z_1),
            .ltout(),
            .carryin(clkdiv_cry_0),
            .carryout(clkdiv_cry_1),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_2_LC_1_13_2.C_ON=1'b1;
    defparam clkdiv_2_LC_1_13_2.SEQ_MODE=4'b1000;
    defparam clkdiv_2_LC_1_13_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_2_LC_1_13_2 (
            .in0(_gnd_net_),
            .in1(N__6164),
            .in2(_gnd_net_),
            .in3(N__6158),
            .lcout(clkdivZ0Z_2),
            .ltout(),
            .carryin(clkdiv_cry_1),
            .carryout(clkdiv_cry_2),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_3_LC_1_13_3.C_ON=1'b1;
    defparam clkdiv_3_LC_1_13_3.SEQ_MODE=4'b1000;
    defparam clkdiv_3_LC_1_13_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_3_LC_1_13_3 (
            .in0(_gnd_net_),
            .in1(N__6155),
            .in2(_gnd_net_),
            .in3(N__6149),
            .lcout(clkdivZ0Z_3),
            .ltout(),
            .carryin(clkdiv_cry_2),
            .carryout(clkdiv_cry_3),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_4_LC_1_13_4.C_ON=1'b1;
    defparam clkdiv_4_LC_1_13_4.SEQ_MODE=4'b1000;
    defparam clkdiv_4_LC_1_13_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_4_LC_1_13_4 (
            .in0(_gnd_net_),
            .in1(N__6146),
            .in2(_gnd_net_),
            .in3(N__6140),
            .lcout(clkdivZ0Z_4),
            .ltout(),
            .carryin(clkdiv_cry_3),
            .carryout(clkdiv_cry_4),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_5_LC_1_13_5.C_ON=1'b1;
    defparam clkdiv_5_LC_1_13_5.SEQ_MODE=4'b1000;
    defparam clkdiv_5_LC_1_13_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_5_LC_1_13_5 (
            .in0(_gnd_net_),
            .in1(N__6137),
            .in2(_gnd_net_),
            .in3(N__6131),
            .lcout(clkdivZ0Z_5),
            .ltout(),
            .carryin(clkdiv_cry_4),
            .carryout(clkdiv_cry_5),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_6_LC_1_13_6.C_ON=1'b1;
    defparam clkdiv_6_LC_1_13_6.SEQ_MODE=4'b1000;
    defparam clkdiv_6_LC_1_13_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_6_LC_1_13_6 (
            .in0(_gnd_net_),
            .in1(N__6128),
            .in2(_gnd_net_),
            .in3(N__6122),
            .lcout(clkdivZ0Z_6),
            .ltout(),
            .carryin(clkdiv_cry_5),
            .carryout(clkdiv_cry_6),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_7_LC_1_13_7.C_ON=1'b1;
    defparam clkdiv_7_LC_1_13_7.SEQ_MODE=4'b1000;
    defparam clkdiv_7_LC_1_13_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_7_LC_1_13_7 (
            .in0(_gnd_net_),
            .in1(N__6119),
            .in2(_gnd_net_),
            .in3(N__6113),
            .lcout(clkdivZ0Z_7),
            .ltout(),
            .carryin(clkdiv_cry_6),
            .carryout(clkdiv_cry_7),
            .clk(N__16122),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_8_LC_1_14_0.C_ON=1'b1;
    defparam clkdiv_8_LC_1_14_0.SEQ_MODE=4'b1000;
    defparam clkdiv_8_LC_1_14_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_8_LC_1_14_0 (
            .in0(_gnd_net_),
            .in1(N__6263),
            .in2(_gnd_net_),
            .in3(N__6257),
            .lcout(clkdivZ0Z_8),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(clkdiv_cry_8),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_9_LC_1_14_1.C_ON=1'b1;
    defparam clkdiv_9_LC_1_14_1.SEQ_MODE=4'b1000;
    defparam clkdiv_9_LC_1_14_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_9_LC_1_14_1 (
            .in0(_gnd_net_),
            .in1(N__6254),
            .in2(_gnd_net_),
            .in3(N__6248),
            .lcout(clkdivZ0Z_9),
            .ltout(),
            .carryin(clkdiv_cry_8),
            .carryout(clkdiv_cry_9),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_10_LC_1_14_2.C_ON=1'b1;
    defparam clkdiv_10_LC_1_14_2.SEQ_MODE=4'b1000;
    defparam clkdiv_10_LC_1_14_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_10_LC_1_14_2 (
            .in0(_gnd_net_),
            .in1(N__6245),
            .in2(_gnd_net_),
            .in3(N__6239),
            .lcout(clkdivZ0Z_10),
            .ltout(),
            .carryin(clkdiv_cry_9),
            .carryout(clkdiv_cry_10),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_11_LC_1_14_3.C_ON=1'b1;
    defparam clkdiv_11_LC_1_14_3.SEQ_MODE=4'b1000;
    defparam clkdiv_11_LC_1_14_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_11_LC_1_14_3 (
            .in0(_gnd_net_),
            .in1(N__6236),
            .in2(_gnd_net_),
            .in3(N__6230),
            .lcout(clkdivZ0Z_11),
            .ltout(),
            .carryin(clkdiv_cry_10),
            .carryout(clkdiv_cry_11),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_12_LC_1_14_4.C_ON=1'b1;
    defparam clkdiv_12_LC_1_14_4.SEQ_MODE=4'b1000;
    defparam clkdiv_12_LC_1_14_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_12_LC_1_14_4 (
            .in0(_gnd_net_),
            .in1(N__6227),
            .in2(_gnd_net_),
            .in3(N__6221),
            .lcout(clkdivZ0Z_12),
            .ltout(),
            .carryin(clkdiv_cry_11),
            .carryout(clkdiv_cry_12),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_13_LC_1_14_5.C_ON=1'b1;
    defparam clkdiv_13_LC_1_14_5.SEQ_MODE=4'b1000;
    defparam clkdiv_13_LC_1_14_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_13_LC_1_14_5 (
            .in0(_gnd_net_),
            .in1(N__6218),
            .in2(_gnd_net_),
            .in3(N__6212),
            .lcout(clkdivZ0Z_13),
            .ltout(),
            .carryin(clkdiv_cry_12),
            .carryout(clkdiv_cry_13),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_14_LC_1_14_6.C_ON=1'b1;
    defparam clkdiv_14_LC_1_14_6.SEQ_MODE=4'b1000;
    defparam clkdiv_14_LC_1_14_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_14_LC_1_14_6 (
            .in0(_gnd_net_),
            .in1(N__6209),
            .in2(_gnd_net_),
            .in3(N__6203),
            .lcout(clkdivZ0Z_14),
            .ltout(),
            .carryin(clkdiv_cry_13),
            .carryout(clkdiv_cry_14),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_15_LC_1_14_7.C_ON=1'b1;
    defparam clkdiv_15_LC_1_14_7.SEQ_MODE=4'b1000;
    defparam clkdiv_15_LC_1_14_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_15_LC_1_14_7 (
            .in0(_gnd_net_),
            .in1(N__6200),
            .in2(_gnd_net_),
            .in3(N__6194),
            .lcout(clkdivZ0Z_15),
            .ltout(),
            .carryin(clkdiv_cry_14),
            .carryout(clkdiv_cry_15),
            .clk(N__16123),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_16_LC_1_15_0.C_ON=1'b1;
    defparam clkdiv_16_LC_1_15_0.SEQ_MODE=4'b1000;
    defparam clkdiv_16_LC_1_15_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_16_LC_1_15_0 (
            .in0(_gnd_net_),
            .in1(N__6191),
            .in2(_gnd_net_),
            .in3(N__6185),
            .lcout(clkdivZ0Z_16),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(clkdiv_cry_16),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_17_LC_1_15_1.C_ON=1'b1;
    defparam clkdiv_17_LC_1_15_1.SEQ_MODE=4'b1000;
    defparam clkdiv_17_LC_1_15_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_17_LC_1_15_1 (
            .in0(_gnd_net_),
            .in1(N__6338),
            .in2(_gnd_net_),
            .in3(N__6332),
            .lcout(clkdivZ0Z_17),
            .ltout(),
            .carryin(clkdiv_cry_16),
            .carryout(clkdiv_cry_17),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_18_LC_1_15_2.C_ON=1'b1;
    defparam clkdiv_18_LC_1_15_2.SEQ_MODE=4'b1000;
    defparam clkdiv_18_LC_1_15_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_18_LC_1_15_2 (
            .in0(_gnd_net_),
            .in1(N__6329),
            .in2(_gnd_net_),
            .in3(N__6323),
            .lcout(clkdivZ0Z_18),
            .ltout(),
            .carryin(clkdiv_cry_17),
            .carryout(clkdiv_cry_18),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_19_LC_1_15_3.C_ON=1'b1;
    defparam clkdiv_19_LC_1_15_3.SEQ_MODE=4'b1000;
    defparam clkdiv_19_LC_1_15_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_19_LC_1_15_3 (
            .in0(_gnd_net_),
            .in1(N__6320),
            .in2(_gnd_net_),
            .in3(N__6314),
            .lcout(clkdivZ0Z_19),
            .ltout(),
            .carryin(clkdiv_cry_18),
            .carryout(clkdiv_cry_19),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_20_LC_1_15_4.C_ON=1'b1;
    defparam clkdiv_20_LC_1_15_4.SEQ_MODE=4'b1000;
    defparam clkdiv_20_LC_1_15_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_20_LC_1_15_4 (
            .in0(_gnd_net_),
            .in1(N__6311),
            .in2(_gnd_net_),
            .in3(N__6305),
            .lcout(clkdivZ0Z_20),
            .ltout(),
            .carryin(clkdiv_cry_19),
            .carryout(clkdiv_cry_20),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_21_LC_1_15_5.C_ON=1'b1;
    defparam clkdiv_21_LC_1_15_5.SEQ_MODE=4'b1000;
    defparam clkdiv_21_LC_1_15_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_21_LC_1_15_5 (
            .in0(_gnd_net_),
            .in1(N__6302),
            .in2(_gnd_net_),
            .in3(N__6296),
            .lcout(clkdivZ0Z_21),
            .ltout(),
            .carryin(clkdiv_cry_20),
            .carryout(clkdiv_cry_21),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_22_LC_1_15_6.C_ON=1'b1;
    defparam clkdiv_22_LC_1_15_6.SEQ_MODE=4'b1000;
    defparam clkdiv_22_LC_1_15_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_22_LC_1_15_6 (
            .in0(_gnd_net_),
            .in1(N__6293),
            .in2(_gnd_net_),
            .in3(N__6287),
            .lcout(clkdivZ0Z_22),
            .ltout(),
            .carryin(clkdiv_cry_21),
            .carryout(clkdiv_cry_22),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_23_LC_1_15_7.C_ON=1'b0;
    defparam clkdiv_23_LC_1_15_7.SEQ_MODE=4'b1000;
    defparam clkdiv_23_LC_1_15_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 clkdiv_23_LC_1_15_7 (
            .in0(_gnd_net_),
            .in1(N__6274),
            .in2(_gnd_net_),
            .in3(N__6284),
            .lcout(GPIO3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16124),
            .ce(),
            .sr(_gnd_net_));
    defparam a_14_LC_9_10_1.C_ON=1'b0;
    defparam a_14_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam a_14_LC_9_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_14_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14318),
            .lcout(aZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16108),
            .ce(N__12244),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_LC_9_10_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_LC_9_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_LC_9_10_2  (
            .in0(N__7282),
            .in1(N__7945),
            .in2(N__13783),
            .in3(N__12025),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_8_LC_9_10_5 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_8_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_8_LC_9_10_5 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.overflow_RNO_8_LC_9_10_5  (
            .in0(N__12026),
            .in1(N__7281),
            .in2(N__7962),
            .in3(N__11833),
            .lcout(\ALU.regsA_result_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_15_LC_9_10_6.C_ON=1'b0;
    defparam a_15_LC_9_10_6.SEQ_MODE=4'b1000;
    defparam a_15_LC_9_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_15_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12119),
            .lcout(aZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16108),
            .ce(N__12244),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_LC_9_11_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_LC_9_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__6590),
            .in2(N__6362),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\ALU.regsA_result_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_1_THRU_LUT4_0_LC_9_11_1 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_1_THRU_LUT4_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_1_THRU_LUT4_0_LC_9_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_1_THRU_LUT4_0_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6353),
            .lcout(\ALU.regsA_result_cry_1_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_LC_9_12_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_LC_9_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__6377),
            .in2(N__6796),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\ALU.regsA_result_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNIA939H_LC_9_12_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNIA939H_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNIA939H_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNIA939H_LC_9_12_1  (
            .in0(N__8255),
            .in1(N__6605),
            .in2(N__6506),
            .in3(N__6350),
            .lcout(\ALU.regsA_result_cry_4_c_RNIA939H ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4 ),
            .carryout(\ALU.regsA_result_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_5_c_RNIKCNNP_LC_9_12_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_5_c_RNIKCNNP_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_5_c_RNIKCNNP_LC_9_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_5_c_RNIKCNNP_LC_9_12_2  (
            .in0(N__8609),
            .in1(N__6371),
            .in2(N__6488),
            .in3(N__6347),
            .lcout(\ALU.regsA_result_cry_5_c_RNIKCNNP ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5 ),
            .carryout(\ALU.regsA_result_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_6_c_RNICICNO_LC_9_12_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_6_c_RNICICNO_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_6_c_RNICICNO_LC_9_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_6_c_RNICICNO_LC_9_12_3  (
            .in0(N__8585),
            .in1(N__6637),
            .in2(N__6626),
            .in3(N__6344),
            .lcout(\ALU.regsA_result_cry_6_c_RNICICNO ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6 ),
            .carryout(\ALU.regsA_result_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_7_THRU_LUT4_0_LC_9_12_4 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_7_THRU_LUT4_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_7_THRU_LUT4_0_LC_9_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_7_THRU_LUT4_0_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6341),
            .lcout(\ALU.regsA_result_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNO_LC_9_12_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNO_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNO_LC_9_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNO_LC_9_12_5  (
            .in0(N__7361),
            .in1(N__6792),
            .in2(_gnd_net_),
            .in3(N__13724),
            .lcout(\ALU.regsA_result_cry_4_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNIKGQO9_LC_9_12_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNIKGQO9_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNIKGQO9_LC_9_12_6 .LUT_INIT=16'b0110110001101100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNIKGQO9_LC_9_12_6  (
            .in0(N__13725),
            .in1(N__6565),
            .in2(N__7976),
            .in3(N__6487),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNIKGQO9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNO_LC_9_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNO_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNO_LC_9_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNO_LC_9_12_7  (
            .in0(N__6566),
            .in1(N__7963),
            .in2(_gnd_net_),
            .in3(N__13723),
            .lcout(\ALU.regsA_result_cry_2_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_12_LC_9_13_1.C_ON=1'b0;
    defparam a_12_LC_9_13_1.SEQ_MODE=4'b1000;
    defparam a_12_LC_9_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_12_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10970),
            .lcout(aZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16116),
            .ce(N__12242),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_LC_9_13_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_LC_9_13_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_LC_9_13_2  (
            .in0(N__13782),
            .in1(N__14660),
            .in2(N__12067),
            .in3(N__7353),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_2_l_ofx_LC_9_13_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_2_l_ofx_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_2_l_ofx_LC_9_13_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_2_l_ofx_LC_9_13_3  (
            .in0(N__12057),
            .in1(N__14659),
            .in2(N__7372),
            .in3(N__11831),
            .lcout(\ALU.regsA_result_axb_2_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_0_LC_9_15_1 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_0_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_0_LC_9_15_1 .LUT_INIT=16'b0111111100001111;
    LogicCell40 \FTDI.TXstate_RNO_0_0_LC_9_15_1  (
            .in0(N__14020),
            .in1(N__6770),
            .in2(N__15388),
            .in3(N__6727),
            .lcout(),
            .ltout(\FTDI.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_0_LC_9_15_2 .C_ON=1'b0;
    defparam \FTDI.TXstate_0_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_0_LC_9_15_2 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \FTDI.TXstate_0_LC_9_15_2  (
            .in0(N__6728),
            .in1(_gnd_net_),
            .in2(N__6365),
            .in3(N__12745),
            .lcout(\FTDI.TXstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_fast_3_LC_9_15_4 .C_ON=1'b0;
    defparam \FTDI.TXstate_fast_3_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_fast_3_LC_9_15_4 .LUT_INIT=16'b0111111100000100;
    LogicCell40 \FTDI.TXstate_fast_3_LC_9_15_4  (
            .in0(N__6731),
            .in1(N__6386),
            .in2(N__6776),
            .in3(N__6745),
            .lcout(\FTDI.TXstate_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNIE1MM_2_LC_9_15_5 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNIE1MM_2_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNIE1MM_2_LC_9_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FTDI.TXstate_RNIE1MM_2_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__12741),
            .in2(_gnd_net_),
            .in3(N__14019),
            .lcout(\FTDI.TXstate_RNIE1MMZ0Z_2 ),
            .ltout(\FTDI.TXstate_RNIE1MMZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_3_LC_9_15_6 .C_ON=1'b0;
    defparam \FTDI.TXstate_3_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_3_LC_9_15_6 .LUT_INIT=16'b0111111100010000;
    LogicCell40 \FTDI.TXstate_3_LC_9_15_6  (
            .in0(N__6730),
            .in1(N__6775),
            .in2(N__6380),
            .in3(N__15377),
            .lcout(\FTDI.TXstateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_1_LC_9_15_7 .C_ON=1'b0;
    defparam \FTDI.TXstate_1_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_1_LC_9_15_7 .LUT_INIT=16'b0110010011000100;
    LogicCell40 \FTDI.TXstate_1_LC_9_15_7  (
            .in0(N__12744),
            .in1(N__6771),
            .in2(N__15389),
            .in3(N__6729),
            .lcout(\FTDI.TXstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_15_l_ofx_LC_9_16_2 .C_ON=1'b0;
    defparam \ALU.addsub_axb_15_l_ofx_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_15_l_ofx_LC_9_16_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ALU.addsub_axb_15_l_ofx_LC_9_16_2  (
            .in0(N__14464),
            .in1(N__8180),
            .in2(_gnd_net_),
            .in3(N__7294),
            .lcout(\ALU.addsub_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_0_LC_9_17_3.C_ON=1'b0;
    defparam TXbuffer_RNO_0_0_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_0_LC_9_17_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 TXbuffer_RNO_0_0_LC_9_17_3 (
            .in0(N__7583),
            .in1(N__7546),
            .in2(_gnd_net_),
            .in3(N__15914),
            .lcout(N_91),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_1_LC_10_9_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_1_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_1_LC_10_9_0 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_1_LC_10_9_0  (
            .in0(N__8697),
            .in1(N__13768),
            .in2(N__6980),
            .in3(N__12062),
            .lcout(\ALU.mult_AdderTree2_bigtree_704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_LC_10_9_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_LC_10_9_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_LC_10_9_2  (
            .in0(N__8698),
            .in1(N__13769),
            .in2(N__12066),
            .in3(N__6976),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_11_LC_10_9_3.C_ON=1'b0;
    defparam a_11_LC_10_9_3.SEQ_MODE=4'b1000;
    defparam a_11_LC_10_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_11_LC_10_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10427),
            .lcout(aZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16099),
            .ce(N__12241),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_0_LC_10_9_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_0_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_0_LC_10_9_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_0_LC_10_9_4  (
            .in0(N__8691),
            .in1(N__13767),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_ma_LC_10_9_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_ma_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_ma_LC_10_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_ma_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__8692),
            .in2(_gnd_net_),
            .in3(N__12053),
            .lcout(\ALU.regsA_result_cry_2_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_ma_LC_10_9_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_ma_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_ma_LC_10_9_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_ma_LC_10_9_6  (
            .in0(N__11824),
            .in1(_gnd_net_),
            .in2(N__8719),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_3_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_ma_LC_10_9_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_ma_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_ma_LC_10_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_ma_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__8696),
            .in2(_gnd_net_),
            .in3(N__13344),
            .lcout(\ALU.regsA_result_cry_4_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_LC_10_10_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_LC_10_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__6449),
            .in2(N__6443),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\ALU.regsA_result_cry_1_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNI2J0N2_LC_10_10_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNI2J0N2_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNI2J0N2_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNI2J0N2_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__6434),
            .in2(N__6965),
            .in3(N__6425),
            .lcout(\ALU.mult_AdderTree2_bigtree_705 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_5 ),
            .carryout(\ALU.regsA_result_cry_2_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_0_c_RNI6Q6R2_LC_10_10_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_0_c_RNI6Q6R2_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_0_c_RNI6Q6R2_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_0_c_RNI6Q6R2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__6422),
            .in2(N__6956),
            .in3(N__6413),
            .lcout(\ALU.mult_AdderTree2_bigtree_706 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_7 ),
            .carryout(\ALU.regsA_result_cry_3_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_0_c_RNIA1DV2_LC_10_10_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_0_c_RNIA1DV2_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_0_c_RNIA1DV2_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_0_c_RNIA1DV2_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__6410),
            .in2(N__6395),
            .in3(N__6404),
            .lcout(\ALU.mult_AdderTree2_bigtree_707 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_7 ),
            .carryout(\ALU.regsA_result_cry_4_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_0_c_RNIE8JJ2_LC_10_10_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_0_c_RNIE8JJ2_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_0_c_RNIE8JJ2_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_0_c_RNIE8JJ2_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__6542),
            .in2(N__6947),
            .in3(N__6401),
            .lcout(\ALU.mult_AdderTree2_bigtree_708 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_6 ),
            .carryout(\ALU.regsA_result_cry_5_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_5_0_THRU_LUT4_0_LC_10_10_5 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_5_0_THRU_LUT4_0_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_5_0_THRU_LUT4_0_LC_10_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_5_0_THRU_LUT4_0_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6398),
            .lcout(\ALU.regsA_result_cry_5_0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_4_l_ofx_LC_10_10_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_4_l_ofx_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_4_l_ofx_LC_10_10_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_4_l_ofx_LC_10_10_6  (
            .in0(N__11657),
            .in1(N__8723),
            .in2(N__7445),
            .in3(N__13317),
            .lcout(\ALU.regsA_result_axb_4_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_5_ma_LC_10_10_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_5_ma_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_5_ma_LC_10_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_5_ma_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__11658),
            .in2(_gnd_net_),
            .in3(N__8699),
            .lcout(\ALU.regsA_result_cry_5_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_LC_10_11_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_LC_10_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__7082),
            .in2(N__7105),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\ALU.regsA_result_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNIHNOEF_LC_10_11_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNIHNOEF_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNIHNOEF_LC_10_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNIHNOEF_LC_10_11_1  (
            .in0(N__8318),
            .in1(N__6536),
            .in2(N__7037),
            .in3(N__6527),
            .lcout(\ALU.regsA_result_cry_2_c_RNIHNOEF ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_0 ),
            .carryout(\ALU.regsA_result_cry_3_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_3_c_RNIHID36_LC_10_11_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_3_c_RNIHID36_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_3_c_RNIHID36_LC_10_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_3_c_RNIHID36_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__6524),
            .in2(N__7016),
            .in3(N__6518),
            .lcout(\ALU.mult_AdderTree2_bigtree_870 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_4 ),
            .carryout(\ALU.regsA_result_cry_4_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_4_c_RNIQ2RR5_LC_10_11_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_4_c_RNIQ2RR5_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_4_c_RNIQ2RR5_LC_10_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_4_c_RNIQ2RR5_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__6515),
            .in2(N__6995),
            .in3(N__6497),
            .lcout(\ALU.mult_AdderTree2_bigtree_871 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_3 ),
            .carryout(\ALU.regsA_result_cry_5_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_5_c_RNI3J846_LC_10_11_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_5_c_RNI3J846_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_5_c_RNI3J846_LC_10_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_5_c_RNI3J846_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__6494),
            .in2(N__7157),
            .in3(N__6473),
            .lcout(\ALU.mult_AdderTree2_bigtree_872 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_4 ),
            .carryout(\ALU.regsA_result_cry_6_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_6_c_RNIC3MS5_LC_10_11_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_6_c_RNIC3MS5_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_6_c_RNIC3MS5_LC_10_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_6_c_RNIC3MS5_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__7145),
            .in2(N__6470),
            .in3(N__6461),
            .lcout(\ALU.mult_AdderTree2_bigtree_873 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_3 ),
            .carryout(\ALU.regsA_result_cry_7_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_2_LC_10_11_6 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_2_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_2_LC_10_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_2_LC_10_11_6  (
            .in0(N__6611),
            .in1(N__6665),
            .in2(N__7127),
            .in3(N__6458),
            .lcout(\ALU.regsA_result_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_LC_10_12_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_LC_10_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__6455),
            .in2(N__6564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\ALU.regsA_result_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNIC59KA_LC_10_12_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNIC59KA_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNIC59KA_LC_10_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNIC59KA_LC_10_12_1  (
            .in0(N__6638),
            .in1(N__6698),
            .in2(N__6599),
            .in3(N__6617),
            .lcout(\ALU.regsA_result_cry_2_c_RNIC59KA ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2 ),
            .carryout(\ALU.regsA_result_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_3_0_THRU_LUT4_0_LC_10_12_2 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_3_0_THRU_LUT4_0_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_3_0_THRU_LUT4_0_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_3_0_THRU_LUT4_0_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6614),
            .lcout(\ALU.regsA_result_cry_3_0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_1_LC_10_12_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_1_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_1_LC_10_12_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_1_LC_10_12_3  (
            .in0(N__12064),
            .in1(N__7362),
            .in2(N__13766),
            .in3(N__14648),
            .lcout(\ALU.mult_AdderTree2_bigtree_739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_axb_1_LC_10_12_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_axb_1_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_axb_1_LC_10_12_4 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_axb_1_LC_10_12_4  (
            .in0(N__7290),
            .in1(N__13717),
            .in2(N__7977),
            .in3(N__12063),
            .lcout(\ALU.mult_AdderTree2_bigtree_774 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_0_LC_10_12_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_0_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_0_LC_10_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_0_LC_10_12_6  (
            .in0(N__7289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13716),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_5_l_ofx_LC_10_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_5_l_ofx_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_5_l_ofx_LC_10_12_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_5_l_ofx_LC_10_12_7  (
            .in0(N__7788),
            .in1(N__11661),
            .in2(N__15041),
            .in3(N__7881),
            .lcout(\ALU.regsA_result_axb_5_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_LC_10_13_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_LC_10_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__7175),
            .in2(N__6584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\ALU.regsA_result_cry_1_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNI9GUP2_LC_10_13_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNI9GUP2_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNI9GUP2_LC_10_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNI9GUP2_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__11138),
            .in2(N__6575),
            .in3(N__6545),
            .lcout(\ALU.mult_AdderTree2_bigtree_740 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_4 ),
            .carryout(\ALU.regsA_result_cry_2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_0_c_RNIDN4U2_LC_10_13_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_0_c_RNIDN4U2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_0_c_RNIDN4U2_LC_10_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_0_c_RNIDN4U2_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__7073),
            .in2(N__6656),
            .in3(N__6692),
            .lcout(\ALU.mult_AdderTree2_bigtree_741 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_6 ),
            .carryout(\ALU.regsA_result_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_4_LC_10_13_3 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_4_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_4_LC_10_13_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_4_LC_10_13_3  (
            .in0(N__6689),
            .in1(N__6677),
            .in2(N__6647),
            .in3(N__6668),
            .lcout(\ALU.regsA_result_axb_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_3_l_ofx_LC_10_13_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_3_l_ofx_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_3_l_ofx_LC_10_13_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_3_l_ofx_LC_10_13_4  (
            .in0(N__13342),
            .in1(N__7357),
            .in2(N__11834),
            .in3(N__14656),
            .lcout(\ALU.regsA_result_axb_3_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_9_LC_10_13_5 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_9_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_9_LC_10_13_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.overflow_RNO_9_LC_10_13_5  (
            .in0(N__14655),
            .in1(N__11659),
            .in2(N__7373),
            .in3(N__13343),
            .lcout(\ALU.regsA_result_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_FirstStep_AB_1_128_LC_10_13_7 .C_ON=1'b0;
    defparam \ALU.mult_FirstStep_AB_1_128_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_FirstStep_AB_1_128_LC_10_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_FirstStep_AB_1_128_LC_10_13_7  (
            .in0(N__13772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7896),
            .lcout(\ALU.mult_ab_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_2_l_ofx_LC_10_14_0 .C_ON=1'b0;
    defparam \ALU.addsub_axb_2_l_ofx_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_2_l_ofx_LC_10_14_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ALU.addsub_axb_2_l_ofx_LC_10_14_0  (
            .in0(N__14446),
            .in1(N__11832),
            .in2(_gnd_net_),
            .in3(N__9803),
            .lcout(\ALU.addsub_axb_2_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_0_LC_10_14_1 .C_ON=1'b0;
    defparam \FTDI.baudAcc_0_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_0_LC_10_14_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \FTDI.baudAcc_0_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__6825),
            .in2(_gnd_net_),
            .in3(N__16173),
            .lcout(\FTDI.baudAccZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_1_LC_10_14_2 .C_ON=1'b0;
    defparam \FTDI.baudAcc_1_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_1_LC_10_14_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \FTDI.baudAcc_1_LC_10_14_2  (
            .in0(N__16174),
            .in1(_gnd_net_),
            .in2(N__6832),
            .in3(N__6814),
            .lcout(\FTDI.baudAccZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_10_l_ofx_LC_10_14_4 .C_ON=1'b0;
    defparam \ALU.addsub_axb_10_l_ofx_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_10_l_ofx_LC_10_14_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.addsub_axb_10_l_ofx_LC_10_14_4  (
            .in0(N__14447),
            .in1(_gnd_net_),
            .in2(N__7451),
            .in3(N__14161),
            .lcout(\ALU.addsub_axb_10_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_1_LC_10_14_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_1_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_1_LC_10_14_5 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_1_LC_10_14_5  (
            .in0(N__7789),
            .in1(N__13771),
            .in2(N__7907),
            .in3(N__12048),
            .lcout(\ALU.mult_AdderTree2_bigtree_669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_2_LC_10_14_6 .C_ON=1'b0;
    defparam \FTDI.baudAcc_2_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_2_LC_10_14_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \FTDI.baudAcc_2_LC_10_14_6  (
            .in0(N__16175),
            .in1(_gnd_net_),
            .in2(N__6833),
            .in3(N__6815),
            .lcout(\FTDI.baudAccZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNI073QE_LC_10_14_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNI073QE_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNI073QE_LC_10_14_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNI073QE_LC_10_14_7  (
            .in0(N__7109),
            .in1(N__7446),
            .in2(N__8351),
            .in3(N__13770),
            .lcout(\ALU.regsA_result_cry_5_c_RNI073QE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_1_2_LC_10_15_0 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_1_2_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_1_2_LC_10_15_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \FTDI.TXstate_RNO_1_2_LC_10_15_0  (
            .in0(N__12742),
            .in1(N__6769),
            .in2(_gnd_net_),
            .in3(N__6726),
            .lcout(),
            .ltout(\FTDI.N_170_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_2_LC_10_15_1 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_2_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_2_LC_10_15_1 .LUT_INIT=16'b1100010001011111;
    LogicCell40 \FTDI.TXstate_RNO_0_2_LC_10_15_1  (
            .in0(N__15381),
            .in1(N__12743),
            .in2(N__6803),
            .in3(N__14018),
            .lcout(),
            .ltout(\FTDI.TXstate_cnst_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_2_LC_10_15_2 .C_ON=1'b0;
    defparam \FTDI.TXstate_2_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_2_LC_10_15_2 .LUT_INIT=16'b1100111100001111;
    LogicCell40 \FTDI.TXstate_2_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__12689),
            .in2(N__6800),
            .in3(N__16172),
            .lcout(\FTDI.un3_TX_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNI8EG3H_LC_10_15_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNI8EG3H_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNI8EG3H_LC_10_15_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNI8EG3H_LC_10_15_3  (
            .in0(N__7374),
            .in1(N__13780),
            .in2(N__8285),
            .in3(N__6797),
            .lcout(\ALU.regsA_result_cry_7_c_RNI8EG3H ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_fast_RNIRJI91_3_LC_10_15_4 .C_ON=1'b0;
    defparam \FTDI.TXstate_fast_RNIRJI91_3_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_fast_RNIRJI91_3_LC_10_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \FTDI.TXstate_fast_RNIRJI91_3_LC_10_15_4  (
            .in0(N__14017),
            .in1(N__6768),
            .in2(N__6746),
            .in3(N__6725),
            .lcout(FTDI_TXready),
            .ltout(FTDI_TXready_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXstart_esr_RNO_0_LC_10_15_5.C_ON=1'b0;
    defparam TXstart_esr_RNO_0_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam TXstart_esr_RNO_0_LC_10_15_5.LUT_INIT=16'b1010100010001000;
    LogicCell40 TXstart_esr_RNO_0_LC_10_15_5 (
            .in0(N__15778),
            .in1(N__15661),
            .in2(N__6704),
            .in3(N__15902),
            .lcout(),
            .ltout(un1_testState31_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXstart_esr_RNO_LC_10_15_6.C_ON=1'b0;
    defparam TXstart_esr_RNO_LC_10_15_6.SEQ_MODE=4'b0000;
    defparam TXstart_esr_RNO_LC_10_15_6.LUT_INIT=16'b1111101011111010;
    LogicCell40 TXstart_esr_RNO_LC_10_15_6 (
            .in0(N__15947),
            .in1(_gnd_net_),
            .in2(N__6701),
            .in3(_gnd_net_),
            .lcout(un1_testState31_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_4_m1_forloop_1_1_regsA_result_cry_0_c_LC_10_16_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_4_m1_forloop_1_1_regsA_result_cry_0_c_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_4_m1_forloop_1_1_regsA_result_cry_0_c_LC_10_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_4_m1_forloop_1_1_regsA_result_cry_0_c_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__7613),
            .in2(N__8393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\ALU.regsA_result_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_9_LC_10_16_1 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_9_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_9_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_9_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__6935),
            .in2(N__8369),
            .in3(N__6926),
            .lcout(\ALU.mult_9 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_0_0 ),
            .carryout(\ALU.regsA_result_cry_1_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_10_LC_10_16_2 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_10_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_10_LC_10_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_10_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__6923),
            .in2(N__8350),
            .in3(N__6911),
            .lcout(\ALU.mult_10 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_1 ),
            .carryout(\ALU.regsA_result_cry_2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_11_LC_10_16_3 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_11_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_11_LC_10_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_11_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__6908),
            .in2(N__8317),
            .in3(N__6899),
            .lcout(\ALU.mult_11 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_2 ),
            .carryout(\ALU.regsA_result_cry_3_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_12_LC_10_16_4 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_12_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_12_LC_10_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_12_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__6896),
            .in2(N__8281),
            .in3(N__6890),
            .lcout(\ALU.mult_12 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_2 ),
            .carryout(\ALU.regsA_result_cry_4_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_13_LC_10_16_5 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_13_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_13_LC_10_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_13_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__8254),
            .in2(N__6887),
            .in3(N__6872),
            .lcout(\ALU.mult_13 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_1 ),
            .carryout(\ALU.regsA_result_cry_5_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_14_LC_10_16_6 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_14_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_14_LC_10_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_14_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__8602),
            .in2(N__6869),
            .in3(N__6854),
            .lcout(\ALU.mult_14 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_2 ),
            .carryout(\ALU.regsA_result_cry_6_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_15_LC_10_16_7 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_15_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_15_LC_10_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_15_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__8581),
            .in2(N__6851),
            .in3(N__6836),
            .lcout(\ALU.mult_15 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_1 ),
            .carryout(\ALU.regsA_result_cry_7_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_0_LC_10_17_0 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_0_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_0_LC_10_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.overflow_RNO_0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__8525),
            .in2(_gnd_net_),
            .in3(N__6983),
            .lcout(\ALU.mult_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_30_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_30_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_30_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_fast_10_LC_11_8_5.C_ON=1'b0;
    defparam a_fast_10_LC_11_8_5.SEQ_MODE=4'b1000;
    defparam a_fast_10_LC_11_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_fast_10_LC_11_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11095),
            .lcout(a_fastZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16088),
            .ce(N__12245),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_2_l_ofx_LC_11_9_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_2_l_ofx_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_2_l_ofx_LC_11_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_2_l_ofx_LC_11_9_0  (
            .in0(N__12065),
            .in1(N__11825),
            .in2(N__8743),
            .in3(N__7419),
            .lcout(\ALU.regsA_result_axb_2_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_10_LC_11_9_1.C_ON=1'b0;
    defparam a_10_LC_11_9_1.SEQ_MODE=4'b1000;
    defparam a_10_LC_11_9_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_10_LC_11_9_1 (
            .in0(N__11106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16094),
            .ce(N__12199),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_3_l_ofx_LC_11_9_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_3_l_ofx_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_3_l_ofx_LC_11_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_3_l_ofx_LC_11_9_2  (
            .in0(N__13334),
            .in1(N__11826),
            .in2(N__8744),
            .in3(N__7420),
            .lcout(\ALU.regsA_result_axb_3_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_5_l_ofx_LC_11_9_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_5_l_ofx_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_5_l_ofx_LC_11_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_5_l_ofx_LC_11_9_4  (
            .in0(N__11611),
            .in1(N__7421),
            .in2(N__8745),
            .in3(N__15039),
            .lcout(\ALU.regsA_result_axb_5_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_8_LC_11_10_1.C_ON=1'b0;
    defparam a_8_LC_11_10_1.SEQ_MODE=4'b1000;
    defparam a_8_LC_11_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_8_LC_11_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14514),
            .lcout(aZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16100),
            .ce(N__12243),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_LC_11_10_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_LC_11_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_LC_11_10_2  (
            .in0(N__7763),
            .in1(N__13744),
            .in2(N__12061),
            .in3(N__7851),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_2_l_ofx_LC_11_10_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_2_l_ofx_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_2_l_ofx_LC_11_10_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_2_l_ofx_LC_11_10_3  (
            .in0(N__12034),
            .in1(N__7759),
            .in2(N__7878),
            .in3(N__11785),
            .lcout(\ALU.regsA_result_axb_2_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_3_l_ofx_LC_11_10_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_3_l_ofx_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_3_l_ofx_LC_11_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_3_l_ofx_LC_11_10_4  (
            .in0(N__7760),
            .in1(N__13315),
            .in2(N__11814),
            .in3(N__7855),
            .lcout(\ALU.regsA_result_axb_3_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_4_l_ofx_LC_11_10_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_4_l_ofx_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_4_l_ofx_LC_11_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_4_l_ofx_LC_11_10_5  (
            .in0(N__13316),
            .in1(N__7761),
            .in2(N__7879),
            .in3(N__11602),
            .lcout(\ALU.regsA_result_axb_4_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_6_l_ofx_LC_11_10_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_6_l_ofx_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_6_l_ofx_LC_11_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_6_l_ofx_LC_11_10_7  (
            .in0(N__15040),
            .in1(N__7762),
            .in2(N__7880),
            .in3(N__13081),
            .lcout(\ALU.regsA_result_axb_6_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_LC_11_11_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__8024),
            .in2(N__7067),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\ALU.regsA_result_cry_1_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNI6MAO2_LC_11_11_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNI6MAO2_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNI6MAO2_LC_11_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNI6MAO2_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__8015),
            .in2(N__7058),
            .in3(N__7049),
            .lcout(\ALU.mult_AdderTree2_bigtree_670 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_6 ),
            .carryout(\ALU.regsA_result_cry_2_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_0_c_RNIATGS2_LC_11_11_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_0_c_RNIATGS2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_0_c_RNIATGS2_LC_11_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_0_c_RNIATGS2_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__8003),
            .in2(N__7046),
            .in3(N__7028),
            .lcout(\ALU.mult_AdderTree2_bigtree_671 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_8 ),
            .carryout(\ALU.regsA_result_cry_3_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_0_c_RNIE4N03_LC_11_11_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_0_c_RNIE4N03_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_0_c_RNIE4N03_LC_11_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_0_c_RNIE4N03_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__7994),
            .in2(N__7025),
            .in3(N__7007),
            .lcout(\ALU.mult_AdderTree2_bigtree_672 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_8 ),
            .carryout(\ALU.regsA_result_cry_4_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_0_c_RNIIBTK2_LC_11_11_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_0_c_RNIIBTK2_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_0_c_RNIIBTK2_LC_11_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_0_c_RNIIBTK2_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__7004),
            .in2(N__7688),
            .in3(N__6986),
            .lcout(\ALU.mult_AdderTree2_bigtree_673 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_7 ),
            .carryout(\ALU.regsA_result_cry_5_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_0_c_RNIMI3P2_LC_11_11_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_0_c_RNIMI3P2_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_0_c_RNIMI3P2_LC_11_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_0_c_RNIMI3P2_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__7118),
            .in2(N__7166),
            .in3(N__7148),
            .lcout(\ALU.mult_AdderTree2_bigtree_674 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_7 ),
            .carryout(\ALU.regsA_result_cry_6_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_0_c_RNIQP9T2_LC_11_11_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_0_c_RNIQP9T2_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_0_c_RNIQP9T2_LC_11_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_0_c_RNIQP9T2_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__7640),
            .in2(N__7631),
            .in3(N__7139),
            .lcout(\ALU.mult_AdderTree2_bigtree_675 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_6 ),
            .carryout(\ALU.regsA_result_cry_7_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_5_LC_11_11_7 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_5_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_5_LC_11_11_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_5_LC_11_11_7  (
            .in0(N__7136),
            .in1(N__7181),
            .in2(N__7622),
            .in3(N__7130),
            .lcout(\ALU.regsA_result_axb_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_7_l_ofx_LC_11_12_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_7_l_ofx_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_7_l_ofx_LC_11_12_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_7_l_ofx_LC_11_12_0  (
            .in0(N__14867),
            .in1(N__13183),
            .in2(N__12626),
            .in3(N__12844),
            .lcout(\ALU.regsA_result_axb_7_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_12_l_ofx_LC_11_12_1 .C_ON=1'b0;
    defparam \ALU.addsub_axb_12_l_ofx_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_12_l_ofx_LC_11_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_12_l_ofx_LC_11_12_1  (
            .in0(N__7382),
            .in1(N__14459),
            .in2(_gnd_net_),
            .in3(N__9599),
            .lcout(\ALU.addsub_axb_12_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_2_l_ofx_LC_11_12_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_2_l_ofx_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_2_l_ofx_LC_11_12_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_2_l_ofx_LC_11_12_2  (
            .in0(N__14866),
            .in1(N__13345),
            .in2(N__12625),
            .in3(N__11798),
            .lcout(\ALU.regsA_result_axb_2_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_ma_LC_11_12_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_ma_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_ma_LC_11_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_ma_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__7781),
            .in2(_gnd_net_),
            .in3(N__15031),
            .lcout(\ALU.regsA_result_cry_6_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNO_LC_11_12_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNO_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNO_LC_11_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNO_LC_11_12_4  (
            .in0(N__13722),
            .in1(N__7104),
            .in2(_gnd_net_),
            .in3(N__7435),
            .lcout(\ALU.regsA_result_cry_2_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_3_ma_LC_11_12_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_3_ma_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_3_ma_LC_11_12_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_3_ma_LC_11_12_5  (
            .in0(N__11799),
            .in1(_gnd_net_),
            .in2(N__14658),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_3_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_10_LC_11_12_6 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_10_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_10_LC_11_12_6 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.overflow_RNO_10_LC_11_12_6  (
            .in0(N__15032),
            .in1(N__7436),
            .in2(N__13091),
            .in3(N__8739),
            .lcout(\ALU.regsA_result_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_0_LC_11_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_0_LC_11_12_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_0_LC_11_12_7  (
            .in0(N__14644),
            .in1(N__13721),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_1_LC_11_13_1.C_ON=1'b0;
    defparam a_1_LC_11_13_1.SEQ_MODE=4'b1000;
    defparam a_1_LC_11_13_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_1_LC_11_13_1 (
            .in0(N__11336),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16109),
            .ce(N__15295),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_LC_11_13_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_LC_11_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_LC_11_13_2  (
            .in0(N__12036),
            .in1(N__13755),
            .in2(N__14898),
            .in3(N__12608),
            .lcout(\ALU.regsA_result_cry_0_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_1_l_ofx_LC_11_13_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_1_l_ofx_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_1_l_ofx_LC_11_13_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_1_l_ofx_LC_11_13_3  (
            .in0(N__14876),
            .in1(N__11827),
            .in2(N__12639),
            .in3(N__12035),
            .lcout(\ALU.regsA_result_axb_1_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_3_l_ofx_LC_11_13_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_3_l_ofx_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_3_l_ofx_LC_11_13_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_3_l_ofx_LC_11_13_5  (
            .in0(N__14877),
            .in1(N__11660),
            .in2(N__12640),
            .in3(N__13325),
            .lcout(\ALU.regsA_result_axb_3_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_4_l_ofx_LC_11_13_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_4_l_ofx_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_4_l_ofx_LC_11_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_4_l_ofx_LC_11_13_6  (
            .in0(N__15038),
            .in1(N__11606),
            .in2(N__14897),
            .in3(N__12615),
            .lcout(\ALU.regsA_result_axb_4_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_5_l_ofx_LC_11_13_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_5_l_ofx_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_5_l_ofx_LC_11_13_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_5_l_ofx_LC_11_13_7  (
            .in0(N__14878),
            .in1(N__13089),
            .in2(N__12641),
            .in3(N__15037),
            .lcout(\ALU.regsA_result_axb_5_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_0_c_THRU_CRY_0_LC_11_14_0 .C_ON=1'b1;
    defparam \ALU.addsub_cry_0_c_THRU_CRY_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_0_c_THRU_CRY_0_LC_11_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.addsub_cry_0_c_THRU_CRY_0_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__14448),
            .in2(N__14463),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\ALU.addsub_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_0_LC_11_14_1 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_0_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_0_LC_11_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_0_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__14889),
            .in2(N__8141),
            .in3(N__7169),
            .lcout(\ALU.addsub_0 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_0_c_THRU_CO ),
            .carryout(\ALU.addsub_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_1_LC_11_14_2 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_1_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_1_LC_11_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_1_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__12603),
            .in2(N__8189),
            .in3(N__7217),
            .lcout(\ALU.addsub_1 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_0 ),
            .carryout(\ALU.addsub_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_2_LC_11_14_3 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_2_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_2_LC_11_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_2_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__9802),
            .in2(N__7214),
            .in3(N__7205),
            .lcout(\ALU.addsub_2 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_1 ),
            .carryout(\ALU.addsub_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_3_LC_11_14_4 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_3_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_3_LC_11_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_3_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__13523),
            .in2(N__13196),
            .in3(N__7202),
            .lcout(\ALU.addsub_3 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_2 ),
            .carryout(\ALU.addsub_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_4_LC_11_14_5 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_4_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_4_LC_11_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_4_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__10901),
            .in2(N__10856),
            .in3(N__7199),
            .lcout(\ALU.addsub_4 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_3 ),
            .carryout(\ALU.addsub_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_5_LC_11_14_6 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_5_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_5_LC_11_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_5_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__15204),
            .in2(N__14918),
            .in3(N__7196),
            .lcout(\ALU.addsub_5 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_4 ),
            .carryout(\ALU.addsub_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_6_LC_11_14_7 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_6_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_6_LC_11_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_6_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__13879),
            .in2(N__13928),
            .in3(N__7193),
            .lcout(\ALU.addsub_6 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_5 ),
            .carryout(\ALU.addsub_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_7_LC_11_15_0 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_7_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_7_LC_11_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_7_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__12967),
            .in2(N__8222),
            .in3(N__7190),
            .lcout(\ALU.addsub_7 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\ALU.addsub_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_8_LC_11_15_1 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_8_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_8_LC_11_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_8_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__7906),
            .in2(N__7820),
            .in3(N__7187),
            .lcout(\ALU.addsub_8 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_7 ),
            .carryout(\ALU.addsub_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_9_LC_11_15_2 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_9_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_9_LC_11_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_9_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__7805),
            .in2(N__7793),
            .in3(N__7184),
            .lcout(\ALU.addsub_9 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_8 ),
            .carryout(\ALU.addsub_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_10_LC_11_15_3 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_10_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_10_LC_11_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_10_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__7450),
            .in2(N__7397),
            .in3(N__7388),
            .lcout(\ALU.addsub_10 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_9 ),
            .carryout(\ALU.addsub_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_11_LC_11_15_4 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_11_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_11_LC_11_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_11_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__8747),
            .in2(N__8651),
            .in3(N__7385),
            .lcout(\ALU.addsub_11 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_10 ),
            .carryout(\ALU.addsub_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_12_LC_11_15_5 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_12_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_12_LC_11_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_12_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__7381),
            .in2(N__7316),
            .in3(N__7304),
            .lcout(\ALU.addsub_12 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_11 ),
            .carryout(\ALU.addsub_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_13_LC_11_15_6 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_13_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_13_LC_11_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_13_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__14657),
            .in2(N__14534),
            .in3(N__7301),
            .lcout(\ALU.addsub_13 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_12 ),
            .carryout(\ALU.addsub_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_14_LC_11_15_7 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_14_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_14_LC_11_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_14_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__7984),
            .in2(N__7922),
            .in3(N__7298),
            .lcout(\ALU.addsub_14 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_13 ),
            .carryout(\ALU.addsub_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_0_15_LC_11_16_0 .C_ON=1'b1;
    defparam \ALU.res_RNO_0_15_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_0_15_LC_11_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_0_15_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__7295),
            .in2(N__7253),
            .in3(N__7241),
            .lcout(\ALU.addsub_15 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\ALU.addsub_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_LC_11_16_1 .C_ON=1'b0;
    defparam \ALU.overflow_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \ALU.overflow_LC_11_16_1 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \ALU.overflow_LC_11_16_1  (
            .in0(N__11271),
            .in1(N__7238),
            .in2(N__14465),
            .in3(N__7232),
            .lcout(overflow),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_1_LC_11_16_2 .C_ON=1'b0;
    defparam \ALU.res_RNO_1_1_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_1_LC_11_16_2 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.res_RNO_1_1_LC_11_16_2  (
            .in0(N__12049),
            .in1(N__12638),
            .in2(N__14899),
            .in3(N__13781),
            .lcout(\ALU.mult_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_14_LC_11_16_3 .C_ON=1'b0;
    defparam \ALU.res_14_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \ALU.res_14_LC_11_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_14_LC_11_16_3  (
            .in0(N__11276),
            .in1(N__7229),
            .in2(_gnd_net_),
            .in3(N__7223),
            .lcout(res_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_8_LC_11_16_4 .C_ON=1'b0;
    defparam \ALU.res_8_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \ALU.res_8_LC_11_16_4 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ALU.res_8_LC_11_16_4  (
            .in0(N__7612),
            .in1(N__11278),
            .in2(N__7592),
            .in3(N__8386),
            .lcout(res_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_11_LC_11_16_5 .C_ON=1'b0;
    defparam \ALU.res_11_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \ALU.res_11_LC_11_16_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_11_LC_11_16_5  (
            .in0(N__11272),
            .in1(N__7571),
            .in2(_gnd_net_),
            .in3(N__7565),
            .lcout(res_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_0_LC_11_16_6 .C_ON=1'b0;
    defparam \ALU.res_0_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \ALU.res_0_LC_11_16_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ALU.res_0_LC_11_16_6  (
            .in0(N__13784),
            .in1(N__7559),
            .in2(N__14900),
            .in3(N__11277),
            .lcout(GPIO0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_13_LC_11_16_7 .C_ON=1'b0;
    defparam \ALU.res_13_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \ALU.res_13_LC_11_16_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.res_13_LC_11_16_7  (
            .in0(N__7523),
            .in1(_gnd_net_),
            .in2(N__11285),
            .in3(N__7517),
            .lcout(res_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_12_LC_11_17_1 .C_ON=1'b0;
    defparam \ALU.res_12_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \ALU.res_12_LC_11_17_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_12_LC_11_17_1  (
            .in0(N__11280),
            .in1(N__7511),
            .in2(_gnd_net_),
            .in3(N__7502),
            .lcout(res_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16120),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_1_LC_11_17_2 .C_ON=1'b0;
    defparam \ALU.res_1_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \ALU.res_1_LC_11_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.res_1_LC_11_17_2  (
            .in0(N__11284),
            .in1(N__7496),
            .in2(_gnd_net_),
            .in3(N__7490),
            .lcout(GPIO1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16120),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_9_LC_11_17_3 .C_ON=1'b0;
    defparam \ALU.res_9_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \ALU.res_9_LC_11_17_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_9_LC_11_17_3  (
            .in0(N__11282),
            .in1(N__7481),
            .in2(_gnd_net_),
            .in3(N__7472),
            .lcout(res_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16120),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_10_LC_11_17_4 .C_ON=1'b0;
    defparam \ALU.res_10_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \ALU.res_10_LC_11_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_10_LC_11_17_4  (
            .in0(N__11283),
            .in1(N__7466),
            .in2(_gnd_net_),
            .in3(N__7457),
            .lcout(res_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16120),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_15_LC_11_17_7 .C_ON=1'b0;
    defparam \ALU.res_15_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \ALU.res_15_LC_11_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_15_LC_11_17_7  (
            .in0(N__11281),
            .in1(N__7679),
            .in2(_gnd_net_),
            .in3(N__7673),
            .lcout(res_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16120),
            .ce(),
            .sr(_gnd_net_));
    defparam b_15_LC_12_8_6.C_ON=1'b0;
    defparam b_15_LC_12_8_6.SEQ_MODE=4'b1000;
    defparam b_15_LC_12_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_15_LC_12_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12104),
            .lcout(bZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16083),
            .ce(N__14225),
            .sr(_gnd_net_));
    defparam \ALU.res_6_LC_12_9_0 .C_ON=1'b0;
    defparam \ALU.res_6_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \ALU.res_6_LC_12_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_6_LC_12_9_0  (
            .in0(N__11231),
            .in1(N__7667),
            .in2(_gnd_net_),
            .in3(N__8411),
            .lcout(res_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16089),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_2_LC_12_9_1 .C_ON=1'b0;
    defparam \ALU.res_RNO_1_2_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_2_LC_12_9_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALU.res_RNO_1_2_LC_12_9_1  (
            .in0(N__9801),
            .in1(N__9829),
            .in2(_gnd_net_),
            .in3(N__13765),
            .lcout(),
            .ltout(\ALU.mult_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_2_LC_12_9_2 .C_ON=1'b0;
    defparam \ALU.res_2_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \ALU.res_2_LC_12_9_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.res_2_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__11230),
            .in2(N__7655),
            .in3(N__7652),
            .lcout(GPIO2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16089),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_ma_LC_12_9_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_ma_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_ma_LC_12_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_ma_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__11610),
            .in2(_gnd_net_),
            .in3(N__13513),
            .lcout(\ALU.regsA_result_cry_5_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_7_ma_LC_12_9_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_7_ma_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_7_ma_LC_12_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_7_ma_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__7758),
            .in2(_gnd_net_),
            .in3(N__13085),
            .lcout(\ALU.regsA_result_cry_7_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_7_l_ofx_LC_12_10_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_7_l_ofx_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_7_l_ofx_LC_12_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_7_l_ofx_LC_12_10_0  (
            .in0(N__7748),
            .in1(N__12851),
            .in2(N__13090),
            .in3(N__7882),
            .lcout(\ALU.regsA_result_axb_7_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_11_LC_12_10_1 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_11_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_11_LC_12_10_1 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.overflow_RNO_11_LC_12_10_1  (
            .in0(N__12852),
            .in1(N__7747),
            .in2(N__7895),
            .in3(N__13178),
            .lcout(\ALU.regsA_result_axb_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_9_LC_12_10_2.C_ON=1'b0;
    defparam a_9_LC_12_10_2.SEQ_MODE=4'b1000;
    defparam a_9_LC_12_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_9_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11332),
            .lcout(aZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16095),
            .ce(N__12231),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_0_LC_12_10_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_0_LC_12_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__13728),
            .in2(_gnd_net_),
            .in3(N__7739),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_ma_LC_12_10_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_ma_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_ma_LC_12_10_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_ma_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7767),
            .in3(N__12033),
            .lcout(\ALU.regsA_result_cry_2_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_ma_LC_12_10_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_ma_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_ma_LC_12_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_ma_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__11784),
            .in2(_gnd_net_),
            .in3(N__7743),
            .lcout(\ALU.regsA_result_cry_3_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_ma_LC_12_10_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_ma_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_ma_LC_12_10_6 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_ma_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__13318),
            .in2(N__7768),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_4_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_14_l_ofx_LC_12_11_0 .C_ON=1'b0;
    defparam \ALU.addsub_axb_14_l_ofx_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_14_l_ofx_LC_12_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_14_l_ofx_LC_12_11_0  (
            .in0(N__7985),
            .in1(N__14267),
            .in2(_gnd_net_),
            .in3(N__14457),
            .lcout(\ALU.addsub_axb_14_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_8_l_ofx_LC_12_11_1 .C_ON=1'b0;
    defparam \ALU.addsub_axb_8_l_ofx_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_8_l_ofx_LC_12_11_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.addsub_axb_8_l_ofx_LC_12_11_1  (
            .in0(N__14455),
            .in1(N__7877),
            .in2(_gnd_net_),
            .in3(N__13182),
            .lcout(\ALU.addsub_axb_8_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_9_l_ofx_LC_12_11_4 .C_ON=1'b0;
    defparam \ALU.addsub_axb_9_l_ofx_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_9_l_ofx_LC_12_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_9_l_ofx_LC_12_11_4  (
            .in0(N__7750),
            .in1(N__14456),
            .in2(_gnd_net_),
            .in3(N__12383),
            .lcout(\ALU.addsub_axb_9_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_ma_LC_12_11_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_ma_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_ma_LC_12_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_ma_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__11586),
            .in2(_gnd_net_),
            .in3(N__7749),
            .lcout(\ALU.regsA_result_cry_5_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_4_LC_12_11_6.C_ON=1'b0;
    defparam b_4_LC_12_11_6.SEQ_MODE=4'b1000;
    defparam b_4_LC_12_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_4_LC_12_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10955),
            .lcout(bZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16101),
            .ce(N__11394),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_ma_LC_12_11_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_ma_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_ma_LC_12_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_ma_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__11585),
            .in2(_gnd_net_),
            .in3(N__14868),
            .lcout(\ALU.regsA_result_cry_3_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_LC_12_12_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_LC_12_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__8831),
            .in2(N__8096),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\ALU.regsA_result_cry_0_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNI9TCO2_LC_12_12_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNI9TCO2_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNI9TCO2_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNI9TCO2_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__8087),
            .in2(N__12158),
            .in3(N__8081),
            .lcout(\ALU.mult_AdderTree2_bigtree_530 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_0_2 ),
            .carryout(\ALU.regsA_result_cry_1_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_0_c_RNID4JS2_LC_12_12_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_0_c_RNID4JS2_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_0_c_RNID4JS2_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_0_c_RNID4JS2_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__12131),
            .in2(N__8078),
            .in3(N__8069),
            .lcout(\ALU.mult_AdderTree2_bigtree_531 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_3 ),
            .carryout(\ALU.regsA_result_cry_2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_0_c_RNIHBP03_LC_12_12_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_0_c_RNIHBP03_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_0_c_RNIHBP03_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_0_c_RNIHBP03_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__8066),
            .in2(N__8060),
            .in3(N__8051),
            .lcout(\ALU.mult_AdderTree2_bigtree_532 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_5 ),
            .carryout(\ALU.regsA_result_cry_3_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_0_c_RNILIVK2_LC_12_12_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_0_c_RNILIVK2_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_0_c_RNILIVK2_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_0_c_RNILIVK2_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__9737),
            .in2(N__8048),
            .in3(N__8039),
            .lcout(\ALU.mult_AdderTree2_bigtree_533 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_6 ),
            .carryout(\ALU.regsA_result_cry_4_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_0_c_RNIPP5P2_LC_12_12_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_0_c_RNIPP5P2_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_0_c_RNIPP5P2_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_0_c_RNIPP5P2_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__8036),
            .in2(N__9929),
            .in3(N__8030),
            .lcout(\ALU.mult_AdderTree2_bigtree_534 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_5 ),
            .carryout(\ALU.regsA_result_cry_5_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_0_c_RNIT0CT2_LC_12_12_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_0_c_RNIT0CT2_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_0_c_RNIT0CT2_LC_12_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_0_c_RNIT0CT2_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__9878),
            .in2(N__9944),
            .in3(N__8027),
            .lcout(\ALU.mult_AdderTree2_bigtree_535 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_6 ),
            .carryout(\ALU.regsA_result_cry_6_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_0_c_RNI18I13_LC_12_12_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_0_c_RNI18I13_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_0_c_RNI18I13_LC_12_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_0_c_RNI18I13_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__12503),
            .in2(N__8132),
            .in3(N__8123),
            .lcout(\ALU.mult_AdderTree2_bigtree_536 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_5 ),
            .carryout(\ALU.regsA_result_cry_7_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_0_c_RNI5FOL2_LC_12_13_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_0_c_RNI5FOL2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_0_c_RNI5FOL2_LC_12_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_0_c_RNI5FOL2_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__8213),
            .in2(N__12515),
            .in3(N__8120),
            .lcout(\ALU.mult_AdderTree2_bigtree_537 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\ALU.regsA_result_cry_8_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_0_c_RNIN2AT1_LC_12_13_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_0_c_RNIN2AT1_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_0_c_RNIN2AT1_LC_12_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_0_c_RNIN2AT1_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__14078),
            .in2(N__10871),
            .in3(N__8117),
            .lcout(\ALU.mult_AdderTree2_bigtree_538 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_8_2 ),
            .carryout(\ALU.regsA_result_cry_9_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_0_c_RNI206J1_LC_12_13_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_0_c_RNI206J1_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_0_c_RNI206J1_LC_12_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_0_c_RNI206J1_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__9626),
            .in2(N__9494),
            .in3(N__8114),
            .lcout(\ALU.mult_AdderTree2_bigtree_539 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_9_3 ),
            .carryout(\ALU.regsA_result_cry_10_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_0_c_RNIDUIG1_LC_12_13_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_0_c_RNIDUIG1_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_0_c_RNIDUIG1_LC_12_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_0_c_RNIDUIG1_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__8618),
            .in2(N__9641),
            .in3(N__8111),
            .lcout(\ALU.mult_AdderTree2_bigtree_540 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_10_2 ),
            .carryout(\ALU.regsA_result_cry_11_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_0_c_RNIH5PK1_LC_12_13_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_0_c_RNIH5PK1_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_0_c_RNIH5PK1_LC_12_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_0_c_RNIH5PK1_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__8825),
            .in2(N__8633),
            .in3(N__8108),
            .lcout(\ALU.mult_AdderTree2_bigtree_541 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_11_3 ),
            .carryout(\ALU.regsA_result_cry_12_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_0_c_RNILCVO1_LC_12_13_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_0_c_RNILCVO1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_0_c_RNILCVO1_LC_12_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_0_c_RNILCVO1_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__14669),
            .in2(N__8816),
            .in3(N__8105),
            .lcout(\ALU.mult_AdderTree2_bigtree_542 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_12_0 ),
            .carryout(\ALU.regsA_result_cry_13_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_0_c_RNIPJ5D1_LC_12_13_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_0_c_RNIPJ5D1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_0_c_RNIPJ5D1_LC_12_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_0_c_RNIPJ5D1_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__8228),
            .in2(N__8198),
            .in3(N__8102),
            .lcout(\ALU.mult_AdderTree2_bigtree_543 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_13_1 ),
            .carryout(\ALU.regsA_result_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_7_LC_12_13_7 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_7_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_7_LC_12_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_7_LC_12_13_7  (
            .in0(N__8204),
            .in1(N__8147),
            .in2(N__8846),
            .in3(N__8099),
            .lcout(\ALU.regsA_result_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_14_l_ofx_LC_12_14_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_14_l_ofx_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_14_l_ofx_LC_12_14_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_14_l_ofx_LC_12_14_0  (
            .in0(N__14255),
            .in1(N__12600),
            .in2(N__8176),
            .in3(N__14888),
            .lcout(\ALU.regsA_result_axb_14_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_7_l_ofx_LC_12_14_1 .C_ON=1'b0;
    defparam \ALU.addsub_axb_7_l_ofx_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_7_l_ofx_LC_12_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_7_l_ofx_LC_12_14_1  (
            .in0(N__12966),
            .in1(N__14445),
            .in2(_gnd_net_),
            .in3(N__12845),
            .lcout(\ALU.addsub_axb_7_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_ma_LC_12_14_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_ma_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_ma_LC_12_14_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_ma_LC_12_14_2  (
            .in0(N__12378),
            .in1(N__14885),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_8_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_14_LC_12_14_3 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_14_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_14_LC_12_14_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.overflow_RNO_14_LC_12_14_3  (
            .in0(N__13519),
            .in1(N__14578),
            .in2(N__12464),
            .in3(N__14256),
            .lcout(\ALU.regsA_result_axb_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_14_ma_LC_12_14_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_14_ma_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_14_ma_LC_12_14_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_14_ma_LC_12_14_4  (
            .in0(N__8168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14886),
            .lcout(\ALU.regsA_result_cry_14_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_1_l_ofx_LC_12_14_5 .C_ON=1'b0;
    defparam \ALU.addsub_axb_1_l_ofx_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_1_l_ofx_LC_12_14_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.addsub_axb_1_l_ofx_LC_12_14_5  (
            .in0(N__12602),
            .in1(_gnd_net_),
            .in2(N__12068),
            .in3(N__14444),
            .lcout(\ALU.addsub_axb_1_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_15_LC_12_14_6 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_15_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_15_LC_12_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.overflow_RNO_15_LC_12_14_6  (
            .in0(N__8169),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12601),
            .lcout(\ALU.overflow_RNOZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_0_l_ofx_LC_12_14_7 .C_ON=1'b0;
    defparam \ALU.addsub_axb_0_l_ofx_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_0_l_ofx_LC_12_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_0_l_ofx_LC_12_14_7  (
            .in0(N__14887),
            .in1(N__14443),
            .in2(_gnd_net_),
            .in3(N__13776),
            .lcout(\ALU.addsub_axb_0_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_LC_12_15_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_LC_12_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__10331),
            .in2(N__10472),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\ALU.regsA_result_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_5_LC_12_15_1 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_5_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_5_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_5_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__9026),
            .in2(N__10388),
            .in3(N__8414),
            .lcout(\ALU.mult_5 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_0 ),
            .carryout(\ALU.regsA_result_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_6_LC_12_15_2 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_6_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_6_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_6_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__8996),
            .in2(N__9845),
            .in3(N__8399),
            .lcout(\ALU.mult_6 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_0 ),
            .carryout(\ALU.regsA_result_cry_2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_7_LC_12_15_3 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_7_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_7_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_7_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__8966),
            .in2(N__9374),
            .in3(N__8396),
            .lcout(\ALU.mult_7 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_1 ),
            .carryout(\ALU.regsA_result_cry_3_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_3_c_RNI2M12C_LC_12_15_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_3_c_RNI2M12C_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_3_c_RNI2M12C_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_3_c_RNI2M12C_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__8933),
            .in2(N__9362),
            .in3(N__8372),
            .lcout(\ALU.mult_AdderTree2_bigtree_932 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_1 ),
            .carryout(\ALU.regsA_result_cry_4_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_4_c_RNILOTIB_LC_12_15_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_4_c_RNILOTIB_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_4_c_RNILOTIB_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_4_c_RNILOTIB_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__8903),
            .in2(N__9350),
            .in3(N__8354),
            .lcout(\ALU.mult_AdderTree2_bigtree_933 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_0 ),
            .carryout(\ALU.regsA_result_cry_5_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNIM757B_LC_12_15_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNIM757B_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNIM757B_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNIM757B_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__9260),
            .in2(N__9338),
            .in3(N__8321),
            .lcout(\ALU.mult_AdderTree2_bigtree_934 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_1 ),
            .carryout(\ALU.regsA_result_cry_6_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_6_c_RNIG0NPA_LC_12_15_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_6_c_RNIG0NPA_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_6_c_RNIG0NPA_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_6_c_RNIG0NPA_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__9233),
            .in2(N__9326),
            .in3(N__8288),
            .lcout(\ALU.mult_AdderTree2_bigtree_935 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_0 ),
            .carryout(\ALU.regsA_result_cry_7_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNIHGF5A_LC_12_16_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNIHGF5A_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNIHGF5A_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNIHGF5A_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__9206),
            .in2(N__9314),
            .in3(N__8258),
            .lcout(\ALU.mult_AdderTree2_bigtree_936 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\ALU.regsA_result_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_8_c_RNI026D9_LC_12_16_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_8_c_RNI026D9_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_8_c_RNI026D9_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_8_c_RNI026D9_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__9173),
            .in2(N__9302),
            .in3(N__8231),
            .lcout(\ALU.mult_AdderTree2_bigtree_937 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_8 ),
            .carryout(\ALU.regsA_result_cry_9_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_9_c_RNIQQNF9_LC_12_16_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_9_c_RNIQQNF9_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_9_c_RNIQQNF9_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_9_c_RNIQQNF9_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__9143),
            .in2(N__9290),
            .in3(N__8588),
            .lcout(\ALU.mult_AdderTree2_bigtree_938 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_9_0 ),
            .carryout(\ALU.regsA_result_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_10_c_RNIGPFR7_LC_12_16_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_10_c_RNIGPFR7_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_10_c_RNIGPFR7_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_10_c_RNIGPFR7_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__9515),
            .in2(N__9110),
            .in3(N__8561),
            .lcout(\ALU.mult_AdderTree2_bigtree_939 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_10 ),
            .carryout(\ALU.regsA_result_cry_11_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_1_LC_12_16_4 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_1_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_1_LC_12_16_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_1_LC_12_16_4  (
            .in0(N__8558),
            .in1(N__9086),
            .in2(N__8543),
            .in3(N__8528),
            .lcout(\ALU.regsA_result_axb_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_5_LC_12_16_5 .C_ON=1'b0;
    defparam \ALU.res_5_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \ALU.res_5_LC_12_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.res_5_LC_12_16_5  (
            .in0(N__8513),
            .in1(N__11265),
            .in2(_gnd_net_),
            .in3(N__8507),
            .lcout(res_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16114),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_7_LC_12_16_7 .C_ON=1'b0;
    defparam \ALU.res_7_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \ALU.res_7_LC_12_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_7_LC_12_16_7  (
            .in0(N__11279),
            .in1(N__8498),
            .in2(_gnd_net_),
            .in3(N__8489),
            .lcout(res_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16114),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_0_LC_12_17_1.C_ON=1'b0;
    defparam TXbuffer_0_LC_12_17_1.SEQ_MODE=4'b1000;
    defparam TXbuffer_0_LC_12_17_1.LUT_INIT=16'b1101111110000000;
    LogicCell40 TXbuffer_0_LC_12_17_1 (
            .in0(N__15908),
            .in1(N__8483),
            .in2(N__15674),
            .in3(N__8477),
            .lcout(TXbufferZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16119),
            .ce(N__9386),
            .sr(_gnd_net_));
    defparam TXbuffer_5_LC_12_17_3.C_ON=1'b0;
    defparam TXbuffer_5_LC_12_17_3.SEQ_MODE=4'b1000;
    defparam TXbuffer_5_LC_12_17_3.LUT_INIT=16'b0100111001000100;
    LogicCell40 TXbuffer_5_LC_12_17_3 (
            .in0(N__15906),
            .in1(N__8468),
            .in2(N__15675),
            .in3(N__8462),
            .lcout(TXbufferZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16119),
            .ce(N__9386),
            .sr(_gnd_net_));
    defparam TXbuffer_2_LC_12_17_4.C_ON=1'b0;
    defparam TXbuffer_2_LC_12_17_4.SEQ_MODE=4'b1000;
    defparam TXbuffer_2_LC_12_17_4.LUT_INIT=16'b0010001011110000;
    LogicCell40 TXbuffer_2_LC_12_17_4 (
            .in0(N__8437),
            .in1(N__15651),
            .in2(N__8423),
            .in3(N__15909),
            .lcout(TXbufferZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16119),
            .ce(N__9386),
            .sr(_gnd_net_));
    defparam TXbuffer_6_LC_12_17_6.C_ON=1'b0;
    defparam TXbuffer_6_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam TXbuffer_6_LC_12_17_6.LUT_INIT=16'b0011101100001000;
    LogicCell40 TXbuffer_6_LC_12_17_6 (
            .in0(N__8777),
            .in1(N__15910),
            .in2(N__15680),
            .in3(N__8768),
            .lcout(TXbufferZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16119),
            .ce(N__9386),
            .sr(_gnd_net_));
    defparam TXbuffer_7_LC_12_17_7.C_ON=1'b0;
    defparam TXbuffer_7_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam TXbuffer_7_LC_12_17_7.LUT_INIT=16'b0100111001000100;
    LogicCell40 TXbuffer_7_LC_12_17_7 (
            .in0(N__15907),
            .in1(N__8762),
            .in2(N__15676),
            .in3(N__8753),
            .lcout(TXbufferZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16119),
            .ce(N__9386),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_11_l_ofx_LC_13_9_4 .C_ON=1'b0;
    defparam \ALU.addsub_axb_11_l_ofx_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_11_l_ofx_LC_13_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_11_l_ofx_LC_13_9_4  (
            .in0(N__8746),
            .in1(N__14458),
            .in2(_gnd_net_),
            .in3(N__10275),
            .lcout(\ALU.addsub_axb_11_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_12_l_ofx_LC_13_10_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_12_l_ofx_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_12_l_ofx_LC_13_10_0 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_12_l_ofx_LC_13_10_0  (
            .in0(N__14570),
            .in1(N__12650),
            .in2(N__9594),
            .in3(N__14862),
            .lcout(\ALU.regsA_result_axb_12_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_12_LC_13_10_1.C_ON=1'b0;
    defparam b_12_LC_13_10_1.SEQ_MODE=4'b1000;
    defparam b_12_LC_13_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_12_LC_13_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10963),
            .lcout(bZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16090),
            .ce(N__14223),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_ma_LC_13_10_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_ma_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_ma_LC_13_10_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_ma_LC_13_10_2  (
            .in0(N__9582),
            .in1(N__14860),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_11_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_13_ma_LC_13_10_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_13_ma_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_13_ma_LC_13_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_13_ma_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__9583),
            .in2(_gnd_net_),
            .in3(N__13466),
            .lcout(\ALU.regsA_result_cry_13_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_13_l_ofx_LC_13_10_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_13_l_ofx_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_13_l_ofx_LC_13_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_13_l_ofx_LC_13_10_4  (
            .in0(N__13467),
            .in1(N__14560),
            .in2(N__9595),
            .in3(N__12453),
            .lcout(\ALU.regsA_result_axb_13_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_13_LC_13_10_5.C_ON=1'b0;
    defparam b_13_LC_13_10_5.SEQ_MODE=4'b1000;
    defparam b_13_LC_13_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_13_LC_13_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12287),
            .lcout(bZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16090),
            .ce(N__14223),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_ma_LC_13_10_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_ma_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_ma_LC_13_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_ma_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__14559),
            .in2(_gnd_net_),
            .in3(N__14861),
            .lcout(\ALU.regsA_result_cry_12_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_13_l_ofx_LC_13_10_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_13_l_ofx_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_13_l_ofx_LC_13_10_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_13_l_ofx_LC_13_10_7  (
            .in0(N__12651),
            .in1(N__14890),
            .in2(N__14571),
            .in3(N__14266),
            .lcout(\ALU.regsA_result_axb_13_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_LC_13_11_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_LC_13_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__9647),
            .in2(N__9656),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\ALU.regsA_result_cry_1_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNIF6113_LC_13_11_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNIF6113_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNIF6113_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNIF6113_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__9866),
            .in2(N__9713),
            .in3(N__8804),
            .lcout(\ALU.mult_AdderTree2_bigtree_565 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_8 ),
            .carryout(\ALU.regsA_result_cry_2_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_0_c_RNIJD753_LC_13_11_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_0_c_RNIJD753_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_0_c_RNIJD753_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_0_c_RNIJD753_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__9860),
            .in2(N__9704),
            .in3(N__8801),
            .lcout(\ALU.mult_AdderTree2_bigtree_566 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_10 ),
            .carryout(\ALU.regsA_result_cry_3_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_0_c_RNINKDP2_LC_13_11_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_0_c_RNINKDP2_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_0_c_RNINKDP2_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_0_c_RNINKDP2_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__9695),
            .in2(N__9854),
            .in3(N__8798),
            .lcout(\ALU.mult_AdderTree2_bigtree_567 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_10 ),
            .carryout(\ALU.regsA_result_cry_4_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_0_c_RNIRRJT2_LC_13_11_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_0_c_RNIRRJT2_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_0_c_RNIRRJT2_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_0_c_RNIRRJT2_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__8795),
            .in2(N__9689),
            .in3(N__8786),
            .lcout(\ALU.mult_AdderTree2_bigtree_568 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_9 ),
            .carryout(\ALU.regsA_result_cry_5_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_0_c_RNI1R903_LC_13_11_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_0_c_RNI1R903_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_0_c_RNI1R903_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_0_c_RNI1R903_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__9914),
            .in2(N__9728),
            .in3(N__8783),
            .lcout(\ALU.mult_AdderTree2_bigtree_569 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_9 ),
            .carryout(\ALU.regsA_result_cry_6_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_0_c_RNI52GK2_LC_13_11_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_0_c_RNI52GK2_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_0_c_RNI52GK2_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_0_c_RNI52GK2_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__9890),
            .in2(N__9902),
            .in3(N__8780),
            .lcout(\ALU.mult_AdderTree2_bigtree_570 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_8 ),
            .carryout(\ALU.regsA_result_cry_7_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_0_c_RNI99MO2_LC_13_11_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_0_c_RNI99MO2_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_0_c_RNI99MO2_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_0_c_RNI99MO2_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__9992),
            .in2(N__12491),
            .in3(N__8888),
            .lcout(\ALU.mult_AdderTree2_bigtree_571 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_7_7 ),
            .carryout(\ALU.regsA_result_cry_8_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_0_c_RNIDGSS2_LC_13_12_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_0_c_RNIDGSS2_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_0_c_RNIDGSS2_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_0_c_RNIDGSS2_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__12476),
            .in2(N__12404),
            .in3(N__8885),
            .lcout(\ALU.mult_AdderTree2_bigtree_572 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\ALU.regsA_result_cry_9_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_0_c_RNIODOI2_LC_13_12_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_0_c_RNIODOI2_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_0_c_RNIODOI2_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_0_c_RNIODOI2_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__9536),
            .in2(N__11126),
            .in3(N__8882),
            .lcout(\ALU.mult_AdderTree2_bigtree_573 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_9_5 ),
            .carryout(\ALU.regsA_result_cry_10_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_0_c_RNIHP7H1_LC_13_12_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_0_c_RNIHP7H1_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_0_c_RNIHP7H1_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_0_c_RNIHP7H1_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__9527),
            .in2(N__9611),
            .in3(N__8879),
            .lcout(\ALU.mult_AdderTree2_bigtree_574 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_10_4 ),
            .carryout(\ALU.regsA_result_cry_11_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_0_c_RNIL0EL1_LC_13_12_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_0_c_RNIL0EL1_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_0_c_RNIL0EL1_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_0_c_RNIL0EL1_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__8837),
            .in2(N__9551),
            .in3(N__8876),
            .lcout(\ALU.mult_AdderTree2_bigtree_575 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_11_4 ),
            .carryout(\ALU.regsA_result_cry_12_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_0_c_RNIP7K91_LC_13_12_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_0_c_RNIP7K91_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_0_c_RNIP7K91_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_0_c_RNIP7K91_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__8873),
            .in2(N__8864),
            .in3(N__8852),
            .lcout(\ALU.mult_AdderTree2_bigtree_576 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_12_1 ),
            .carryout(\ALU.regsA_result_cry_13_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_13_0_THRU_LUT4_0_LC_13_12_5 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_13_0_THRU_LUT4_0_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_13_0_THRU_LUT4_0_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_13_0_THRU_LUT4_0_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8849),
            .lcout(\ALU.regsA_result_cry_13_0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_ma_LC_13_12_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_ma_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_ma_LC_13_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_ma_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__10287),
            .in2(_gnd_net_),
            .in3(N__13468),
            .lcout(\ALU.regsA_result_cry_12_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_0_LC_13_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_0_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_0_LC_13_12_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_0_LC_13_12_7  (
            .in0(N__12013),
            .in1(N__14819),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_LC_13_13_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_LC_13_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__9743),
            .in2(N__9828),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\ALU.regsA_result_cry_0_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_3_LC_13_13_1 .C_ON=1'b1;
    defparam \ALU.res_RNO_1_3_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_3_LC_13_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.res_RNO_1_3_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__9680),
            .in2(N__9077),
            .in3(N__9068),
            .lcout(\ALU.mult_3 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_0_1 ),
            .carryout(\ALU.regsA_result_cry_1_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_1_c_RNITU8C6_LC_13_13_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_1_c_RNITU8C6_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_1_c_RNITU8C6_LC_13_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_1_c_RNITU8C6_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__9065),
            .in2(N__9059),
            .in3(N__9047),
            .lcout(\ALU.mult_AdderTree2_bigtree_796 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_2 ),
            .carryout(\ALU.regsA_result_cry_2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_2_c_RNI6FM46_LC_13_13_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_2_c_RNI6FM46_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_2_c_RNI6FM46_LC_13_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_2_c_RNI6FM46_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__9044),
            .in2(N__9038),
            .in3(N__9017),
            .lcout(\ALU.mult_AdderTree2_bigtree_797 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_3 ),
            .carryout(\ALU.regsA_result_cry_3_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_3_c_RNIFV3T5_LC_13_13_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_3_c_RNIFV3T5_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_3_c_RNIFV3T5_LC_13_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_3_c_RNIFV3T5_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__9014),
            .in2(N__9008),
            .in3(N__8987),
            .lcout(\ALU.mult_AdderTree2_bigtree_798 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_3 ),
            .carryout(\ALU.regsA_result_cry_4_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_4_c_RNIOFH56_LC_13_13_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_4_c_RNIOFH56_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_4_c_RNIOFH56_LC_13_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_4_c_RNIOFH56_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__8984),
            .in2(N__8978),
            .in3(N__8954),
            .lcout(\ALU.mult_AdderTree2_bigtree_799 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_2 ),
            .carryout(\ALU.regsA_result_cry_5_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_5_c_RNI3OEC6_LC_13_13_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_5_c_RNI3OEC6_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_5_c_RNI3OEC6_LC_13_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_5_c_RNI3OEC6_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__8951),
            .in2(N__8945),
            .in3(N__8924),
            .lcout(\ALU.mult_AdderTree2_bigtree_800 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_3 ),
            .carryout(\ALU.regsA_result_cry_6_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_6_c_RNIC8SK5_LC_13_13_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_6_c_RNIC8SK5_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_6_c_RNIC8SK5_LC_13_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_6_c_RNIC8SK5_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__8921),
            .in2(N__8915),
            .in3(N__8891),
            .lcout(\ALU.mult_AdderTree2_bigtree_801 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_2 ),
            .carryout(\ALU.regsA_result_cry_7_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_7_c_RNI35L05_LC_13_14_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_7_c_RNI35L05_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_7_c_RNI35L05_LC_13_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_7_c_RNI35L05_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__9278),
            .in2(N__9272),
            .in3(N__9254),
            .lcout(\ALU.mult_AdderTree2_bigtree_802 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\ALU.regsA_result_cry_8_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_8_c_RNIJBOQ4_LC_13_14_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_8_c_RNIJBOQ4_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_8_c_RNIJBOQ4_LC_13_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_8_c_RNIJBOQ4_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__9251),
            .in2(N__9245),
            .in3(N__9227),
            .lcout(\ALU.mult_AdderTree2_bigtree_803 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_8_0 ),
            .carryout(\ALU.regsA_result_cry_9_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_9_c_RNIA92E4_LC_13_14_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_9_c_RNIA92E4_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_9_c_RNIA92E4_LC_13_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_9_c_RNIA92E4_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__9224),
            .in2(N__9218),
            .in3(N__9194),
            .lcout(\ALU.mult_AdderTree2_bigtree_804 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_9_1 ),
            .carryout(\ALU.regsA_result_cry_10_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_10_c_RNIF8AD3_LC_13_14_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_10_c_RNIF8AD3_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_10_c_RNIF8AD3_LC_13_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_10_c_RNIF8AD3_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__9191),
            .in2(N__9185),
            .in3(N__9164),
            .lcout(\ALU.mult_AdderTree2_bigtree_805 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_10_0 ),
            .carryout(\ALU.regsA_result_cry_11_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_11_c_RNIOONL3_LC_13_14_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_11_c_RNIOONL3_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_11_c_RNIOONL3_LC_13_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_11_c_RNIOONL3_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__9161),
            .in2(N__9155),
            .in3(N__9134),
            .lcout(\ALU.mult_AdderTree2_bigtree_806 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_11_2 ),
            .carryout(\ALU.regsA_result_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_12_c_RNI195U2_LC_13_14_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_12_c_RNI195U2_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_12_c_RNI195U2_LC_13_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_12_c_RNI195U2_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__9131),
            .in2(N__9125),
            .in3(N__9098),
            .lcout(\ALU.mult_AdderTree2_bigtree_807 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_12 ),
            .carryout(\ALU.regsA_result_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_3_LC_13_14_6 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_3_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_3_LC_13_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_3_LC_13_14_6  (
            .in0(N__9503),
            .in1(N__9095),
            .in2(N__10016),
            .in3(N__9089),
            .lcout(\ALU.regsA_result_axb_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_LC_13_15_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_LC_13_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__13550),
            .in2(N__13905),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\ALU.regsA_result_cry_2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNIS7EJ4_LC_13_15_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNIS7EJ4_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNIS7EJ4_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNIS7EJ4_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__10445),
            .in2(N__9980),
            .in3(N__9365),
            .lcout(\ALU.mult_AdderTree2_bigtree_832 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_4 ),
            .carryout(\ALU.regsA_result_cry_3_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_3_c_RNIV8BJ5_LC_13_15_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_3_c_RNIV8BJ5_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_3_c_RNIV8BJ5_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_3_c_RNIV8BJ5_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__10655),
            .in2(N__9968),
            .in3(N__9353),
            .lcout(\ALU.mult_AdderTree2_bigtree_833 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_5 ),
            .carryout(\ALU.regsA_result_cry_4_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_4_c_RNI8POR5_LC_13_15_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_4_c_RNI8POR5_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_4_c_RNI8POR5_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_4_c_RNI8POR5_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__10631),
            .in2(N__9956),
            .in3(N__9341),
            .lcout(\ALU.mult_AdderTree2_bigtree_834 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_4 ),
            .carryout(\ALU.regsA_result_cry_5_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_5_c_RNIH9646_LC_13_15_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_5_c_RNIH9646_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_5_c_RNIH9646_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_5_c_RNIH9646_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__10610),
            .in2(N__10130),
            .in3(N__9329),
            .lcout(\ALU.mult_AdderTree2_bigtree_835 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_5 ),
            .carryout(\ALU.regsA_result_cry_6_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_6_c_RNIQPJS5_LC_13_15_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_6_c_RNIQPJS5_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_6_c_RNIQPJS5_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_6_c_RNIQPJS5_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__10586),
            .in2(N__10109),
            .in3(N__9317),
            .lcout(\ALU.mult_AdderTree2_bigtree_836 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_4 ),
            .carryout(\ALU.regsA_result_cry_7_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_7_c_RNI3A1L5_LC_13_15_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_7_c_RNI3A1L5_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_7_c_RNI3A1L5_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_7_c_RNI3A1L5_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__10562),
            .in2(N__10076),
            .in3(N__9305),
            .lcout(\ALU.mult_AdderTree2_bigtree_837 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_7_4 ),
            .carryout(\ALU.regsA_result_cry_8_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_8_c_RNICQET5_LC_13_15_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_8_c_RNICQET5_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_8_c_RNICQET5_LC_13_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_8_c_RNICQET5_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__10538),
            .in2(N__10064),
            .in3(N__9293),
            .lcout(\ALU.mult_AdderTree2_bigtree_838 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_8_1 ),
            .carryout(\ALU.regsA_result_cry_9_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_9_c_RNIS0IN5_LC_13_16_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_9_c_RNIS0IN5_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_9_c_RNIS0IN5_LC_13_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_9_c_RNIS0IN5_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__10052),
            .in2(N__10523),
            .in3(N__9281),
            .lcout(\ALU.mult_AdderTree2_bigtree_839 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\ALU.regsA_result_cry_10_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_10_c_RNI126N4_LC_13_16_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_10_c_RNI126N4_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_10_c_RNI126N4_LC_13_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_10_c_RNI126N4_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__10043),
            .in2(N__10766),
            .in3(N__9509),
            .lcout(\ALU.mult_AdderTree2_bigtree_840 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_10_1 ),
            .carryout(\ALU.regsA_result_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_11_THRU_LUT4_0_LC_13_16_2 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_11_THRU_LUT4_0_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_11_THRU_LUT4_0_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_11_THRU_LUT4_0_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9506),
            .lcout(\ALU.regsA_result_cry_11_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_fast_RNIP6NA1_3_LC_13_16_3 .C_ON=1'b0;
    defparam \FTDI.TXstate_fast_RNIP6NA1_3_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_fast_RNIP6NA1_3_LC_13_16_3 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \FTDI.TXstate_fast_RNIP6NA1_3_LC_13_16_3  (
            .in0(N__15662),
            .in1(N__15883),
            .in2(N__15785),
            .in3(N__16188),
            .lcout(TXstate_fast_RNIP6NA1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_10_l_ofx_LC_13_16_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_10_l_ofx_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_10_l_ofx_LC_13_16_4 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_10_l_ofx_LC_13_16_4  (
            .in0(N__14875),
            .in1(N__12649),
            .in2(N__14157),
            .in3(N__10292),
            .lcout(\ALU.regsA_result_axb_10_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_3_LC_13_16_7 .C_ON=1'b0;
    defparam \ALU.res_3_LC_13_16_7 .SEQ_MODE=4'b1000;
    defparam \ALU.res_3_LC_13_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_3_LC_13_16_7  (
            .in0(N__11264),
            .in1(N__9482),
            .in2(_gnd_net_),
            .in3(N__9470),
            .lcout(res_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16111),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_3_LC_13_17_1.C_ON=1'b0;
    defparam TXbuffer_3_LC_13_17_1.SEQ_MODE=4'b1000;
    defparam TXbuffer_3_LC_13_17_1.LUT_INIT=16'b0111001001010000;
    LogicCell40 TXbuffer_3_LC_13_17_1 (
            .in0(N__15911),
            .in1(N__15678),
            .in2(N__9461),
            .in3(N__9446),
            .lcout(TXbufferZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16115),
            .ce(N__9385),
            .sr(_gnd_net_));
    defparam TXbuffer_1_LC_13_17_4.C_ON=1'b0;
    defparam TXbuffer_1_LC_13_17_4.SEQ_MODE=4'b1000;
    defparam TXbuffer_1_LC_13_17_4.LUT_INIT=16'b0010001011110000;
    LogicCell40 TXbuffer_1_LC_13_17_4 (
            .in0(N__9427),
            .in1(N__15677),
            .in2(N__9410),
            .in3(N__15913),
            .lcout(TXbufferZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16115),
            .ce(N__9385),
            .sr(_gnd_net_));
    defparam TXbuffer_4_LC_13_17_5.C_ON=1'b0;
    defparam TXbuffer_4_LC_13_17_5.SEQ_MODE=4'b1000;
    defparam TXbuffer_4_LC_13_17_5.LUT_INIT=16'b0111001001010000;
    LogicCell40 TXbuffer_4_LC_13_17_5 (
            .in0(N__15912),
            .in1(N__15679),
            .in2(N__9398),
            .in3(N__11153),
            .lcout(TXbufferZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16115),
            .ce(N__9385),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_11_l_ofx_LC_14_9_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_11_l_ofx_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_11_l_ofx_LC_14_9_0 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_11_l_ofx_LC_14_9_0  (
            .in0(N__9581),
            .in1(N__12648),
            .in2(N__10276),
            .in3(N__14841),
            .lcout(\ALU.regsA_result_axb_11_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_11_LC_14_9_1.C_ON=1'b0;
    defparam b_11_LC_14_9_1.SEQ_MODE=4'b1000;
    defparam b_11_LC_14_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_11_LC_14_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10417),
            .lcout(bZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16080),
            .ce(N__14199),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_ma_LC_14_9_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_ma_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_ma_LC_14_9_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_ma_LC_14_9_2  (
            .in0(N__10258),
            .in1(N__14840),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_10_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_11_l_ofx_LC_14_9_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_11_l_ofx_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_11_l_ofx_LC_14_9_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_11_l_ofx_LC_14_9_4  (
            .in0(N__10262),
            .in1(N__12444),
            .in2(N__14162),
            .in3(N__13533),
            .lcout(\ALU.regsA_result_axb_11_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_13_LC_14_9_6 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_13_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_13_LC_14_9_6 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.overflow_RNO_13_LC_14_9_6  (
            .in0(N__15189),
            .in1(N__10271),
            .in2(N__9593),
            .in3(N__10852),
            .lcout(\ALU.regsA_result_axb_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_12_l_ofx_LC_14_9_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_12_l_ofx_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_12_l_ofx_LC_14_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_12_l_ofx_LC_14_9_7  (
            .in0(N__12443),
            .in1(N__13512),
            .in2(N__10286),
            .in3(N__9577),
            .lcout(\ALU.regsA_result_axb_12_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_10_l_ofx_LC_14_10_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_10_l_ofx_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_10_l_ofx_LC_14_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_10_l_ofx_LC_14_10_0  (
            .in0(N__12379),
            .in1(N__12442),
            .in2(N__13536),
            .in3(N__14149),
            .lcout(\ALU.regsA_result_axb_10_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_2_LC_14_10_1.C_ON=1'b0;
    defparam a_2_LC_14_10_1.SEQ_MODE=4'b1000;
    defparam a_2_LC_14_10_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_2_LC_14_10_1 (
            .in0(N__11107),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16084),
            .ce(N__15275),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_ma_LC_14_10_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_ma_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_ma_LC_14_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_ma_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__14148),
            .in2(_gnd_net_),
            .in3(N__13463),
            .lcout(\ALU.regsA_result_cry_11_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_2_rep1_LC_14_10_3.C_ON=1'b0;
    defparam a_2_rep1_LC_14_10_3.SEQ_MODE=4'b1000;
    defparam a_2_rep1_LC_14_10_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_2_rep1_LC_14_10_3 (
            .in0(N__11108),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_2_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16084),
            .ce(N__15275),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_2_l_ofx_LC_14_10_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_2_l_ofx_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_2_l_ofx_LC_14_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_2_l_ofx_LC_14_10_4  (
            .in0(N__11946),
            .in1(N__11746),
            .in2(N__13537),
            .in3(N__9769),
            .lcout(\ALU.regsA_result_axb_2_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_3_l_ofx_LC_14_10_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_3_l_ofx_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_3_l_ofx_LC_14_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_3_l_ofx_LC_14_10_5  (
            .in0(N__13464),
            .in1(N__11797),
            .in2(N__9789),
            .in3(N__13285),
            .lcout(\ALU.regsA_result_axb_3_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_4_l_ofx_LC_14_10_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_4_l_ofx_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_4_l_ofx_LC_14_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_4_l_ofx_LC_14_10_6  (
            .in0(N__13286),
            .in1(N__11644),
            .in2(N__13538),
            .in3(N__9773),
            .lcout(\ALU.regsA_result_axb_4_l_ofx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_5_l_ofx_LC_14_10_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_5_l_ofx_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_5_l_ofx_LC_14_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_5_l_ofx_LC_14_10_7  (
            .in0(N__13465),
            .in1(N__11645),
            .in2(N__9790),
            .in3(N__15024),
            .lcout(\ALU.regsA_result_axb_5_l_ofx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_1_LC_14_11_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_1_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_1_LC_14_11_0 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_1_LC_14_11_0  (
            .in0(N__13726),
            .in1(N__13439),
            .in2(N__9671),
            .in3(N__11945),
            .lcout(\ALU.mult_AdderTree2_bigtree_564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_fast_2_LC_14_11_1.C_ON=1'b0;
    defparam a_fast_2_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam a_fast_2_LC_14_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_fast_2_LC_14_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11105),
            .lcout(a_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16091),
            .ce(N__15249),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_LC_14_11_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_LC_14_11_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_LC_14_11_2  (
            .in0(N__13727),
            .in1(N__13440),
            .in2(N__11993),
            .in3(N__9667),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_3_LC_14_11_3.C_ON=1'b0;
    defparam a_3_LC_14_11_3.SEQ_MODE=4'b1000;
    defparam a_3_LC_14_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_3_LC_14_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10420),
            .lcout(aZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16091),
            .ce(N__15249),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_0_LC_14_11_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_0_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_0_LC_14_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_0_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__13642),
            .in2(_gnd_net_),
            .in3(N__13435),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_ma_LC_14_11_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_ma_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_ma_LC_14_11_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_ma_LC_14_11_5  (
            .in0(N__13436),
            .in1(N__11944),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_2_ma_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_ma_LC_14_11_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_ma_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_ma_LC_14_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_ma_LC_14_11_6  (
            .in0(N__11749),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13437),
            .lcout(\ALU.regsA_result_cry_3_ma_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_ma_LC_14_11_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_ma_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_ma_LC_14_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_ma_LC_14_11_7  (
            .in0(N__13438),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13287),
            .lcout(\ALU.regsA_result_cry_4_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNIUA504_LC_14_12_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNIUA504_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNIUA504_LC_14_12_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNIUA504_LC_14_12_0  (
            .in0(N__13906),
            .in1(N__13869),
            .in2(_gnd_net_),
            .in3(N__13670),
            .lcout(\ALU.mult_AdderTree2_bigtree_831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_0_LC_14_12_1.C_ON=1'b0;
    defparam b_0_LC_14_12_1.SEQ_MODE=4'b1000;
    defparam b_0_LC_14_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_0_LC_14_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14503),
            .lcout(bZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16096),
            .ce(N__11396),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_14_12_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_14_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_14_12_2  (
            .in0(N__9830),
            .in1(N__9791),
            .in2(_gnd_net_),
            .in3(N__13669),
            .lcout(\ALU.regsA_result_cry_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_ma_LC_14_12_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_ma_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_ma_LC_14_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_ma_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__14998),
            .in2(_gnd_net_),
            .in3(N__14820),
            .lcout(\ALU.regsA_result_cry_4_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_5_LC_14_12_6.C_ON=1'b0;
    defparam b_5_LC_14_12_6.SEQ_MODE=4'b1000;
    defparam b_5_LC_14_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_5_LC_14_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12282),
            .lcout(bZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16096),
            .ce(N__11396),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_ma_LC_14_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_ma_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_ma_LC_14_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_ma_LC_14_12_7  (
            .in0(N__13434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14999),
            .lcout(\ALU.regsA_result_cry_6_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_6_l_ofx_LC_14_13_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_6_l_ofx_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_6_l_ofx_LC_14_13_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_6_l_ofx_LC_14_13_0  (
            .in0(N__12806),
            .in1(N__14832),
            .in2(N__13068),
            .in3(N__12607),
            .lcout(\ALU.regsA_result_axb_6_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_6_LC_14_13_1.C_ON=1'b0;
    defparam b_6_LC_14_13_1.SEQ_MODE=4'b1000;
    defparam b_6_LC_14_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_6_LC_14_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14307),
            .lcout(bZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16102),
            .ce(N__11387),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_ma_LC_14_13_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_ma_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_ma_LC_14_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_ma_LC_14_13_2  (
            .in0(N__13032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14831),
            .lcout(\ALU.regsA_result_cry_5_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_6_l_ofx_LC_14_13_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_6_l_ofx_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_6_l_ofx_LC_14_13_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_6_l_ofx_LC_14_13_4  (
            .in0(N__15001),
            .in1(N__15188),
            .in2(N__13067),
            .in3(N__10833),
            .lcout(\ALU.regsA_result_axb_6_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_6_l_ofx_LC_14_13_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_6_l_ofx_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_6_l_ofx_LC_14_13_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_6_l_ofx_LC_14_13_5  (
            .in0(N__12454),
            .in1(N__13039),
            .in2(N__13521),
            .in3(N__15000),
            .lcout(\ALU.regsA_result_axb_6_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_ma_LC_14_13_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_ma_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_ma_LC_14_13_6 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_ma_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__13488),
            .in2(N__13069),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_7_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_7_l_ofx_LC_14_13_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_7_l_ofx_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_7_l_ofx_LC_14_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_7_l_ofx_LC_14_13_7  (
            .in0(N__12455),
            .in1(N__13043),
            .in2(N__13522),
            .in3(N__12805),
            .lcout(\ALU.regsA_result_axb_7_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_7_LC_14_14_1.C_ON=1'b0;
    defparam b_7_LC_14_14_1.SEQ_MODE=4'b1000;
    defparam b_7_LC_14_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_7_LC_14_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12115),
            .lcout(bZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16104),
            .ce(N__11395),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_ma_LC_14_14_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_ma_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_ma_LC_14_14_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_ma_LC_14_14_2  (
            .in0(N__12801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14847),
            .lcout(\ALU.regsA_result_cry_6_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_ma_LC_14_14_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_ma_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_ma_LC_14_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_ma_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__12803),
            .in2(_gnd_net_),
            .in3(N__15180),
            .lcout(\ALU.regsA_result_cry_8_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_7_l_ofx_LC_14_14_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_7_l_ofx_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_7_l_ofx_LC_14_14_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_7_l_ofx_LC_14_14_4  (
            .in0(N__15181),
            .in1(N__13054),
            .in2(N__10847),
            .in3(N__12831),
            .lcout(\ALU.regsA_result_axb_7_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_ma_LC_14_14_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_ma_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_ma_LC_14_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_ma_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__12802),
            .in2(_gnd_net_),
            .in3(N__13495),
            .lcout(\ALU.regsA_result_cry_8_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_8_l_ofx_LC_14_14_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_8_l_ofx_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_8_l_ofx_LC_14_14_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_8_l_ofx_LC_14_14_6  (
            .in0(N__15182),
            .in1(N__12832),
            .in2(N__10848),
            .in3(N__13171),
            .lcout(\ALU.regsA_result_axb_8_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_7_l_ofx_LC_14_14_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_7_l_ofx_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_7_l_ofx_LC_14_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_7_l_ofx_LC_14_14_7  (
            .in0(N__13055),
            .in1(N__13867),
            .in2(N__12968),
            .in3(N__12804),
            .lcout(\ALU.regsA_result_axb_7_l_ofx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_LC_14_15_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__10370),
            .in2(N__10700),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\ALU.regsA_result_cry_1_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNI5R443_LC_14_15_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNI5R443_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNI5R443_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNI5R443_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__10358),
            .in2(N__10724),
            .in3(N__9983),
            .lcout(\ALU.mult_AdderTree2_bigtree_600 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_7 ),
            .carryout(\ALU.regsA_result_cry_2_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_0_c_RNI92BO2_LC_14_15_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_0_c_RNI92BO2_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_0_c_RNI92BO2_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_0_c_RNI92BO2_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__12143),
            .in2(N__10346),
            .in3(N__9971),
            .lcout(\ALU.mult_AdderTree2_bigtree_601 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_9 ),
            .carryout(\ALU.regsA_result_cry_3_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_0_c_RNI0ARQ2_LC_14_15_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_0_c_RNI0ARQ2_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_0_c_RNI0ARQ2_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_0_c_RNI0ARQ2_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__10889),
            .in2(N__10682),
            .in3(N__9959),
            .lcout(\ALU.mult_AdderTree2_bigtree_602 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_9 ),
            .carryout(\ALU.regsA_result_cry_4_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_0_c_RNI4H1V2_LC_14_15_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_0_c_RNI4H1V2_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_0_c_RNI4H1V2_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_0_c_RNI4H1V2_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__10883),
            .in2(N__10910),
            .in3(N__9947),
            .lcout(\ALU.mult_AdderTree2_bigtree_603 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_8 ),
            .carryout(\ALU.regsA_result_cry_5_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_0_c_RNI8O733_LC_14_15_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_0_c_RNI8O733_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_0_c_RNI8O733_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_0_c_RNI8O733_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__10877),
            .in2(N__10142),
            .in3(N__10121),
            .lcout(\ALU.mult_AdderTree2_bigtree_604 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_8 ),
            .carryout(\ALU.regsA_result_cry_6_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_0_c_RNICVDN2_LC_14_15_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_0_c_RNICVDN2_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_0_c_RNICVDN2_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_0_c_RNICVDN2_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__10715),
            .in2(N__10118),
            .in3(N__10100),
            .lcout(\ALU.mult_AdderTree2_bigtree_605 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_7 ),
            .carryout(\ALU.regsA_result_cry_7_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_0_c_RNIG6KR2_LC_14_15_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_0_c_RNIG6KR2_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_0_c_RNIG6KR2_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_0_c_RNIG6KR2_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__10097),
            .in2(N__10088),
            .in3(N__10067),
            .lcout(\ALU.mult_AdderTree2_bigtree_606 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_7_6 ),
            .carryout(\ALU.regsA_result_cry_8_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_0_c_RNIKDQV2_LC_14_16_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_0_c_RNIKDQV2_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_0_c_RNIKDQV2_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_0_c_RNIKDQV2_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__10736),
            .in2(N__10775),
            .in3(N__10055),
            .lcout(\ALU.mult_AdderTree2_bigtree_607 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\ALU.regsA_result_cry_9_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_0_c_RNIVAML2_LC_14_16_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_0_c_RNIVAML2_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_0_c_RNIVAML2_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_0_c_RNIVAML2_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__10217),
            .in2(N__10001),
            .in3(N__10046),
            .lcout(\ALU.mult_AdderTree2_bigtree_608 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_9_4 ),
            .carryout(\ALU.regsA_result_cry_10_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_0_c_RNIONSH1_LC_14_16_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_0_c_RNIONSH1_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_0_c_RNIONSH1_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_0_c_RNIONSH1_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__10298),
            .in2(N__10226),
            .in3(N__10037),
            .lcout(\ALU.mult_AdderTree2_bigtree_609 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_10_3 ),
            .carryout(\ALU.regsA_result_cry_11_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_6_LC_14_16_3 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_6_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_6_LC_14_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.overflow_RNO_6_LC_14_16_3  (
            .in0(N__10709),
            .in1(N__10745),
            .in2(N__10034),
            .in3(N__10019),
            .lcout(\ALU.regsA_result_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_10_l_ofx_LC_14_16_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_10_l_ofx_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_10_l_ofx_LC_14_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_10_l_ofx_LC_14_16_4  (
            .in0(N__12355),
            .in1(N__10828),
            .in2(N__15205),
            .in3(N__14127),
            .lcout(\ALU.regsA_result_axb_10_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_11_ma_LC_14_16_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_11_ma_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_11_ma_LC_14_16_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_11_ma_LC_14_16_5  (
            .in0(N__14128),
            .in1(_gnd_net_),
            .in2(N__15206),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_11_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_11_l_ofx_LC_14_16_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_11_l_ofx_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_11_l_ofx_LC_14_16_6 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_11_l_ofx_LC_14_16_6  (
            .in0(N__15199),
            .in1(N__10829),
            .in2(N__10291),
            .in3(N__14129),
            .lcout(\ALU.regsA_result_axb_11_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_ma_LC_14_16_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_ma_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_ma_LC_14_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_ma_LC_14_16_7  (
            .in0(N__15200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12354),
            .lcout(\ALU.regsA_result_cry_10_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_1_LC_14_17_0 .C_ON=1'b0;
    defparam \FTDI.TXshift_1_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_1_LC_14_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \FTDI.TXshift_1_LC_14_17_0  (
            .in0(N__10196),
            .in1(N__15424),
            .in2(_gnd_net_),
            .in3(N__10211),
            .lcout(\FTDI.TXshiftZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_2_LC_14_17_1 .C_ON=1'b0;
    defparam \FTDI.TXshift_2_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_2_LC_14_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_2_LC_14_17_1  (
            .in0(N__15425),
            .in1(N__10148),
            .in2(_gnd_net_),
            .in3(N__10205),
            .lcout(\FTDI.TXshiftZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_6_LC_14_17_2 .C_ON=1'b0;
    defparam \FTDI.TXshift_6_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_6_LC_14_17_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \FTDI.TXshift_6_LC_14_17_2  (
            .in0(N__11030),
            .in1(N__15429),
            .in2(_gnd_net_),
            .in3(N__10190),
            .lcout(\FTDI.TXshiftZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_4_LC_14_17_3 .C_ON=1'b0;
    defparam \FTDI.TXshift_4_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_4_LC_14_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_4_LC_14_17_3  (
            .in0(N__15427),
            .in1(N__10304),
            .in2(_gnd_net_),
            .in3(N__10181),
            .lcout(\FTDI.TXshiftZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_0_LC_14_17_4 .C_ON=1'b0;
    defparam \FTDI.TXshift_0_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_0_LC_14_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \FTDI.TXshift_0_LC_14_17_4  (
            .in0(N__10175),
            .in1(N__15423),
            .in2(_gnd_net_),
            .in3(N__10169),
            .lcout(\FTDI.TXshiftZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_3_LC_14_17_6 .C_ON=1'b0;
    defparam \FTDI.TXshift_3_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_3_LC_14_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_3_LC_14_17_6  (
            .in0(N__10160),
            .in1(N__10154),
            .in2(_gnd_net_),
            .in3(N__15426),
            .lcout(\FTDI.TXshiftZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_5_LC_14_17_7 .C_ON=1'b0;
    defparam \FTDI.TXshift_5_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_5_LC_14_17_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_5_LC_14_17_7  (
            .in0(N__15428),
            .in1(N__10319),
            .in2(_gnd_net_),
            .in3(N__10313),
            .lcout(\FTDI.TXshiftZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__12713),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_2_LC_15_8_2 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_2_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_2_LC_15_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_2_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10418),
            .lcout(RXbuffer_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_2C_net ),
            .ce(N__10993),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_4_LC_15_8_3 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_4_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_4_LC_15_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_4_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12271),
            .lcout(RXbuffer_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_2C_net ),
            .ce(N__10993),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_3_LC_15_8_5 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_3_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_3_LC_15_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_3_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10942),
            .lcout(RXbuffer_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_2C_net ),
            .ce(N__10993),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_7_LC_15_8_7 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_7_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_7_LC_15_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_7_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11024),
            .lcout(RXbuffer_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_2C_net ),
            .ce(N__10993),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_5_LC_15_9_1 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_5_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_5_LC_15_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_5_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14296),
            .lcout(RXbuffer_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_5C_net ),
            .ce(N__10997),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_0_LC_15_9_2 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_0_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_0_LC_15_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_0_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11320),
            .lcout(RXbuffer_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_5C_net ),
            .ce(N__10997),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_6_LC_15_9_3 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_6_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_6_LC_15_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_6_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12103),
            .lcout(RXbuffer_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_5C_net ),
            .ce(N__10997),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_1_LC_15_9_6 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_1_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_1_LC_15_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_1_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11084),
            .lcout(RXbuffer_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_5C_net ),
            .ce(N__10997),
            .sr(_gnd_net_));
    defparam b_1_LC_15_10_0.C_ON=1'b0;
    defparam b_1_LC_15_10_0.SEQ_MODE=4'b1000;
    defparam b_1_LC_15_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_1_LC_15_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11314),
            .lcout(bZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16081),
            .ce(N__11374),
            .sr(_gnd_net_));
    defparam b_2_LC_15_10_1.C_ON=1'b0;
    defparam b_2_LC_15_10_1.SEQ_MODE=4'b1000;
    defparam b_2_LC_15_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_2_LC_15_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11094),
            .lcout(bZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16081),
            .ce(N__11374),
            .sr(_gnd_net_));
    defparam b_3_LC_15_10_2.C_ON=1'b0;
    defparam b_3_LC_15_10_2.SEQ_MODE=4'b1000;
    defparam b_3_LC_15_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_3_LC_15_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10419),
            .lcout(bZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16081),
            .ce(N__11374),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_1_LC_15_11_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_1_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_1_LC_15_11_0 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_1_LC_15_11_0  (
            .in0(N__13671),
            .in1(N__15159),
            .in2(N__11948),
            .in3(N__10505),
            .lcout(\ALU.mult_AdderTree2_bigtree_599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_fast_4_LC_15_11_1.C_ON=1'b0;
    defparam a_fast_4_LC_15_11_1.SEQ_MODE=4'b1000;
    defparam a_fast_4_LC_15_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_fast_4_LC_15_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10943),
            .lcout(a_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16085),
            .ce(N__15264),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_LC_15_11_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_LC_15_11_2 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_LC_15_11_2  (
            .in0(N__13674),
            .in1(N__10491),
            .in2(N__11947),
            .in3(N__15161),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_2_l_ofx_LC_15_11_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_2_l_ofx_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_2_l_ofx_LC_15_11_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_2_l_ofx_LC_15_11_3  (
            .in0(N__15160),
            .in1(N__11904),
            .in2(N__10503),
            .in3(N__11747),
            .lcout(\ALU.regsA_result_axb_2_l_ofx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_3_l_ofx_LC_15_11_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_3_l_ofx_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_3_l_ofx_LC_15_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_3_l_ofx_LC_15_11_4  (
            .in0(N__11748),
            .in1(N__10495),
            .in2(N__15190),
            .in3(N__13252),
            .lcout(\ALU.regsA_result_axb_3_l_ofx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_15_11_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_15_11_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_15_11_5  (
            .in0(N__10471),
            .in1(_gnd_net_),
            .in2(N__10504),
            .in3(N__13672),
            .lcout(\ALU.regsA_result_cry_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_RNO_1_4_LC_15_11_6 .C_ON=1'b0;
    defparam \ALU.res_RNO_1_4_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.res_RNO_1_4_LC_15_11_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ALU.res_RNO_1_4_LC_15_11_6  (
            .in0(N__13673),
            .in1(N__10499),
            .in2(_gnd_net_),
            .in3(N__10470),
            .lcout(\ALU.mult_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_5_LC_15_11_7.C_ON=1'b0;
    defparam a_5_LC_15_11_7.SEQ_MODE=4'b1000;
    defparam a_5_LC_15_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_5_LC_15_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12286),
            .lcout(aZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16085),
            .ce(N__15264),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_1_LC_15_12_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_1_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_1_LC_15_12_0 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_1_LC_15_12_0  (
            .in0(N__12940),
            .in1(N__13643),
            .in2(N__13873),
            .in3(N__11967),
            .lcout(\ALU.mult_AdderTree2_bigtree_634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_6_LC_15_12_1.C_ON=1'b0;
    defparam a_6_LC_15_12_1.SEQ_MODE=4'b1000;
    defparam a_6_LC_15_12_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 a_6_LC_15_12_1 (
            .in0(N__14297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16092),
            .ce(N__15285),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_LC_15_12_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_LC_15_12_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_LC_15_12_2  (
            .in0(N__12948),
            .in1(N__13644),
            .in2(N__11994),
            .in3(N__13828),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_2_l_ofx_LC_15_12_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_2_l_ofx_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_2_l_ofx_LC_15_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_2_l_ofx_LC_15_12_3  (
            .in0(N__11968),
            .in1(N__12941),
            .in2(N__13864),
            .in3(N__11781),
            .lcout(\ALU.regsA_result_axb_2_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_3_l_ofx_LC_15_12_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_3_l_ofx_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_3_l_ofx_LC_15_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_3_l_ofx_LC_15_12_4  (
            .in0(N__11782),
            .in1(N__13297),
            .in2(N__12962),
            .in3(N__13832),
            .lcout(\ALU.regsA_result_axb_3_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_4_l_ofx_LC_15_12_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_4_l_ofx_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_4_l_ofx_LC_15_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_4_l_ofx_LC_15_12_5  (
            .in0(N__13298),
            .in1(N__12945),
            .in2(N__13865),
            .in3(N__11646),
            .lcout(\ALU.regsA_result_axb_4_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_5_l_ofx_LC_15_12_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_5_l_ofx_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_5_l_ofx_LC_15_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_5_l_ofx_LC_15_12_6  (
            .in0(N__12946),
            .in1(N__13836),
            .in2(N__11662),
            .in3(N__14987),
            .lcout(\ALU.regsA_result_axb_5_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_6_l_ofx_LC_15_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_6_l_ofx_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_6_l_ofx_LC_15_12_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_6_l_ofx_LC_15_12_7  (
            .in0(N__14988),
            .in1(N__12947),
            .in2(N__13866),
            .in3(N__13044),
            .lcout(\ALU.regsA_result_axb_6_l_ofx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_LC_15_13_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__10691),
            .in2(N__10673),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\ALU.regsA_result_cry_1_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNIVOCL2_LC_15_13_1 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNIVOCL2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNIVOCL2_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNIVOCL2_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__11840),
            .in2(N__10664),
            .in3(N__10643),
            .lcout(\ALU.mult_AdderTree2_bigtree_635 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_1_9 ),
            .carryout(\ALU.regsA_result_cry_2_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_0_c_RNI30JP2_LC_15_13_2 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_0_c_RNI30JP2_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_0_c_RNI30JP2_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_0_c_RNI30JP2_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__11678),
            .in2(N__10640),
            .in3(N__10619),
            .lcout(\ALU.mult_AdderTree2_bigtree_636 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_2_11 ),
            .carryout(\ALU.regsA_result_cry_3_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_0_c_RNI77PT2_LC_15_13_3 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_0_c_RNI77PT2_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_0_c_RNI77PT2_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_0_c_RNI77PT2_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__10616),
            .in2(N__11672),
            .in3(N__10598),
            .lcout(\ALU.mult_AdderTree2_bigtree_637 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_3_11 ),
            .carryout(\ALU.regsA_result_cry_4_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_0_c_RNIBEV13_LC_15_13_4 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_0_c_RNIBEV13_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_0_c_RNIBEV13_LC_15_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_0_c_RNIBEV13_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__11522),
            .in2(N__10595),
            .in3(N__10574),
            .lcout(\ALU.mult_AdderTree2_bigtree_638 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_4_10 ),
            .carryout(\ALU.regsA_result_cry_5_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_0_c_RNIFL5M2_LC_15_13_5 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_0_c_RNIFL5M2_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_0_c_RNIFL5M2_LC_15_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_0_c_RNIFL5M2_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__12659),
            .in2(N__10571),
            .in3(N__10550),
            .lcout(\ALU.mult_AdderTree2_bigtree_639 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_5_10 ),
            .carryout(\ALU.regsA_result_cry_6_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_0_c_RNIJSBQ2_LC_15_13_6 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_0_c_RNIJSBQ2_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_0_c_RNIJSBQ2_LC_15_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_0_c_RNIJSBQ2_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__12974),
            .in2(N__10547),
            .in3(N__10526),
            .lcout(\ALU.mult_AdderTree2_bigtree_640 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_6_9 ),
            .carryout(\ALU.regsA_result_cry_7_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_0_c_RNIN3IU2_LC_15_13_7 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_0_c_RNIN3IU2_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_0_c_RNIN3IU2_LC_15_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_0_c_RNIN3IU2_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__12389),
            .in2(N__12761),
            .in3(N__10508),
            .lcout(\ALU.mult_AdderTree2_bigtree_641 ),
            .ltout(),
            .carryin(\ALU.regsA_result_cry_7_8 ),
            .carryout(\ALU.regsA_result_cry_8_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_0_c_RNIRAO23_LC_15_14_0 .C_ON=1'b1;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_0_c_RNIRAO23_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_0_c_RNIRAO23_LC_15_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_0_c_RNIRAO23_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__13097),
            .in2(N__12296),
            .in3(N__10751),
            .lcout(\ALU.mult_AdderTree2_bigtree_642 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\ALU.regsA_result_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.regsA_result_cry_9_THRU_LUT4_0_LC_15_14_1 .C_ON=1'b0;
    defparam \ALU.regsA_result_cry_9_THRU_LUT4_0_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.regsA_result_cry_9_THRU_LUT4_0_LC_15_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.regsA_result_cry_9_THRU_LUT4_0_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10748),
            .lcout(\ALU.regsA_result_cry_9_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_ma_LC_15_14_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_ma_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_ma_LC_15_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_ma_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__13153),
            .in2(_gnd_net_),
            .in3(N__15134),
            .lcout(\ALU.regsA_result_cry_9_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_ma_LC_15_14_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_ma_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_ma_LC_15_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_ma_LC_15_14_3  (
            .in0(N__15133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11970),
            .lcout(\ALU.regsA_result_cry_2_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_ma_LC_15_14_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_ma_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_ma_LC_15_14_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_ma_LC_15_14_4  (
            .in0(N__13045),
            .in1(N__15135),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_7_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.overflow_RNO_12_LC_15_14_5 .C_ON=1'b0;
    defparam \ALU.overflow_RNO_12_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.overflow_RNO_12_LC_15_14_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.overflow_RNO_12_LC_15_14_5  (
            .in0(N__12371),
            .in1(N__13868),
            .in2(N__14153),
            .in3(N__12939),
            .lcout(\ALU.regsA_result_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_0_LC_15_14_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_0_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_0_LC_15_14_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_0_LC_15_14_6  (
            .in0(N__13676),
            .in1(N__15132),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_0_LC_15_14_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_0_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_0_LC_15_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_0_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__13675),
            .in2(_gnd_net_),
            .in3(N__12938),
            .lcout(\ALU.regsA_result_cry_1_0_c_RNO_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_4_l_ofx_LC_15_15_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_4_l_ofx_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_4_l_ofx_LC_15_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_4_l_ofx_LC_15_15_0  (
            .in0(N__13346),
            .in1(N__11651),
            .in2(N__15179),
            .in3(N__10822),
            .lcout(\ALU.regsA_result_axb_4_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_4_LC_15_15_1.C_ON=1'b0;
    defparam a_4_LC_15_15_1.SEQ_MODE=4'b1000;
    defparam a_4_LC_15_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_4_LC_15_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10956),
            .lcout(aZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16105),
            .ce(N__15296),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_5_l_ofx_LC_15_15_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_5_l_ofx_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_5_l_ofx_LC_15_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_5_l_ofx_LC_15_15_2  (
            .in0(N__15142),
            .in1(N__10823),
            .in2(N__11663),
            .in3(N__15017),
            .lcout(\ALU.regsA_result_axb_5_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_4_l_ofx_LC_15_15_3 .C_ON=1'b0;
    defparam \ALU.addsub_axb_4_l_ofx_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_4_l_ofx_LC_15_15_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.addsub_axb_4_l_ofx_LC_15_15_3  (
            .in0(N__11653),
            .in1(_gnd_net_),
            .in2(N__10843),
            .in3(N__14426),
            .lcout(\ALU.addsub_axb_4_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_ma_LC_15_15_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_ma_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_ma_LC_15_15_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_ma_LC_15_15_5  (
            .in0(N__13296),
            .in1(N__15136),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_4_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_ma_LC_15_15_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_ma_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_ma_LC_15_15_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_ma_LC_15_15_6  (
            .in0(N__15137),
            .in1(N__11652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_5_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_ma_LC_15_15_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_ma_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_ma_LC_15_15_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_ma_LC_15_15_7  (
            .in0(N__15018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15138),
            .lcout(\ALU.regsA_result_cry_6_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_9_l_ofx_LC_15_16_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_9_l_ofx_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_9_l_ofx_LC_15_16_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_9_l_ofx_LC_15_16_0  (
            .in0(N__14130),
            .in1(N__14874),
            .in2(N__12652),
            .in3(N__12353),
            .lcout(\ALU.regsA_result_axb_9_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_9_LC_15_16_1.C_ON=1'b0;
    defparam b_9_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam b_9_LC_15_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_9_LC_15_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11331),
            .lcout(bZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16107),
            .ce(N__14224),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_9_l_ofx_LC_15_16_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_9_l_ofx_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_9_l_ofx_LC_15_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_9_l_ofx_LC_15_16_3  (
            .in0(N__15195),
            .in1(N__12352),
            .in2(N__13184),
            .in3(N__10827),
            .lcout(\ALU.regsA_result_axb_9_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_ma_LC_15_16_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_ma_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_ma_LC_15_16_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_ma_LC_15_16_6  (
            .in0(N__12351),
            .in1(N__13534),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_10_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_10_LC_15_16_7.C_ON=1'b0;
    defparam b_10_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam b_10_LC_15_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_10_LC_15_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11099),
            .lcout(bZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16107),
            .ce(N__14224),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_7_LC_15_17_4 .C_ON=1'b0;
    defparam \FTDI.TXshift_7_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_7_LC_15_17_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \FTDI.TXshift_7_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__15422),
            .in2(_gnd_net_),
            .in3(N__11039),
            .lcout(\FTDI.TXshiftZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_7C_net ),
            .ce(N__12712),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNIV5TH_0_LC_16_8_0 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNIV5TH_0_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNIV5TH_0_LC_16_8_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \FTDI.RXstate_RNIV5TH_0_LC_16_8_0  (
            .in0(N__11510),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13951),
            .lcout(\FTDI.N_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNO_0_3_LC_16_8_1 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNO_0_3_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNO_0_3_LC_16_8_1 .LUT_INIT=16'b0101000011110001;
    LogicCell40 \FTDI.RXstate_RNO_0_3_LC_16_8_1  (
            .in0(N__11451),
            .in1(N__11023),
            .in2(N__11495),
            .in3(N__11417),
            .lcout(),
            .ltout(\FTDI.m13_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_3_LC_16_8_2 .C_ON=1'b0;
    defparam \FTDI.RXstate_3_LC_16_8_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_3_LC_16_8_2 .LUT_INIT=16'b1111011101010000;
    LogicCell40 \FTDI.RXstate_3_LC_16_8_2  (
            .in0(N__11511),
            .in1(N__13956),
            .in2(N__11000),
            .in3(N__11490),
            .lcout(\FTDI.RXstateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXstate_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_1_LC_16_8_3 .C_ON=1'b0;
    defparam \FTDI.RXstate_1_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_1_LC_16_8_3 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \FTDI.RXstate_1_LC_16_8_3  (
            .in0(N__11489),
            .in1(N__11418),
            .in2(N__13958),
            .in3(N__11513),
            .lcout(\FTDI.RXstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXstate_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_RNI29TH_2_LC_16_8_4 .C_ON=1'b0;
    defparam \FTDI.gap_RNI29TH_2_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \FTDI.gap_RNI29TH_2_LC_16_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FTDI.gap_RNI29TH_2_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__13952),
            .in2(_gnd_net_),
            .in3(N__11488),
            .lcout(\FTDI.N_201_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNI67DS1_0_LC_16_8_5 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNI67DS1_0_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNI67DS1_0_LC_16_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \FTDI.RXstate_RNI67DS1_0_LC_16_8_5  (
            .in0(N__11449),
            .in1(N__11415),
            .in2(N__11494),
            .in3(N__11509),
            .lcout(\FTDI.gap8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNO_0_0_LC_16_8_6 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNO_0_0_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNO_0_0_LC_16_8_6 .LUT_INIT=16'b0111000011111110;
    LogicCell40 \FTDI.RXstate_RNO_0_0_LC_16_8_6  (
            .in0(N__11416),
            .in1(N__11450),
            .in2(N__13957),
            .in3(N__11484),
            .lcout(),
            .ltout(\FTDI.N_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_0_LC_16_8_7 .C_ON=1'b0;
    defparam \FTDI.RXstate_0_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_0_LC_16_8_7 .LUT_INIT=16'b0000111110001000;
    LogicCell40 \FTDI.RXstate_0_LC_16_8_7  (
            .in0(N__11491),
            .in1(N__13950),
            .in2(N__11516),
            .in3(N__11512),
            .lcout(\FTDI.RXstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXstate_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_2_LC_16_9_1 .C_ON=1'b0;
    defparam \FTDI.RXstate_2_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_2_LC_16_9_1 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \FTDI.RXstate_2_LC_16_9_1  (
            .in0(N__11420),
            .in1(N__11431),
            .in2(N__11456),
            .in3(N__11493),
            .lcout(\FTDI.RXstateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXstate_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXready_LC_16_9_4 .C_ON=1'b0;
    defparam \FTDI.RXready_LC_16_9_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXready_LC_16_9_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \FTDI.RXready_LC_16_9_4  (
            .in0(N__11492),
            .in1(N__11452),
            .in2(N__11432),
            .in3(N__11419),
            .lcout(RXready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXstate_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXready_RNIICV7_1_LC_16_9_6 .C_ON=1'b0;
    defparam \FTDI.RXready_RNIICV7_1_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXready_RNIICV7_1_LC_16_9_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \FTDI.RXready_RNIICV7_1_LC_16_9_6  (
            .in0(N__15605),
            .in1(N__15881),
            .in2(N__15783),
            .in3(N__15498),
            .lcout(RXready_RNIICV7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXready_RNIICV7_0_LC_16_10_0 .C_ON=1'b0;
    defparam \FTDI.RXready_RNIICV7_0_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXready_RNIICV7_0_LC_16_10_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \FTDI.RXready_RNIICV7_0_LC_16_10_0  (
            .in0(N__15584),
            .in1(N__15880),
            .in2(N__15782),
            .in3(N__15499),
            .lcout(RXready_RNIICV7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam op_1_LC_16_10_3.C_ON=1'b0;
    defparam op_1_LC_16_10_3.SEQ_MODE=4'b1000;
    defparam op_1_LC_16_10_3.LUT_INIT=16'b1101111110000000;
    LogicCell40 op_1_LC_16_10_3 (
            .in0(N__15500),
            .in1(N__11321),
            .in2(N__15962),
            .in3(N__11203),
            .lcout(opZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.res_4_LC_16_10_6 .C_ON=1'b0;
    defparam \ALU.res_4_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \ALU.res_4_LC_16_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.res_4_LC_16_10_6  (
            .in0(N__11202),
            .in1(N__11174),
            .in2(_gnd_net_),
            .in3(N__11159),
            .lcout(res_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_ma_LC_16_11_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_ma_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_ma_LC_16_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_ma_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__14603),
            .in2(_gnd_net_),
            .in3(N__11940),
            .lcout(\ALU.regsA_result_cry_2_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_13_LC_16_11_3.C_ON=1'b0;
    defparam a_13_LC_16_11_3.SEQ_MODE=4'b1000;
    defparam a_13_LC_16_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_13_LC_16_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12281),
            .lcout(aZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16079),
            .ce(N__12213),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_ma_LC_16_11_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_ma_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_ma_LC_16_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_ma_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__11729),
            .in2(_gnd_net_),
            .in3(N__14740),
            .lcout(\ALU.regsA_result_cry_1_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_ma_LC_16_11_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_ma_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_ma_LC_16_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_ma_LC_16_11_6  (
            .in0(N__11730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15099),
            .lcout(\ALU.regsA_result_cry_3_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_ma_LC_16_11_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_ma_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_ma_LC_16_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_ma_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__13264),
            .in2(_gnd_net_),
            .in3(N__14741),
            .lcout(\ALU.regsA_result_cry_2_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_7_LC_16_12_1.C_ON=1'b0;
    defparam a_7_LC_16_12_1.SEQ_MODE=4'b1000;
    defparam a_7_LC_16_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_7_LC_16_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12114),
            .lcout(aZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16082),
            .ce(N__15274),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_ma_LC_16_12_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_ma_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_ma_LC_16_12_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_ma_LC_16_12_3  (
            .in0(N__11969),
            .in1(N__12926),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_2_ma_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_ma_LC_16_12_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_ma_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_ma_LC_16_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_ma_LC_16_12_4  (
            .in0(N__12927),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11783),
            .lcout(\ALU.regsA_result_cry_3_ma_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_ma_LC_16_12_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_ma_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_ma_LC_16_12_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_ma_LC_16_12_5  (
            .in0(N__13299),
            .in1(N__12928),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_4_ma_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_ma_LC_16_12_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_ma_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_ma_LC_16_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_ma_LC_16_12_6  (
            .in0(N__12929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11650),
            .lcout(\ALU.regsA_result_cry_5_ma_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_ma_LC_16_12_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_ma_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_ma_LC_16_12_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_ma_LC_16_12_7  (
            .in0(N__15005),
            .in1(N__12930),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_6_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_8_l_ofx_LC_16_13_0 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_8_l_ofx_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_8_l_ofx_LC_16_13_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_8_l_ofx_LC_16_13_0  (
            .in0(N__13152),
            .in1(N__14753),
            .in2(N__12653),
            .in3(N__12370),
            .lcout(\ALU.regsA_result_axb_8_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_8_LC_16_13_1.C_ON=1'b0;
    defparam b_8_LC_16_13_1.SEQ_MODE=4'b1000;
    defparam b_8_LC_16_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_8_LC_16_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14516),
            .lcout(bZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16087),
            .ce(N__14219),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_ma_LC_16_13_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_ma_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_ma_LC_16_13_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_ma_LC_16_13_2  (
            .in0(N__13148),
            .in1(N__14752),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_7_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_8_l_ofx_LC_16_13_3 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_8_l_ofx_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_8_l_ofx_LC_16_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_8_l_ofx_LC_16_13_3  (
            .in0(N__13515),
            .in1(N__12456),
            .in2(N__12857),
            .in3(N__13149),
            .lcout(\ALU.regsA_result_axb_8_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_ma_LC_16_13_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_ma_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_ma_LC_16_13_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_ma_LC_16_13_4  (
            .in0(N__13151),
            .in1(N__13514),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_9_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_9_l_ofx_LC_16_13_5 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_9_l_ofx_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_9_l_ofx_LC_16_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_9_l_ofx_LC_16_13_5  (
            .in0(N__13155),
            .in1(N__12457),
            .in2(N__13535),
            .in3(N__12368),
            .lcout(\ALU.regsA_result_axb_9_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_8_l_ofx_LC_16_13_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_8_l_ofx_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_8_l_ofx_LC_16_13_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_8_l_ofx_LC_16_13_6  (
            .in0(N__13150),
            .in1(N__12934),
            .in2(N__13878),
            .in3(N__12856),
            .lcout(\ALU.regsA_result_axb_8_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_9_l_ofx_LC_16_13_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_9_l_ofx_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_9_l_ofx_LC_16_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_9_l_ofx_LC_16_13_7  (
            .in0(N__13156),
            .in1(N__12369),
            .in2(N__12961),
            .in3(N__13863),
            .lcout(\ALU.regsA_result_axb_9_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_6_l_ofx_LC_16_14_1 .C_ON=1'b0;
    defparam \ALU.addsub_axb_6_l_ofx_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_6_l_ofx_LC_16_14_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.addsub_axb_6_l_ofx_LC_16_14_1  (
            .in0(N__13080),
            .in1(_gnd_net_),
            .in2(N__13880),
            .in3(N__14372),
            .lcout(\ALU.addsub_axb_6_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNO_LC_16_14_2 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNO_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNO_LC_16_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNO_LC_16_14_2  (
            .in0(N__13913),
            .in1(N__13874),
            .in2(_gnd_net_),
            .in3(N__13748),
            .lcout(\ALU.regsA_result_cry_2_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_3_l_ofx_LC_16_14_3 .C_ON=1'b0;
    defparam \ALU.addsub_axb_3_l_ofx_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_3_l_ofx_LC_16_14_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.addsub_axb_3_l_ofx_LC_16_14_3  (
            .in0(N__14371),
            .in1(N__13520),
            .in2(_gnd_net_),
            .in3(N__13338),
            .lcout(\ALU.addsub_axb_3_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_9_ma_LC_16_14_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_9_ma_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_9_ma_LC_16_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_9_ma_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__13154),
            .in2(_gnd_net_),
            .in3(N__12951),
            .lcout(\ALU.regsA_result_cry_9_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_ma_LC_16_14_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_ma_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_ma_LC_16_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_ma_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__12949),
            .in2(_gnd_net_),
            .in3(N__13079),
            .lcout(\ALU.regsA_result_cry_7_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_ma_LC_16_14_7 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_ma_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_ma_LC_16_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_ma_LC_16_14_7  (
            .in0(N__12950),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12830),
            .lcout(\ALU.regsA_result_cry_8_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_RNID8HD2_2_LC_16_15_0 .C_ON=1'b0;
    defparam \FTDI.baudAcc_RNID8HD2_2_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.baudAcc_RNID8HD2_2_LC_16_15_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \FTDI.baudAcc_RNID8HD2_2_LC_16_15_0  (
            .in0(N__16186),
            .in1(N__12752),
            .in2(N__15435),
            .in3(N__12682),
            .lcout(\FTDI.un1_TXstate_0_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXstart_esr_LC_16_15_1.C_ON=1'b0;
    defparam TXstart_esr_LC_16_15_1.SEQ_MODE=4'b1000;
    defparam TXstart_esr_LC_16_15_1.LUT_INIT=16'b1100100000000000;
    LogicCell40 TXstart_esr_LC_16_15_1 (
            .in0(N__15849),
            .in1(N__15768),
            .in2(N__15650),
            .in3(N__16185),
            .lcout(TXstartZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16098),
            .ce(N__12671),
            .sr(N__15961));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_ma_LC_16_15_6 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_ma_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_ma_LC_16_15_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_ma_LC_16_15_6  (
            .in0(N__14112),
            .in1(N__14821),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.regsA_result_cry_9_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_16_16_2 .C_ON=1'b0;
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_16_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \FTDI.un3_TX_cry_2_c_inv_LC_16_16_2  (
            .in0(N__14063),
            .in1(N__15454),
            .in2(_gnd_net_),
            .in3(N__14027),
            .lcout(\FTDI.un3_TX_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_1_LC_17_8_1 .C_ON=1'b0;
    defparam \FTDI.gap_1_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.gap_1_LC_17_8_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \FTDI.gap_1_LC_17_8_1  (
            .in0(N__13981),
            .in1(N__13969),
            .in2(_gnd_net_),
            .in3(N__13993),
            .lcout(\FTDI.gapZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_0_LC_17_8_3 .C_ON=1'b0;
    defparam \FTDI.gap_0_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.gap_0_LC_17_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \FTDI.gap_0_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__13968),
            .in2(_gnd_net_),
            .in3(N__13992),
            .lcout(\FTDI.gapZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_2_LC_17_8_6 .C_ON=1'b0;
    defparam \FTDI.gap_2_LC_17_8_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.gap_2_LC_17_8_6 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \FTDI.gap_2_LC_17_8_6  (
            .in0(N__13994),
            .in1(N__13982),
            .in2(N__13973),
            .in3(_gnd_net_),
            .lcout(\FTDI.gapZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXready_RNIICV7_LC_17_9_3 .C_ON=1'b0;
    defparam \FTDI.RXready_RNIICV7_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXready_RNIICV7_LC_17_9_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \FTDI.RXready_RNIICV7_LC_17_9_3  (
            .in0(N__15606),
            .in1(N__15882),
            .in2(N__15784),
            .in3(N__15501),
            .lcout(RXready_RNIICV7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_10_2_0__m7_x1_LC_17_11_1.C_ON=1'b0;
    defparam testState_10_2_0__m7_x1_LC_17_11_1.SEQ_MODE=4'b0000;
    defparam testState_10_2_0__m7_x1_LC_17_11_1.LUT_INIT=16'b0110011001101010;
    LogicCell40 testState_10_2_0__m7_x1_LC_17_11_1 (
            .in0(N__15573),
            .in1(N__15853),
            .in2(N__15760),
            .in3(N__15502),
            .lcout(m7_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXready_RNIICV7_2_LC_17_11_4 .C_ON=1'b0;
    defparam \FTDI.RXready_RNIICV7_2_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXready_RNIICV7_2_LC_17_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \FTDI.RXready_RNIICV7_2_LC_17_11_4  (
            .in0(N__15504),
            .in1(N__15735),
            .in2(N__15879),
            .in3(N__15572),
            .lcout(RXready_RNIICV7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_10_2_0__m7_x0_LC_17_11_5.C_ON=1'b0;
    defparam testState_10_2_0__m7_x0_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam testState_10_2_0__m7_x0_LC_17_11_5.LUT_INIT=16'b1010011010101010;
    LogicCell40 testState_10_2_0__m7_x0_LC_17_11_5 (
            .in0(N__15574),
            .in1(N__15854),
            .in2(N__15761),
            .in3(N__15503),
            .lcout(),
            .ltout(m7_x0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_1_LC_17_11_6.C_ON=1'b0;
    defparam testState_1_LC_17_11_6.SEQ_MODE=4'b1000;
    defparam testState_1_LC_17_11_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 testState_1_LC_17_11_6 (
            .in0(_gnd_net_),
            .in1(N__15305),
            .in2(N__15299),
            .in3(N__16196),
            .lcout(testStateZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16086),
            .ce(),
            .sr(_gnd_net_));
    defparam a_0_LC_17_12_0.C_ON=1'b0;
    defparam a_0_LC_17_12_0.SEQ_MODE=4'b1000;
    defparam a_0_LC_17_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 a_0_LC_17_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14510),
            .lcout(aZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16093),
            .ce(N__15273),
            .sr(_gnd_net_));
    defparam testState_RNIJBO_1_LC_17_13_0.C_ON=1'b0;
    defparam testState_RNIJBO_1_LC_17_13_0.SEQ_MODE=4'b0000;
    defparam testState_RNIJBO_1_LC_17_13_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 testState_RNIJBO_1_LC_17_13_0 (
            .in0(_gnd_net_),
            .in1(N__15601),
            .in2(_gnd_net_),
            .in3(N__15872),
            .lcout(),
            .ltout(testState30_testState30_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_2_LC_17_13_1.C_ON=1'b0;
    defparam testState_2_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam testState_2_LC_17_13_1.LUT_INIT=16'b0100101011101010;
    LogicCell40 testState_2_LC_17_13_1 (
            .in0(N__15731),
            .in1(N__15518),
            .in2(N__15209),
            .in3(N__16195),
            .lcout(testStateZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16097),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_5_l_ofx_LC_17_13_3 .C_ON=1'b0;
    defparam \ALU.addsub_axb_5_l_ofx_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_5_l_ofx_LC_17_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_5_l_ofx_LC_17_13_3  (
            .in0(N__15191),
            .in1(N__14368),
            .in2(_gnd_net_),
            .in3(N__15036),
            .lcout(\ALU.addsub_axb_5_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_ma_LC_17_13_4 .C_ON=1'b0;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_ma_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_ma_LC_17_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_ma_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__14243),
            .in2(_gnd_net_),
            .in3(N__14754),
            .lcout(\ALU.regsA_result_cry_13_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_axb_13_l_ofx_LC_17_13_5 .C_ON=1'b0;
    defparam \ALU.addsub_axb_13_l_ofx_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_axb_13_l_ofx_LC_17_13_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.addsub_axb_13_l_ofx_LC_17_13_5  (
            .in0(N__14622),
            .in1(N__14579),
            .in2(_gnd_net_),
            .in3(N__14369),
            .lcout(\ALU.addsub_axb_13_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam op_0_LC_17_13_7.C_ON=1'b0;
    defparam op_0_LC_17_13_7.SEQ_MODE=4'b1000;
    defparam op_0_LC_17_13_7.LUT_INIT=16'b1111011110000000;
    LogicCell40 op_0_LC_17_13_7 (
            .in0(N__15954),
            .in1(N__15517),
            .in2(N__14515),
            .in3(N__14370),
            .lcout(opZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16097),
            .ce(),
            .sr(_gnd_net_));
    defparam b_14_LC_17_14_2.C_ON=1'b0;
    defparam b_14_LC_17_14_2.SEQ_MODE=4'b1000;
    defparam b_14_LC_17_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 b_14_LC_17_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14317),
            .lcout(bZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16103),
            .ce(N__14215),
            .sr(_gnd_net_));
    defparam testState_10_2_0__i3_mux_i_x0_LC_17_15_1.C_ON=1'b0;
    defparam testState_10_2_0__i3_mux_i_x0_LC_17_15_1.SEQ_MODE=4'b0000;
    defparam testState_10_2_0__i3_mux_i_x0_LC_17_15_1.LUT_INIT=16'b1001110110101010;
    LogicCell40 testState_10_2_0__i3_mux_i_x0_LC_17_15_1 (
            .in0(N__15828),
            .in1(N__15734),
            .in2(N__15646),
            .in3(N__15516),
            .lcout(),
            .ltout(i3_mux_i_x0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_0_LC_17_15_2.C_ON=1'b0;
    defparam testState_0_LC_17_15_2.SEQ_MODE=4'b1000;
    defparam testState_0_LC_17_15_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 testState_0_LC_17_15_2 (
            .in0(_gnd_net_),
            .in1(N__15461),
            .in2(N__16199),
            .in3(N__16187),
            .lcout(testStateZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16106),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_RNIUI41_2_LC_17_15_6.C_ON=1'b0;
    defparam testState_RNIUI41_2_LC_17_15_6.SEQ_MODE=4'b0000;
    defparam testState_RNIUI41_2_LC_17_15_6.LUT_INIT=16'b0000000000010001;
    LogicCell40 testState_RNIUI41_2_LC_17_15_6 (
            .in0(N__15732),
            .in1(N__15612),
            .in2(_gnd_net_),
            .in3(N__15826),
            .lcout(testState27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_10_2_0__i3_mux_i_x1_LC_17_15_7.C_ON=1'b0;
    defparam testState_10_2_0__i3_mux_i_x1_LC_17_15_7.SEQ_MODE=4'b0000;
    defparam testState_10_2_0__i3_mux_i_x1_LC_17_15_7.LUT_INIT=16'b0101010101100010;
    LogicCell40 testState_10_2_0__i3_mux_i_x1_LC_17_15_7 (
            .in0(N__15827),
            .in1(N__15733),
            .in2(N__15645),
            .in3(N__15515),
            .lcout(i3_mux_i_x1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_2_c_LC_17_16_0 .C_ON=1'b1;
    defparam \FTDI.un3_TX_cry_2_c_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_2_c_LC_17_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \FTDI.un3_TX_cry_2_c_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__15455),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\FTDI.un3_TX_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_17_16_1 .C_ON=1'b1;
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_17_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \FTDI.un3_TX_cry_3_c_inv_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__15443),
            .in2(_gnd_net_),
            .in3(N__15437),
            .lcout(\FTDI.un3_TX_axb_3 ),
            .ltout(),
            .carryin(\FTDI.un3_TX_cry_2 ),
            .carryout(\FTDI.un3_TX_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_17_16_2 .C_ON=1'b0;
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_17_16_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_17_16_2  (
            .in0(N__15436),
            .in1(N__15341),
            .in2(_gnd_net_),
            .in3(N__15329),
            .lcout(FTDI_TX_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
