
module gpu(
    output reg [7:0] red,
    output reg [7:0] green,
    output reg [7:0] blue,

    input wire [7:0] address,
    
  );

endmodule
