module promdata(
    input wire CLK,
    input wire [15:0] address,
    output wire [31:0] data
  );

  // Xilinx style block ram directive
  (* rom_style = "block" *) reg [31:0] dintern = 32'b0;

  always @( * ) begin
    case (address)
      16'h0000: dintern = 32'h00000007;
      16'h0001: dintern = 32'h04000008;
      16'h0002: dintern = 32'h04010008;
      16'h0003: dintern = 32'h20100007;
      16'h0004: dintern = 32'h04020008;
      16'h0005: dintern = 32'h00840054;
      16'h0006: dintern = 32'h00110054;
      16'h0007: dintern = 32'h00160054;
      16'h0008: dintern = 32'h001A0054;
      16'h0009: dintern = 32'h028AC007;
      16'h000A: dintern = 32'h0C20E007;
      16'h000B: dintern = 32'h00038007;
      16'h000C: dintern = 32'h0000A007;
      16'h000D: dintern = 32'h003D0054;
      16'h000E: dintern = 32'h006D0054;
      16'h000F: dintern = 32'h00060050;
      16'h0010: dintern = 32'h00100050;
      16'h0011: dintern = 32'hFFFFE007;
      16'h0012: dintern = 32'h0000000E;
      16'h0013: dintern = 32'h00010017;
      16'h0014: dintern = 32'h00000464;
      16'h0015: dintern = 32'h00110050;
      16'h0016: dintern = 32'hFFFFE007;
      16'h0017: dintern = 32'h0000C007;
      16'h0018: dintern = 32'h00000311;
      16'h0019: dintern = 32'h00000058;
      16'h001A: dintern = 32'h04000004;
      16'h001B: dintern = 32'h0001001B;
      16'h001C: dintern = 32'h04000008;
      16'h001D: dintern = 32'h00010017;
      16'h001E: dintern = 32'h00001064;
      16'h001F: dintern = 32'h00000007;
      16'h0020: dintern = 32'h04000008;
      16'h0021: dintern = 32'h00000058;
      16'h0022: dintern = 32'h0003C323;
      16'h0023: dintern = 32'h0000C31B;
      16'h0024: dintern = 32'h0000000D;
      16'h0025: dintern = 32'h00004007;
      16'h0026: dintern = 32'h00006007;
      16'h0027: dintern = 32'h00060117;
      16'h0028: dintern = 32'h0034045C;
      16'h0029: dintern = 32'h0001411B;
      16'h002A: dintern = 32'h0001202F;
      16'h002B: dintern = 32'h00010043;
      16'h002C: dintern = 32'h00000097;
      16'h002D: dintern = 32'h0031045C;
      16'h002E: dintern = 32'h00000211;
      16'h002F: dintern = 32'h0100E39B;
      16'h0030: dintern = 32'h00270050;
      16'h0031: dintern = 32'h00000291;
      16'h0032: dintern = 32'h0100E39B;
      16'h0033: dintern = 32'h00270050;
      16'h0034: dintern = 32'h00020197;
      16'h0035: dintern = 32'h00000464;
      16'h0036: dintern = 32'h0001619B;
      16'h0037: dintern = 32'h0001C31B;
      16'h0038: dintern = 32'h0000000D;
      16'h0039: dintern = 32'h00004007;
      16'h003A: dintern = 32'h0001E39B;
      16'h003B: dintern = 32'h0600E39F;
      16'h003C: dintern = 32'h00270050;
      16'h003D: dintern = 32'h04030308;
      16'h003E: dintern = 32'h0000000D;
      16'h003F: dintern = 32'h00000017;
      16'h0040: dintern = 32'h00000464;
      16'h0041: dintern = 32'h0000C01B;
      16'h0042: dintern = 32'h00220054;
      16'h0043: dintern = 32'h0002E39B;
      16'h0044: dintern = 32'h0600E39F;
      16'h0045: dintern = 32'h0403C004;
      16'h0046: dintern = 32'h0001C31B;
      16'h0047: dintern = 32'h003D0050;
      16'h0048: dintern = 32'h04050288;
      16'h0049: dintern = 32'h04040208;
      16'h004A: dintern = 32'h00004007;
      16'h004B: dintern = 32'h00006007;
      16'h004C: dintern = 32'h0000000D;
      16'h004D: dintern = 32'h04048004;
      16'h004E: dintern = 32'h00FF822F;
      16'h004F: dintern = 32'h00001115;
      16'h0050: dintern = 32'h0061045C;
      16'h0051: dintern = 32'h0001202F;
      16'h0052: dintern = 32'h005A00DC;
      16'h0053: dintern = 32'h0405A004;
      16'h0054: dintern = 32'h00FFA2AF;
      16'h0055: dintern = 32'h00000291;
      16'h0056: dintern = 32'h0100E39B;
      16'h0057: dintern = 32'h0001411B;
      16'h0058: dintern = 32'h00010043;
      16'h0059: dintern = 32'h004D0050;
      16'h005A: dintern = 32'h0405A004;
      16'h005B: dintern = 32'h0008A2C3;
      16'h005C: dintern = 32'h00000291;
      16'h005D: dintern = 32'h0100E39B;
      16'h005E: dintern = 32'h0001411B;
      16'h005F: dintern = 32'h00010043;
      16'h0060: dintern = 32'h004D0050;
      16'h0061: dintern = 32'h04048004;
      16'h0062: dintern = 32'h00088243;
      16'h0063: dintern = 32'h00001195;
      16'h0064: dintern = 32'h00000464;
      16'h0065: dintern = 32'h0001619B;
      16'h0066: dintern = 32'h01004123;
      16'h0067: dintern = 32'h0000EB9D;
      16'h0068: dintern = 32'h0001C31B;
      16'h0069: dintern = 32'h0000000D;
      16'h006A: dintern = 32'h0001E39B;
      16'h006B: dintern = 32'h00004007;
      16'h006C: dintern = 32'h004D0050;
      16'h006D: dintern = 32'h04000004;
      16'h006E: dintern = 32'h00000017;
      16'h006F: dintern = 32'h0071045C;
      16'h0070: dintern = 32'h00000058;
      16'h0071: dintern = 32'h10108007;
      16'h0072: dintern = 32'h0004A007;
      16'h0073: dintern = 32'h0401C004;
      16'h0074: dintern = 32'h0010C323;
      16'h0075: dintern = 32'h0180C31B;
      16'h0076: dintern = 32'h0402E004;
      16'h0077: dintern = 32'h00480054;
      16'h0078: dintern = 32'h04020004;
      16'h0079: dintern = 32'h0002001B;
      16'h007A: dintern = 32'h04020008;
      16'h007B: dintern = 32'h04010004;
      16'h007C: dintern = 32'h0001001B;
      16'h007D: dintern = 32'h000E0017;
      16'h007E: dintern = 32'h0081045C;
      16'h007F: dintern = 32'h04010008;
      16'h0080: dintern = 32'h00000058;
      16'h0081: dintern = 32'h00000007;
      16'h0082: dintern = 32'h04010008;
      16'h0083: dintern = 32'h00000058;
      16'h0084: dintern = 32'h0280C007;
      16'h0085: dintern = 32'h9900E007;
      16'h0086: dintern = 32'h00002007;
      16'h0087: dintern = 32'h000A0097;
      16'h0088: dintern = 32'h00000464;
      16'h0089: dintern = 32'h0001209B;
      16'h008A: dintern = 32'h0000000D;
      16'h008B: dintern = 32'h00000011;
      16'h008C: dintern = 32'h0001C31B;
      16'h008D: dintern = 32'h0001E39B;
      16'h008E: dintern = 32'h00870050;
      default: dintern = 32'h0;
    endcase
  end

  assign data = dintern;

endmodule
