module promdata(
    input wire CLK,
    input wire [15:0] address,
    output wire [31:0] data
  );

  // Xilinx style block ram directive
  (* rom_style = "block" *) reg [31:0] dintern = 32'b0;

  always @( * ) begin
    case (address)
      16'h0000: dintern = 32'h00080007;
      16'h0001: dintern = 32'h04000008;
      16'h0002: dintern = 32'h00002005;
      16'h0003: dintern = 32'h00004007;
      16'h0004: dintern = 32'h00000419;
      16'h0005: dintern = 32'h0000043D;
      16'h0006: dintern = 32'h00080017;
      16'h0007: dintern = 32'h0009085C;
      16'h0008: dintern = 32'h00080050;
      16'h0009: dintern = 32'h00030008;
      16'h000A: dintern = 32'h00080043;
      16'h000B: dintern = 32'h00030008;
      16'h000C: dintern = 32'h00080050;
      default: dintern = 32'h0;
    endcase
  end

  assign data = dintern;

endmodule
