-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Aug 15 2020 12:51:42

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    TX : out std_logic;
    GPIO11 : out std_logic;
    CLK : in std_logic;
    RX : in std_logic;
    GPIO9 : out std_logic;
    GPIO3 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__57007\ : std_logic;
signal \N__57006\ : std_logic;
signal \N__57005\ : std_logic;
signal \N__56996\ : std_logic;
signal \N__56995\ : std_logic;
signal \N__56994\ : std_logic;
signal \N__56987\ : std_logic;
signal \N__56986\ : std_logic;
signal \N__56985\ : std_logic;
signal \N__56978\ : std_logic;
signal \N__56977\ : std_logic;
signal \N__56976\ : std_logic;
signal \N__56969\ : std_logic;
signal \N__56968\ : std_logic;
signal \N__56967\ : std_logic;
signal \N__56950\ : std_logic;
signal \N__56949\ : std_logic;
signal \N__56948\ : std_logic;
signal \N__56947\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56945\ : std_logic;
signal \N__56942\ : std_logic;
signal \N__56937\ : std_logic;
signal \N__56932\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56920\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56908\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56900\ : std_logic;
signal \N__56897\ : std_logic;
signal \N__56896\ : std_logic;
signal \N__56895\ : std_logic;
signal \N__56894\ : std_logic;
signal \N__56891\ : std_logic;
signal \N__56888\ : std_logic;
signal \N__56885\ : std_logic;
signal \N__56882\ : std_logic;
signal \N__56877\ : std_logic;
signal \N__56866\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56864\ : std_logic;
signal \N__56863\ : std_logic;
signal \N__56862\ : std_logic;
signal \N__56861\ : std_logic;
signal \N__56858\ : std_logic;
signal \N__56851\ : std_logic;
signal \N__56846\ : std_logic;
signal \N__56839\ : std_logic;
signal \N__56838\ : std_logic;
signal \N__56837\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56835\ : std_logic;
signal \N__56834\ : std_logic;
signal \N__56833\ : std_logic;
signal \N__56832\ : std_logic;
signal \N__56831\ : std_logic;
signal \N__56826\ : std_logic;
signal \N__56817\ : std_logic;
signal \N__56816\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56810\ : std_logic;
signal \N__56807\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56801\ : std_logic;
signal \N__56800\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56798\ : std_logic;
signal \N__56797\ : std_logic;
signal \N__56796\ : std_logic;
signal \N__56795\ : std_logic;
signal \N__56792\ : std_logic;
signal \N__56789\ : std_logic;
signal \N__56786\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56773\ : std_logic;
signal \N__56768\ : std_logic;
signal \N__56763\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56741\ : std_logic;
signal \N__56740\ : std_logic;
signal \N__56739\ : std_logic;
signal \N__56738\ : std_logic;
signal \N__56737\ : std_logic;
signal \N__56732\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56720\ : std_logic;
signal \N__56713\ : std_logic;
signal \N__56710\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56704\ : std_logic;
signal \N__56703\ : std_logic;
signal \N__56702\ : std_logic;
signal \N__56701\ : std_logic;
signal \N__56696\ : std_logic;
signal \N__56695\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56689\ : std_logic;
signal \N__56686\ : std_logic;
signal \N__56681\ : std_logic;
signal \N__56674\ : std_logic;
signal \N__56673\ : std_logic;
signal \N__56670\ : std_logic;
signal \N__56669\ : std_logic;
signal \N__56666\ : std_logic;
signal \N__56661\ : std_logic;
signal \N__56656\ : std_logic;
signal \N__56655\ : std_logic;
signal \N__56652\ : std_logic;
signal \N__56649\ : std_logic;
signal \N__56644\ : std_logic;
signal \N__56641\ : std_logic;
signal \N__56640\ : std_logic;
signal \N__56635\ : std_logic;
signal \N__56632\ : std_logic;
signal \N__56629\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56623\ : std_logic;
signal \N__56620\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56614\ : std_logic;
signal \N__56611\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56605\ : std_logic;
signal \N__56602\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56596\ : std_logic;
signal \N__56593\ : std_logic;
signal \N__56590\ : std_logic;
signal \N__56587\ : std_logic;
signal \N__56586\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56580\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56573\ : std_logic;
signal \N__56570\ : std_logic;
signal \N__56567\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56558\ : std_logic;
signal \N__56555\ : std_logic;
signal \N__56550\ : std_logic;
signal \N__56545\ : std_logic;
signal \N__56542\ : std_logic;
signal \N__56539\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56533\ : std_logic;
signal \N__56530\ : std_logic;
signal \N__56527\ : std_logic;
signal \N__56524\ : std_logic;
signal \N__56521\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56507\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56505\ : std_logic;
signal \N__56504\ : std_logic;
signal \N__56501\ : std_logic;
signal \N__56498\ : std_logic;
signal \N__56495\ : std_logic;
signal \N__56492\ : std_logic;
signal \N__56489\ : std_logic;
signal \N__56488\ : std_logic;
signal \N__56485\ : std_logic;
signal \N__56482\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56477\ : std_logic;
signal \N__56476\ : std_logic;
signal \N__56475\ : std_logic;
signal \N__56472\ : std_logic;
signal \N__56469\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56463\ : std_logic;
signal \N__56460\ : std_logic;
signal \N__56457\ : std_logic;
signal \N__56454\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56448\ : std_logic;
signal \N__56445\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56437\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56431\ : std_logic;
signal \N__56426\ : std_logic;
signal \N__56423\ : std_logic;
signal \N__56420\ : std_logic;
signal \N__56417\ : std_logic;
signal \N__56414\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56399\ : std_logic;
signal \N__56398\ : std_logic;
signal \N__56397\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56389\ : std_logic;
signal \N__56386\ : std_logic;
signal \N__56381\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56375\ : std_logic;
signal \N__56372\ : std_logic;
signal \N__56369\ : std_logic;
signal \N__56366\ : std_logic;
signal \N__56363\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56351\ : std_logic;
signal \N__56348\ : std_logic;
signal \N__56343\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56331\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56319\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56311\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56303\ : std_logic;
signal \N__56302\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56300\ : std_logic;
signal \N__56299\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56296\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56294\ : std_logic;
signal \N__56293\ : std_logic;
signal \N__56292\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56290\ : std_logic;
signal \N__56289\ : std_logic;
signal \N__56288\ : std_logic;
signal \N__56287\ : std_logic;
signal \N__56286\ : std_logic;
signal \N__56285\ : std_logic;
signal \N__56284\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56282\ : std_logic;
signal \N__56281\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56277\ : std_logic;
signal \N__56276\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56274\ : std_logic;
signal \N__56273\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56270\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56267\ : std_logic;
signal \N__56266\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56264\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56262\ : std_logic;
signal \N__56261\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56258\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56255\ : std_logic;
signal \N__56254\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56252\ : std_logic;
signal \N__56251\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56249\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56246\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56243\ : std_logic;
signal \N__56242\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56240\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56238\ : std_logic;
signal \N__56237\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56235\ : std_logic;
signal \N__56234\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56232\ : std_logic;
signal \N__56231\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56226\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56058\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56055\ : std_logic;
signal \N__56054\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56052\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56049\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56046\ : std_logic;
signal \N__56045\ : std_logic;
signal \N__56044\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56042\ : std_logic;
signal \N__56041\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56039\ : std_logic;
signal \N__56038\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56036\ : std_logic;
signal \N__55987\ : std_logic;
signal \N__55984\ : std_logic;
signal \N__55981\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55972\ : std_logic;
signal \N__55969\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55962\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55958\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55955\ : std_logic;
signal \N__55952\ : std_logic;
signal \N__55951\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55947\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55942\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55939\ : std_logic;
signal \N__55934\ : std_logic;
signal \N__55933\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55930\ : std_logic;
signal \N__55929\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55927\ : std_logic;
signal \N__55924\ : std_logic;
signal \N__55921\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55910\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55904\ : std_logic;
signal \N__55903\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55896\ : std_logic;
signal \N__55893\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55879\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55871\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55861\ : std_logic;
signal \N__55858\ : std_logic;
signal \N__55853\ : std_logic;
signal \N__55848\ : std_logic;
signal \N__55847\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55841\ : std_logic;
signal \N__55840\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55834\ : std_logic;
signal \N__55831\ : std_logic;
signal \N__55826\ : std_logic;
signal \N__55819\ : std_logic;
signal \N__55818\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55814\ : std_logic;
signal \N__55809\ : std_logic;
signal \N__55808\ : std_logic;
signal \N__55807\ : std_logic;
signal \N__55806\ : std_logic;
signal \N__55805\ : std_logic;
signal \N__55802\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55799\ : std_logic;
signal \N__55798\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55784\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55776\ : std_logic;
signal \N__55773\ : std_logic;
signal \N__55772\ : std_logic;
signal \N__55769\ : std_logic;
signal \N__55766\ : std_logic;
signal \N__55763\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55759\ : std_logic;
signal \N__55754\ : std_logic;
signal \N__55749\ : std_logic;
signal \N__55744\ : std_logic;
signal \N__55741\ : std_logic;
signal \N__55738\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55736\ : std_logic;
signal \N__55731\ : std_logic;
signal \N__55730\ : std_logic;
signal \N__55729\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55723\ : std_logic;
signal \N__55722\ : std_logic;
signal \N__55719\ : std_logic;
signal \N__55716\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55701\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55693\ : std_logic;
signal \N__55690\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55679\ : std_logic;
signal \N__55676\ : std_logic;
signal \N__55671\ : std_logic;
signal \N__55666\ : std_logic;
signal \N__55663\ : std_logic;
signal \N__55660\ : std_logic;
signal \N__55659\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55642\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55640\ : std_logic;
signal \N__55631\ : std_logic;
signal \N__55626\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55609\ : std_logic;
signal \N__55604\ : std_logic;
signal \N__55601\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55586\ : std_logic;
signal \N__55585\ : std_logic;
signal \N__55582\ : std_logic;
signal \N__55579\ : std_logic;
signal \N__55574\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55555\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55536\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55533\ : std_logic;
signal \N__55530\ : std_logic;
signal \N__55529\ : std_logic;
signal \N__55528\ : std_logic;
signal \N__55527\ : std_logic;
signal \N__55524\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55521\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55517\ : std_logic;
signal \N__55514\ : std_logic;
signal \N__55513\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55507\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55503\ : std_logic;
signal \N__55500\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55491\ : std_logic;
signal \N__55490\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55488\ : std_logic;
signal \N__55485\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55481\ : std_logic;
signal \N__55480\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55476\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55468\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55458\ : std_logic;
signal \N__55449\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55446\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55434\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55428\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55417\ : std_logic;
signal \N__55414\ : std_logic;
signal \N__55411\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55401\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55388\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55381\ : std_logic;
signal \N__55378\ : std_logic;
signal \N__55375\ : std_logic;
signal \N__55366\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55348\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55342\ : std_logic;
signal \N__55337\ : std_logic;
signal \N__55334\ : std_logic;
signal \N__55331\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55325\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55316\ : std_logic;
signal \N__55311\ : std_logic;
signal \N__55306\ : std_logic;
signal \N__55303\ : std_logic;
signal \N__55282\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55279\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55269\ : std_logic;
signal \N__55268\ : std_logic;
signal \N__55265\ : std_logic;
signal \N__55264\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55262\ : std_logic;
signal \N__55261\ : std_logic;
signal \N__55260\ : std_logic;
signal \N__55259\ : std_logic;
signal \N__55256\ : std_logic;
signal \N__55253\ : std_logic;
signal \N__55250\ : std_logic;
signal \N__55247\ : std_logic;
signal \N__55244\ : std_logic;
signal \N__55241\ : std_logic;
signal \N__55238\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55227\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55216\ : std_logic;
signal \N__55205\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55199\ : std_logic;
signal \N__55196\ : std_logic;
signal \N__55193\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55189\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55176\ : std_logic;
signal \N__55173\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55153\ : std_logic;
signal \N__55150\ : std_logic;
signal \N__55143\ : std_logic;
signal \N__55142\ : std_logic;
signal \N__55139\ : std_logic;
signal \N__55138\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55130\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55114\ : std_logic;
signal \N__55111\ : std_logic;
signal \N__55108\ : std_logic;
signal \N__55105\ : std_logic;
signal \N__55102\ : std_logic;
signal \N__55099\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55072\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55062\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55048\ : std_logic;
signal \N__55045\ : std_logic;
signal \N__55042\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55030\ : std_logic;
signal \N__55027\ : std_logic;
signal \N__55024\ : std_logic;
signal \N__55021\ : std_logic;
signal \N__55018\ : std_logic;
signal \N__55015\ : std_logic;
signal \N__55008\ : std_logic;
signal \N__55003\ : std_logic;
signal \N__54998\ : std_logic;
signal \N__54991\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54972\ : std_logic;
signal \N__54969\ : std_logic;
signal \N__54966\ : std_logic;
signal \N__54961\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54957\ : std_logic;
signal \N__54956\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54940\ : std_logic;
signal \N__54937\ : std_logic;
signal \N__54936\ : std_logic;
signal \N__54933\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54923\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54921\ : std_logic;
signal \N__54920\ : std_logic;
signal \N__54919\ : std_logic;
signal \N__54916\ : std_logic;
signal \N__54915\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54907\ : std_logic;
signal \N__54906\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54902\ : std_logic;
signal \N__54901\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54899\ : std_logic;
signal \N__54898\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54891\ : std_logic;
signal \N__54890\ : std_logic;
signal \N__54889\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54887\ : std_logic;
signal \N__54886\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54878\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54864\ : std_logic;
signal \N__54861\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54858\ : std_logic;
signal \N__54855\ : std_logic;
signal \N__54850\ : std_logic;
signal \N__54843\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54834\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54830\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54824\ : std_logic;
signal \N__54823\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54821\ : std_logic;
signal \N__54818\ : std_logic;
signal \N__54817\ : std_logic;
signal \N__54814\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54812\ : std_logic;
signal \N__54811\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54805\ : std_logic;
signal \N__54804\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54802\ : std_logic;
signal \N__54801\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54797\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54795\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54791\ : std_logic;
signal \N__54790\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54788\ : std_logic;
signal \N__54787\ : std_logic;
signal \N__54786\ : std_logic;
signal \N__54785\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54783\ : std_logic;
signal \N__54782\ : std_logic;
signal \N__54781\ : std_logic;
signal \N__54780\ : std_logic;
signal \N__54779\ : std_logic;
signal \N__54778\ : std_logic;
signal \N__54777\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54765\ : std_logic;
signal \N__54760\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54749\ : std_logic;
signal \N__54746\ : std_logic;
signal \N__54739\ : std_logic;
signal \N__54734\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54725\ : std_logic;
signal \N__54720\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54715\ : std_logic;
signal \N__54708\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54701\ : std_logic;
signal \N__54698\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54681\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54664\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54658\ : std_logic;
signal \N__54655\ : std_logic;
signal \N__54652\ : std_logic;
signal \N__54651\ : std_logic;
signal \N__54648\ : std_logic;
signal \N__54645\ : std_logic;
signal \N__54642\ : std_logic;
signal \N__54641\ : std_logic;
signal \N__54640\ : std_logic;
signal \N__54639\ : std_logic;
signal \N__54638\ : std_logic;
signal \N__54633\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54630\ : std_logic;
signal \N__54629\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54627\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54622\ : std_logic;
signal \N__54619\ : std_logic;
signal \N__54618\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54616\ : std_logic;
signal \N__54615\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54608\ : std_logic;
signal \N__54607\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54605\ : std_logic;
signal \N__54604\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54597\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54595\ : std_logic;
signal \N__54594\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54592\ : std_logic;
signal \N__54591\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54587\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54584\ : std_logic;
signal \N__54583\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54577\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54563\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54557\ : std_logic;
signal \N__54556\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54554\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54552\ : std_logic;
signal \N__54547\ : std_logic;
signal \N__54540\ : std_logic;
signal \N__54533\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54521\ : std_logic;
signal \N__54520\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54496\ : std_logic;
signal \N__54489\ : std_logic;
signal \N__54484\ : std_logic;
signal \N__54479\ : std_logic;
signal \N__54478\ : std_logic;
signal \N__54475\ : std_logic;
signal \N__54470\ : std_logic;
signal \N__54467\ : std_logic;
signal \N__54464\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54448\ : std_logic;
signal \N__54447\ : std_logic;
signal \N__54442\ : std_logic;
signal \N__54439\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54429\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54409\ : std_logic;
signal \N__54406\ : std_logic;
signal \N__54403\ : std_logic;
signal \N__54396\ : std_logic;
signal \N__54393\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54383\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54365\ : std_logic;
signal \N__54362\ : std_logic;
signal \N__54359\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54349\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54325\ : std_logic;
signal \N__54322\ : std_logic;
signal \N__54319\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54301\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54295\ : std_logic;
signal \N__54290\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__54260\ : std_logic;
signal \N__54257\ : std_logic;
signal \N__54250\ : std_logic;
signal \N__54247\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54233\ : std_logic;
signal \N__54230\ : std_logic;
signal \N__54219\ : std_logic;
signal \N__54216\ : std_logic;
signal \N__54215\ : std_logic;
signal \N__54212\ : std_logic;
signal \N__54209\ : std_logic;
signal \N__54204\ : std_logic;
signal \N__54193\ : std_logic;
signal \N__54188\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54167\ : std_logic;
signal \N__54164\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54129\ : std_logic;
signal \N__54128\ : std_logic;
signal \N__54125\ : std_logic;
signal \N__54120\ : std_logic;
signal \N__54111\ : std_logic;
signal \N__54108\ : std_logic;
signal \N__54105\ : std_logic;
signal \N__54102\ : std_logic;
signal \N__54099\ : std_logic;
signal \N__54096\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54066\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54062\ : std_logic;
signal \N__54061\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54059\ : std_logic;
signal \N__54058\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54056\ : std_logic;
signal \N__54055\ : std_logic;
signal \N__54054\ : std_logic;
signal \N__54053\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54051\ : std_logic;
signal \N__54050\ : std_logic;
signal \N__54049\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54047\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54041\ : std_logic;
signal \N__54040\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54038\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54033\ : std_logic;
signal \N__54032\ : std_logic;
signal \N__54029\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54027\ : std_logic;
signal \N__54026\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54023\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54020\ : std_logic;
signal \N__54017\ : std_logic;
signal \N__54014\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54003\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__54000\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53985\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53975\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53973\ : std_logic;
signal \N__53972\ : std_logic;
signal \N__53971\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53959\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53955\ : std_logic;
signal \N__53952\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53950\ : std_logic;
signal \N__53949\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53946\ : std_logic;
signal \N__53945\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53930\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53928\ : std_logic;
signal \N__53927\ : std_logic;
signal \N__53926\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53923\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53914\ : std_logic;
signal \N__53913\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53901\ : std_logic;
signal \N__53900\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53897\ : std_logic;
signal \N__53896\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53893\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53887\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53873\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53864\ : std_logic;
signal \N__53861\ : std_logic;
signal \N__53858\ : std_logic;
signal \N__53857\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53826\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53804\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53781\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53759\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53748\ : std_logic;
signal \N__53743\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53732\ : std_logic;
signal \N__53725\ : std_logic;
signal \N__53718\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53702\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53687\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53681\ : std_logic;
signal \N__53680\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53675\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53657\ : std_logic;
signal \N__53652\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53646\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53644\ : std_logic;
signal \N__53641\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53625\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53613\ : std_logic;
signal \N__53610\ : std_logic;
signal \N__53607\ : std_logic;
signal \N__53594\ : std_logic;
signal \N__53591\ : std_logic;
signal \N__53590\ : std_logic;
signal \N__53587\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53579\ : std_logic;
signal \N__53576\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53559\ : std_logic;
signal \N__53552\ : std_logic;
signal \N__53543\ : std_logic;
signal \N__53540\ : std_logic;
signal \N__53535\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53516\ : std_logic;
signal \N__53513\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53505\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53495\ : std_logic;
signal \N__53486\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53480\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53447\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53422\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53396\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53377\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53327\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53317\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53305\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53257\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53251\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53242\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53240\ : std_logic;
signal \N__53239\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53236\ : std_logic;
signal \N__53233\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53231\ : std_logic;
signal \N__53230\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53224\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53216\ : std_logic;
signal \N__53215\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53213\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53208\ : std_logic;
signal \N__53207\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53197\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53193\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53183\ : std_logic;
signal \N__53182\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53169\ : std_logic;
signal \N__53168\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53166\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53164\ : std_logic;
signal \N__53163\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53159\ : std_logic;
signal \N__53158\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53153\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53146\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53143\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53139\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53135\ : std_logic;
signal \N__53134\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53123\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53120\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53111\ : std_logic;
signal \N__53108\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53102\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53098\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53091\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53081\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53074\ : std_logic;
signal \N__53069\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53018\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52985\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52972\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52967\ : std_logic;
signal \N__52964\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52945\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52941\ : std_logic;
signal \N__52940\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52938\ : std_logic;
signal \N__52937\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52915\ : std_logic;
signal \N__52912\ : std_logic;
signal \N__52909\ : std_logic;
signal \N__52906\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52884\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52873\ : std_logic;
signal \N__52870\ : std_logic;
signal \N__52867\ : std_logic;
signal \N__52864\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52855\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52841\ : std_logic;
signal \N__52838\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52819\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52808\ : std_logic;
signal \N__52803\ : std_logic;
signal \N__52800\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52766\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52741\ : std_logic;
signal \N__52738\ : std_logic;
signal \N__52735\ : std_logic;
signal \N__52732\ : std_logic;
signal \N__52729\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52720\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52718\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52657\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52633\ : std_logic;
signal \N__52630\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52617\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52581\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52550\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52537\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52517\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52466\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52382\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52360\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52354\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52325\ : std_logic;
signal \N__52324\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52321\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52317\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52310\ : std_logic;
signal \N__52309\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52299\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52256\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52250\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52152\ : std_logic;
signal \N__52151\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52139\ : std_logic;
signal \N__52136\ : std_logic;
signal \N__52131\ : std_logic;
signal \N__52128\ : std_logic;
signal \N__52123\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52103\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52079\ : std_logic;
signal \N__52070\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51988\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51941\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51936\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51902\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51839\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51832\ : std_logic;
signal \N__51831\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51828\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51822\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51807\ : std_logic;
signal \N__51806\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51796\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51736\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51713\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51575\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51534\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51527\ : std_logic;
signal \N__51524\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51509\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51485\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51423\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51337\ : std_logic;
signal \N__51334\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51305\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51302\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51202\ : std_logic;
signal \N__51199\ : std_logic;
signal \N__51196\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51088\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51058\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51034\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51028\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50992\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50965\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50958\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50942\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50926\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50894\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50728\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50683\ : std_logic;
signal \N__50680\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50503\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50115\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48915\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45325\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19051\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \ALU.N_675_0_0_cascade_\ : std_logic;
signal \ALU.N_703_0_0_0_cascade_\ : std_logic;
signal \ALU.N_681_0_0_0\ : std_logic;
signal \ALU.g0_0_2_cascade_\ : std_logic;
signal \ALU.N_699_0\ : std_logic;
signal \ALU.madd_167_cascade_\ : std_logic;
signal \ALU.madd_167\ : std_logic;
signal \ALU.g0_2\ : std_logic;
signal \ALU.a5_b_4_cascade_\ : std_logic;
signal \ALU.madd_139\ : std_logic;
signal \ALU.a2_b_8_cascade_\ : std_logic;
signal \ALU.madd_181_cascade_\ : std_logic;
signal \ALU.a3_b_8\ : std_logic;
signal \ALU.a3_b_8_cascade_\ : std_logic;
signal \ALU.madd_181\ : std_logic;
signal \ALU.madd_234_cascade_\ : std_logic;
signal \ALU.a7_b_8_cascade_\ : std_logic;
signal \ALU.madd_490_3\ : std_logic;
signal \ALU.madd_171_0_tz_cascade_\ : std_logic;
signal \ALU.madd_97\ : std_logic;
signal \ALU.madd_171_x_cascade_\ : std_logic;
signal \ALU.madd_171_0_tz\ : std_logic;
signal \ALU.madd_171_cascade_\ : std_logic;
signal \ALU.madd_315_0_tz_cascade_\ : std_logic;
signal \ALU.madd_214\ : std_logic;
signal \ALU.madd_311_cascade_\ : std_logic;
signal \ALU.madd_268\ : std_logic;
signal \ALU.madd_268_cascade_\ : std_logic;
signal \ALU.madd_311\ : std_logic;
signal \ALU.madd_316\ : std_logic;
signal \ALU.a8_b_5\ : std_logic;
signal \ALU.a1_b_13_cascade_\ : std_logic;
signal \ALU.madd_388_cascade_\ : std_logic;
signal \ALU.madd_403_cascade_\ : std_logic;
signal \ALU.a1_b_13\ : std_logic;
signal \ALU.madd_403_0_cascade_\ : std_logic;
signal \ALU.a_6_ns_1_2_cascade_\ : std_logic;
signal \TXbuffer_18_13_ns_1_2_cascade_\ : std_logic;
signal \TXbuffer_18_6_ns_1_2_cascade_\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_2_cascade_\ : std_logic;
signal \ALU.madd_417\ : std_logic;
signal \ALU.madd_490_1_0_cascade_\ : std_logic;
signal \ALU.madd_378_0\ : std_logic;
signal \ALU.madd_388\ : std_logic;
signal \ALU.madd_402_cascade_\ : std_logic;
signal \ALU.madd_330\ : std_logic;
signal \ALU.madd_490_21\ : std_logic;
signal \ALU.madd_397\ : std_logic;
signal \ALU.a6_b_9_cascade_\ : std_logic;
signal \ALU.madd_490_10_cascade_\ : std_logic;
signal \ALU.madd_490_7_cascade_\ : std_logic;
signal \ALU.madd_490_11\ : std_logic;
signal \ALU.a2_b_13\ : std_logic;
signal \TXbuffer_18_13_ns_1_0_cascade_\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_4_cascade_\ : std_logic;
signal \TXbuffer_18_15_ns_1_4_cascade_\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_0\ : std_logic;
signal \TXbuffer_18_15_ns_1_0_cascade_\ : std_logic;
signal \TXbuffer_18_10_ns_1_3_cascade_\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \TXbuffer_18_10_ns_1_4_cascade_\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_4\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_3\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal clkdiv_cry_0 : std_logic;
signal clkdiv_cry_1 : std_logic;
signal clkdiv_cry_2 : std_logic;
signal clkdiv_cry_3 : std_logic;
signal clkdiv_cry_4 : std_logic;
signal clkdiv_cry_5 : std_logic;
signal clkdiv_cry_6 : std_logic;
signal clkdiv_cry_7 : std_logic;
signal \clkdivZ0Z_8\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \clkdivZ0Z_9\ : std_logic;
signal clkdiv_cry_8 : std_logic;
signal \clkdivZ0Z_10\ : std_logic;
signal clkdiv_cry_9 : std_logic;
signal \clkdivZ0Z_11\ : std_logic;
signal clkdiv_cry_10 : std_logic;
signal \clkdivZ0Z_12\ : std_logic;
signal clkdiv_cry_11 : std_logic;
signal \clkdivZ0Z_13\ : std_logic;
signal clkdiv_cry_12 : std_logic;
signal \clkdivZ0Z_14\ : std_logic;
signal clkdiv_cry_13 : std_logic;
signal \clkdivZ0Z_15\ : std_logic;
signal clkdiv_cry_14 : std_logic;
signal clkdiv_cry_15 : std_logic;
signal \clkdivZ0Z_16\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \clkdivZ0Z_17\ : std_logic;
signal clkdiv_cry_16 : std_logic;
signal \clkdivZ0Z_18\ : std_logic;
signal clkdiv_cry_17 : std_logic;
signal \clkdivZ0Z_19\ : std_logic;
signal clkdiv_cry_18 : std_logic;
signal \clkdivZ0Z_20\ : std_logic;
signal clkdiv_cry_19 : std_logic;
signal \clkdivZ0Z_21\ : std_logic;
signal clkdiv_cry_20 : std_logic;
signal \clkdivZ0Z_22\ : std_logic;
signal clkdiv_cry_21 : std_logic;
signal clkdiv_cry_22 : std_logic;
signal \GPIO3_c\ : std_logic;
signal \ALU.madd_154_cascade_\ : std_logic;
signal \ALU.N_703_1_cascade_\ : std_logic;
signal \ALU.g0_cascade_\ : std_logic;
signal \ALU.madd_206\ : std_logic;
signal \ALU.madd_334_cascade_\ : std_logic;
signal \ALU.N_724_0_0_0\ : std_logic;
signal \ALU.madd_192_0\ : std_logic;
signal \ALU.madd_144\ : std_logic;
signal \ALU.g0_1\ : std_logic;
signal \ALU.N_695_0\ : std_logic;
signal \ALU.g0_4\ : std_logic;
signal \ALU.madd_197\ : std_logic;
signal \ALU.madd_112\ : std_logic;
signal \ALU.madd_191\ : std_logic;
signal \ALU.madd_234\ : std_logic;
signal \ALU.madd_112_cascade_\ : std_logic;
signal \ALU.madd_196_0\ : std_logic;
signal \ALU.madd_187\ : std_logic;
signal \ALU.madd_154\ : std_logic;
signal \ALU.madd_134\ : std_logic;
signal \ALU.g2_0_1\ : std_logic;
signal \ALU.madd_182_0\ : std_logic;
signal \ALU.a3_b_7\ : std_logic;
signal \ALU.a2_b_8\ : std_logic;
signal \ALU.madd_177\ : std_logic;
signal \ALU.madd_229\ : std_logic;
signal \ALU.madd_243_cascade_\ : std_logic;
signal \ALU.madd_219_0\ : std_logic;
signal \ALU.madd_181_0\ : std_logic;
signal \ALU.madd_315_0\ : std_logic;
signal \ALU.madd_320\ : std_logic;
signal \ALU.madd_393_cascade_\ : std_logic;
signal \ALU.madd_412\ : std_logic;
signal \ALU.madd_308_0_tz_0\ : std_logic;
signal \ALU.madd_299\ : std_logic;
signal \ALU.madd_209\ : std_logic;
signal \ALU.madd_243\ : std_logic;
signal \ALU.a0_b_13_cascade_\ : std_logic;
signal \ALU.madd_356\ : std_logic;
signal \ALU.madd_303_0\ : std_logic;
signal \ALU.madd_356_cascade_\ : std_logic;
signal \ALU.madd_175\ : std_logic;
signal \ALU.madd_388_0\ : std_logic;
signal \ALU.madd_393\ : std_logic;
signal \ALU.madd_340\ : std_logic;
signal \ALU.madd_355_cascade_\ : std_logic;
signal \ALU.madd_418\ : std_logic;
signal \ALU.madd_413_0\ : std_logic;
signal \ALU.madd_418_cascade_\ : std_logic;
signal \ALU.madd_293\ : std_logic;
signal \ALU.madd_336_0\ : std_logic;
signal \ALU.madd_351\ : std_logic;
signal \ALU.madd_346\ : std_logic;
signal \ALU.madd_172\ : std_logic;
signal \ALU.madd_346_cascade_\ : std_logic;
signal \ALU.madd_298_0\ : std_logic;
signal \ALU.madd_360\ : std_logic;
signal \ALU.madd_190\ : std_logic;
signal \ALU.madd_330_0_tz\ : std_logic;
signal \ALU.madd_326\ : std_logic;
signal \ALU.madd_326_cascade_\ : std_logic;
signal \ALU.madd_350_0\ : std_logic;
signal \ALU.madd_355\ : std_logic;
signal \ALU.madd_408\ : std_logic;
signal \ALU.madd_350_0_cascade_\ : std_logic;
signal \ALU.madd_422\ : std_logic;
signal \ALU.a7_b_7_cascade_\ : std_logic;
signal \ALU.madd_383\ : std_logic;
signal \ALU.b_9_cascade_\ : std_logic;
signal \ALU.madd_326_0\ : std_logic;
signal \ALU.a5_b_9_cascade_\ : std_logic;
signal \ALU.a6_b_8\ : std_logic;
signal \ALU.a5_b_9\ : std_logic;
signal \ALU.a6_b_8_cascade_\ : std_logic;
signal \ALU.madd_378\ : std_logic;
signal \ALU.b_i_3_cascade_\ : std_logic;
signal \ALU.a3_b_11\ : std_logic;
signal \ALU.madd_382\ : std_logic;
signal \ALU.a4_b_10\ : std_logic;
signal \ALU.a11_b_3_cascade_\ : std_logic;
signal \ALU.madd_373\ : std_logic;
signal \ALU.a11_b_3\ : std_logic;
signal \ALU.madd_392\ : std_logic;
signal \ALU.madd_490_16\ : std_logic;
signal \ALU.madd_490_15_cascade_\ : std_logic;
signal \ALU.madd_490_19\ : std_logic;
signal \ALU.madd_339\ : std_logic;
signal \ALU.madd_340_0\ : std_logic;
signal \ALU.madd_490_1\ : std_logic;
signal \ALU.madd_490_9\ : std_logic;
signal \ALU.madd_490_0_cascade_\ : std_logic;
signal \ALU.madd_490_13\ : std_logic;
signal \ALU.madd_490_14\ : std_logic;
signal \ALU.r2_RNIFR6TZ0Z_15_cascade_\ : std_logic;
signal \ALU.b_15_cascade_\ : std_logic;
signal \TXbuffer_18_13_ns_1_3\ : std_logic;
signal \ALU.r1_RNIAFSRZ0Z_15\ : std_logic;
signal \ALU.r5_RNIJBVTZ0Z_15_cascade_\ : std_logic;
signal \ALU.b_7_ns_1_15\ : std_logic;
signal \ALU.a_15_cascade_\ : std_logic;
signal \ALU.lshift_3_ns_1_15_cascade_\ : std_logic;
signal \ALU.b_6_ns_1_13_cascade_\ : std_logic;
signal \ALU.r6_RNIC9GA2Z0Z_13_cascade_\ : std_logic;
signal \ALU.b_13_cascade_\ : std_logic;
signal \TXbuffer_18_13_ns_1_4_cascade_\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_4\ : std_logic;
signal \ALU.N_661_0\ : std_logic;
signal \ALU.madd_155_cascade_\ : std_logic;
signal \ALU.madd_109_0_tz_cascade_\ : std_logic;
signal \ALU.madd_109_cascade_\ : std_logic;
signal \ALU.N_687_0\ : std_logic;
signal \ALU.madd_159_N_2L1\ : std_logic;
signal \ALU.madd_159\ : std_logic;
signal \ALU.madd_150\ : std_logic;
signal \ALU.madd_155\ : std_logic;
signal \ALU.a7_b_1_cascade_\ : std_logic;
signal \ALU.a6_b_2\ : std_logic;
signal \ALU.a6_b_2_cascade_\ : std_logic;
signal \ALU.a7_b_1\ : std_logic;
signal \ALU.madd_99_cascade_\ : std_logic;
signal \ALU.madd_149\ : std_logic;
signal \ALU.madd_99\ : std_logic;
signal \ALU.madd_145\ : std_logic;
signal \ALU.madd_244\ : std_logic;
signal \ALU.madd_201\ : std_logic;
signal \ALU.madd_239\ : std_logic;
signal \ALU.a3_b_9_cascade_\ : std_logic;
signal \ALU.a3_b_9\ : std_logic;
signal \ALU.a4_b_8\ : std_logic;
signal \ALU.a4_b_8_cascade_\ : std_logic;
signal \ALU.madd_269\ : std_logic;
signal \ALU.madd_274\ : std_logic;
signal \ALU.madd_269_cascade_\ : std_logic;
signal \ALU.madd_289\ : std_logic;
signal \ALU.madd_185_1_cascade_\ : std_logic;
signal \ALU.madd_106\ : std_logic;
signal \ALU.g0_2_N_2L1_cascade_\ : std_logic;
signal \ALU.madd_186_0\ : std_logic;
signal \ALU.madd_228\ : std_logic;
signal \ALU.madd_338\ : std_logic;
signal \ALU.madd_337\ : std_logic;
signal \ALU.a0_b_13\ : std_logic;
signal \ALU.madd_335_0\ : std_logic;
signal \ALU.madd_233\ : std_logic;
signal \ALU.madd_238\ : std_logic;
signal \ALU.madd_294\ : std_logic;
signal \ALU.madd_304\ : std_logic;
signal \ALU.madd_253\ : std_logic;
signal \ALU.madd_341\ : std_logic;
signal \ALU.madd_336\ : std_logic;
signal \ALU.madd_335\ : std_logic;
signal \ALU.madd_283\ : std_logic;
signal \ALU.madd_124_0\ : std_logic;
signal \ALU.madd_218_0_tz\ : std_logic;
signal \ALU.madd_218_cascade_\ : std_logic;
signal \ALU.madd_346_1\ : std_logic;
signal \ALU.a2_b_10\ : std_logic;
signal \ALU.a0_b_12_cascade_\ : std_logic;
signal \ALU.madd_279_0\ : std_logic;
signal \ALU.madd_331_0\ : std_logic;
signal \ALU.a0_b_12\ : std_logic;
signal \ALU.madd_218\ : std_logic;
signal \ALU.madd_202\ : std_logic;
signal \ALU.a12_b_0_cascade_\ : std_logic;
signal \ALU.madd_263\ : std_logic;
signal \ALU.madd_264_cascade_\ : std_logic;
signal \ALU.madd_288\ : std_logic;
signal \ALU.a12_b_0\ : std_logic;
signal \ALU.a10_b_2\ : std_logic;
signal \ALU.madd_259\ : std_logic;
signal \ALU.a7_b_5\ : std_logic;
signal \ALU.madd_259_cascade_\ : std_logic;
signal \ALU.madd_284_0\ : std_logic;
signal \ALU.b_3_ns_1_9_cascade_\ : std_logic;
signal \ALU.r4_RNIM58R1Z0Z_9\ : std_logic;
signal \ALU.b_3_ns_1_10_cascade_\ : std_logic;
signal \ALU.b_3_ns_1_11_cascade_\ : std_logic;
signal \ALU.r5_RNIQGFS1Z0Z_11_cascade_\ : std_logic;
signal \ALU.b_6_ns_1_10_cascade_\ : std_logic;
signal \ALU.b_6_ns_1_11_cascade_\ : std_logic;
signal \ALU.r6_RNI2H0U1Z0Z_11\ : std_logic;
signal \ALU.b_6_ns_1_9_cascade_\ : std_logic;
signal \ALU.r6_RNIUT042Z0Z_9\ : std_logic;
signal \ALU.r5_RNIH9VTZ0Z_14\ : std_logic;
signal \ALU.r1_RNI8DSRZ0Z_14_cascade_\ : std_logic;
signal \ALU.r2_RNIDP6TZ0Z_14\ : std_logic;
signal \ALU.b_7_ns_1_14_cascade_\ : std_logic;
signal \ALU.r6_RNILPNUZ0Z_14\ : std_logic;
signal \ALU.b_14_cascade_\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \ALU.r0_12_prm_8_11_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_11_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_11_s1\ : std_logic;
signal \ALU.r0_12_prm_7_11_s1\ : std_logic;
signal \ALU.r0_12_prm_5_11_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_11_s1\ : std_logic;
signal \ALU.r0_12_prm_5_11_s1\ : std_logic;
signal \ALU.r0_12_prm_4_11_s1\ : std_logic;
signal \ALU.r0_12_prm_3_11_s1\ : std_logic;
signal \ALU.r0_12_prm_2_11_s1\ : std_logic;
signal \ALU.r0_12_prm_1_11_s1_c_RNOZ0\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \ALU.r0_12_s1_11\ : std_logic;
signal \ALU.b_3_ns_1_12_cascade_\ : std_logic;
signal \ALU.b_6_ns_1_12_cascade_\ : std_logic;
signal \ALU.r6_RNI85GA2Z0Z_12\ : std_logic;
signal \ALU.r5_RNI05V82Z0Z_12\ : std_logic;
signal \ALU.r6_RNI85GA2Z0Z_12_cascade_\ : std_logic;
signal \ALU.b_3_ns_1_13_cascade_\ : std_logic;
signal \ALU.r5_RNI49V82Z0Z_13\ : std_logic;
signal \ALU.a_6_ns_1_15_cascade_\ : std_logic;
signal \ALU.r6_RNIH8772Z0Z_15\ : std_logic;
signal \ALU.r6_RNINRNUZ0Z_15\ : std_logic;
signal \TXbuffer_18_6_ns_1_0_cascade_\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_0\ : std_logic;
signal \TXbuffer_18_13_ns_1_7\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \ALU.r0_12_prm_8_11_s0_cy\ : std_logic;
signal \ALU.r5_RNIE0AK8_0Z0Z_11\ : std_logic;
signal \ALU.r0_12_prm_8_11_s0\ : std_logic;
signal \ALU.r0_12_prm_7_11_s0\ : std_logic;
signal \ALU.r5_RNIE0AK8_1Z0Z_11\ : std_logic;
signal \ALU.r0_12_prm_6_11_s0\ : std_logic;
signal \ALU.a_i_11\ : std_logic;
signal \ALU.r0_12_prm_5_11_s0\ : std_logic;
signal \ALU.r0_12_prm_3_11_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_11_s0\ : std_logic;
signal \ALU.r0_12_prm_3_11_s0\ : std_logic;
signal \ALU.r0_12_prm_2_11_s0\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \ALU.r0_12_s0_11\ : std_logic;
signal \ALU.r0_12_s0_11_THRU_CO\ : std_logic;
signal \ALU.g1_7_cascade_\ : std_logic;
signal \ALU.a4_b_0_0_5\ : std_logic;
signal \ALU.N_663_0_cascade_\ : std_logic;
signal \ALU.madd_109\ : std_logic;
signal \ALU.N_683_0_0_0\ : std_logic;
signal \ALU.madd_43_0_cascade_\ : std_logic;
signal \ALU.madd_77_0_tz\ : std_logic;
signal \ALU.madd_278\ : std_logic;
signal \ALU.madd_273\ : std_logic;
signal \ALU.madd_345\ : std_logic;
signal \ALU.madd_159_N_3L3\ : std_logic;
signal \ALU.madd_61\ : std_logic;
signal \ALU.madd_140_0\ : std_logic;
signal \ALU.madd_140_0_cascade_\ : std_logic;
signal \ALU.madd_155_1\ : std_logic;
signal \ALU.madd_144_0_tz\ : std_logic;
signal \ALU.a4_b_5\ : std_logic;
signal \ALU.g0_6_1\ : std_logic;
signal \ALU.r6_RNIUC0U1Z0Z_10\ : std_logic;
signal \ALU.r5_RNIMCFS1Z0Z_10\ : std_logic;
signal \ALU.a0_b_10\ : std_logic;
signal \ALU.a5_b_8_cascade_\ : std_logic;
signal \ALU.madd_325\ : std_logic;
signal \ALU.b_7_cascade_\ : std_logic;
signal \ALU.a5_b_7\ : std_logic;
signal \ALU.a5_b_5_cascade_\ : std_logic;
signal \ALU.madd_176\ : std_logic;
signal \ALU.a5_b_8\ : std_logic;
signal \ALU.a6_b_7\ : std_logic;
signal \ALU.madd_321\ : std_logic;
signal \ALU.b_6_ns_1_6_cascade_\ : std_logic;
signal \ALU.r6_RNIIH042Z0Z_6_cascade_\ : std_logic;
signal \ALU.b_6_cascade_\ : std_logic;
signal \ALU.g0_2_N_3L3\ : std_logic;
signal \bZ0Z_2\ : std_logic;
signal \ALU.b_3_ns_1_6_cascade_\ : std_logic;
signal \ALU.r4_RNIAP7R1Z0Z_6\ : std_logic;
signal \ALU.a0_b_14\ : std_logic;
signal \ALU.g2_0\ : std_logic;
signal \ALU.g0_2_N_4L5\ : std_logic;
signal \ALU.madd_134_0_tz\ : std_logic;
signal \ALU.madd_130_0\ : std_logic;
signal \ALU.madd_130\ : std_logic;
signal \ALU.madd_171_sx\ : std_logic;
signal \ALU.madd_213\ : std_logic;
signal \ALU.a9_b_3\ : std_logic;
signal \ALU.madd_167_0\ : std_logic;
signal \ALU.b_6_ns_1_5_cascade_\ : std_logic;
signal \ALU.b_3_ns_1_5_cascade_\ : std_logic;
signal \ALU.r6_RNIBP2O1Z0Z_5\ : std_logic;
signal \ALU.r4_RNI0QNE1Z0Z_5_cascade_\ : std_logic;
signal \ALU.b_5_cascade_\ : std_logic;
signal \TXbuffer_18_3_ns_1_1_cascade_\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_1_cascade_\ : std_logic;
signal r6_9 : std_logic;
signal \TXbuffer_18_6_ns_1_1_cascade_\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_1\ : std_logic;
signal r0_5 : std_logic;
signal \ALU.a_3_ns_1_5_cascade_\ : std_logic;
signal r2_10 : std_logic;
signal \ALU.a_6_ns_1_10_cascade_\ : std_logic;
signal \ALU.a_6_ns_1_11_cascade_\ : std_logic;
signal \ALU.r6_RNIT7372Z0Z_11_cascade_\ : std_logic;
signal \ALU.a_6_ns_1_7_cascade_\ : std_logic;
signal \ALU.b_6_ns_1_7_cascade_\ : std_logic;
signal \ALU.r6_RNIJ13O1Z0Z_7\ : std_logic;
signal r2_15 : std_logic;
signal r2_7 : std_logic;
signal \TXbuffer_18_6_ns_1_7_cascade_\ : std_logic;
signal r3_10 : std_logic;
signal r3_11 : std_logic;
signal r3_15 : std_logic;
signal r3_7 : std_logic;
signal \TXbuffer_18_13_ns_1_6_cascade_\ : std_logic;
signal \TXbuffer_18_3_ns_1_2_cascade_\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_2\ : std_logic;
signal \TXbuffer_18_3_ns_1_4\ : std_logic;
signal r6_10 : std_logic;
signal r6_15 : std_logic;
signal r7_10 : std_logic;
signal r7_11 : std_logic;
signal r7_15 : std_logic;
signal \TXbuffer_18_10_ns_1_6_cascade_\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_6\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \TXbuffer_18_6_ns_1_6\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_6_cascade_\ : std_logic;
signal \TXbuffer_18_15_ns_1_6\ : std_logic;
signal \TXbuffer_18_3_ns_1_6_cascade_\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_6\ : std_logic;
signal \ALU.r0_12_prm_4_11_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNIAFVE5Z0Z_11\ : std_logic;
signal \ALU.r0_12_prm_5_11_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_11_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_11_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_11_s1_c_RNOZ0\ : std_logic;
signal \TXbuffer_18_3_ns_1_5\ : std_logic;
signal \ALU.a4_b_4_cascade_\ : std_logic;
signal \ALU.madd_104\ : std_logic;
signal \ALU.madd_68_cascade_\ : std_logic;
signal \ALU.madd_82_0_cascade_\ : std_logic;
signal \ALU.madd_119\ : std_logic;
signal \ALU.a_6_cascade_\ : std_logic;
signal \ALU.g3\ : std_logic;
signal \ALU.madd_72_0_tz\ : std_logic;
signal \ALU.madd_40_cascade_\ : std_logic;
signal \ALU.madd_72\ : std_logic;
signal \ALU.madd_95\ : std_logic;
signal \ALU.madd_72_cascade_\ : std_logic;
signal \ALU.madd_77\ : std_logic;
signal \ALU.b_8_cascade_\ : std_logic;
signal \ALU.madd_82\ : std_logic;
signal \ALU.madd_127_cascade_\ : std_logic;
signal \ALU.madd_223\ : std_logic;
signal \ALU.madd_223_0_tz\ : std_logic;
signal \ALU.madd_105_0\ : std_logic;
signal \ALU.r4_RNIU5NK1Z0Z_8\ : std_logic;
signal \ALU.un9_addsub_axb_1_cascade_\ : std_logic;
signal \ALU.a7_b_3\ : std_logic;
signal \ALU.a_1_cascade_\ : std_logic;
signal \ALU.madd_228_0_tz\ : std_logic;
signal \ALU.a_9_cascade_\ : std_logic;
signal \ALU.N_675_1\ : std_logic;
signal \ALU.bZ0Z_0_cascade_\ : std_logic;
signal \ALU.madd_130_0_0\ : std_logic;
signal \ALU.r6_RNIGC3D2Z0Z_7\ : std_logic;
signal \ALU.a_7_cascade_\ : std_logic;
signal \ALU.madd_76\ : std_logic;
signal \ALU.madd_213_0_tz\ : std_logic;
signal \ALU.madd_209_0\ : std_logic;
signal \ALU.a8_b_4\ : std_logic;
signal \ALU.g0_7_x1_cascade_\ : std_logic;
signal \ALU.madd_76_1\ : std_logic;
signal \ALU.r6_RNIPK3D2Z0Z_9\ : std_logic;
signal \ALU.a9_b_4\ : std_logic;
signal \ALU.a_8_cascade_\ : std_logic;
signal \ALU.madd_224_0\ : std_logic;
signal \ALU.madd_224\ : std_logic;
signal \ALU.madd_121\ : std_logic;
signal \ALU.b_3_ns_1_8\ : std_logic;
signal r2_2 : std_logic;
signal r3_2 : std_logic;
signal \ALU.b_6_ns_1_2_cascade_\ : std_logic;
signal \ALU.b_6_ns_1_3_cascade_\ : std_logic;
signal r7_0 : std_logic;
signal \ALU.b_6_ns_1_0_cascade_\ : std_logic;
signal r6_0 : std_logic;
signal \ALU.a_3_ns_1_6_cascade_\ : std_logic;
signal r0_6 : std_logic;
signal \ALU.a_6_ns_1_5_cascade_\ : std_logic;
signal r3_6 : std_logic;
signal \ALU.a_6_ns_1_6_cascade_\ : std_logic;
signal \ALU.a_6_ns_1_9\ : std_logic;
signal \ALU.a_6_ns_1_8_cascade_\ : std_logic;
signal \ALU.r6_RNIKG3D2Z0Z_8\ : std_logic;
signal r2_8 : std_logic;
signal r3_8 : std_logic;
signal \ALU.b_6_ns_1_8_cascade_\ : std_logic;
signal \ALU.r6_RNIN53O1Z0Z_8\ : std_logic;
signal \ALU.a_6_ns_1_1_cascade_\ : std_logic;
signal \ALU.a_3_ns_1_10_cascade_\ : std_logic;
signal \ALU.r5_RNIVQN52Z0Z_10_cascade_\ : std_logic;
signal \ALU.a_3_ns_1_11_cascade_\ : std_logic;
signal \ALU.r5_RNI3VN52Z0Z_11\ : std_logic;
signal r3_3 : std_logic;
signal \ALU.a_6_ns_1_3_cascade_\ : std_logic;
signal \ALU.a_3_ns_1_12_cascade_\ : std_logic;
signal r7_12 : std_logic;
signal \ALU.a_6_ns_1_12_cascade_\ : std_logic;
signal \ALU.r6_RNI5S672Z0Z_12_cascade_\ : std_logic;
signal \ALU.r5_RNIS3672Z0Z_12\ : std_logic;
signal r2_5 : std_logic;
signal r2_6 : std_logic;
signal r2_9 : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \ALU.r0_12_prm_8_15_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_15_s1\ : std_logic;
signal \ALU.r0_12_prm_6_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_15_s1\ : std_logic;
signal \ALU.r0_12_prm_6_15_s1\ : std_logic;
signal \ALU.r0_12_prm_4_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_15_s1\ : std_logic;
signal \ALU.r0_12_prm_4_15_s1\ : std_logic;
signal \ALU.r0_12_prm_3_15_s1\ : std_logic;
signal \ALU.r0_12_prm_2_15_s1\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \ALU.madd_axb_14\ : std_logic;
signal \ALU.r0_12_s1_15\ : std_logic;
signal \ALU.a_3_ns_1_13_cascade_\ : std_logic;
signal r2_13 : std_logic;
signal \ALU.a_6_ns_1_13_cascade_\ : std_logic;
signal \ALU.r6_RNI90772Z0Z_13_cascade_\ : std_logic;
signal \ALU.r5_RNI10M52Z0Z_13\ : std_logic;
signal \ALU.r5_RNIPV8A9Z0Z_13_cascade_\ : std_logic;
signal r3_12 : std_logic;
signal r3_5 : std_logic;
signal r3_13 : std_logic;
signal r6_13 : std_logic;
signal \TXbuffer_18_6_ns_1_5\ : std_logic;
signal r6_5 : std_logic;
signal \TXbuffer_RNO_5Z0Z_5\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_5_cascade_\ : std_logic;
signal r7_13 : std_logic;
signal r7_5 : std_logic;
signal \TXbuffer_18_13_ns_1_5\ : std_logic;
signal \TXbuffer_18_10_ns_1_5\ : std_logic;
signal \ALU.madd_68_0\ : std_logic;
signal \ALU.madd_46_0\ : std_logic;
signal \ALU.madd_100\ : std_logic;
signal \ALU.madd_105\ : std_logic;
signal \ALU.madd_46_0_cascade_\ : std_logic;
signal \ALU.madd_82_0\ : std_logic;
signal \ALU.a5_b_3\ : std_logic;
signal \ALU.g2_0_0_0\ : std_logic;
signal \ALU.a0_b_7\ : std_logic;
signal \ALU.a5_b_0\ : std_logic;
signal \ALU.madd_38_cascade_\ : std_logic;
signal \ALU.madd_87_cascade_\ : std_logic;
signal \ALU.madd_92_cascade_\ : std_logic;
signal \ALU.madd_78_0\ : std_logic;
signal \ALU.madd_68\ : std_logic;
signal \ALU.madd_78_0_cascade_\ : std_logic;
signal \ALU.madd_60\ : std_logic;
signal \ALU.madd_332_cascade_\ : std_logic;
signal \ALU.r6_RNIA0841Z0Z_0\ : std_logic;
signal \ALU.madd_92\ : std_logic;
signal \ALU.madd_120\ : std_logic;
signal \ALU.r6_RNII9FT1Z0Z_3\ : std_logic;
signal \ALU.b_3_cascade_\ : std_logic;
signal \ALU.un2_addsub_axb_3\ : std_logic;
signal \ALU.b_1_cascade_\ : std_logic;
signal \ALU.a4_b_1\ : std_logic;
signal \ALU.a_3_cascade_\ : std_logic;
signal \ALU.g1_1\ : std_logic;
signal \ALU.b_4_cascade_\ : std_logic;
signal \ALU.madd_214_0\ : std_logic;
signal \ALU.b_2_cascade_\ : std_logic;
signal \ALU.madd_134_0_tz_0\ : std_logic;
signal \ALU.madd_172_0\ : std_logic;
signal \ALU.madd_368\ : std_logic;
signal \ALU.a12_b_2\ : std_logic;
signal \ALU.a12_b_2_cascade_\ : std_logic;
signal \ALU.madd_372\ : std_logic;
signal \ALU.g1_2\ : std_logic;
signal \ALU.madd_311_0\ : std_logic;
signal \b_1_repZ0Z1\ : std_logic;
signal \b_1_repZ0Z2\ : std_logic;
signal r0_11 : std_logic;
signal \TXbuffer_18_3_ns_1_3_cascade_\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_3_cascade_\ : std_logic;
signal \TXbuffer_18_15_ns_1_3\ : std_logic;
signal r2_11 : std_logic;
signal r2_3 : std_logic;
signal r6_11 : std_logic;
signal \TXbuffer_18_6_ns_1_3_cascade_\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_3\ : std_logic;
signal r4_11 : std_logic;
signal \bZ0Z_0\ : std_logic;
signal \a_0_repZ0Z1\ : std_logic;
signal \ALU.a_6_ns_1_4_cascade_\ : std_logic;
signal r3_4 : std_logic;
signal \b_0_repZ0Z1\ : std_logic;
signal \ALU.b_6_ns_1_4_cascade_\ : std_logic;
signal \ALU.r6_RNI7L2O1Z0Z_4\ : std_logic;
signal \ALU.r6_RNI7L2O1Z0Z_4_cascade_\ : std_logic;
signal r2_12 : std_logic;
signal r2_4 : std_logic;
signal \TXbuffer_18_6_ns_1_4_cascade_\ : std_logic;
signal r6_12 : std_logic;
signal \TXbuffer_RNO_6Z0Z_4\ : std_logic;
signal r1_11 : std_logic;
signal r1_12 : std_logic;
signal r1_13 : std_logic;
signal r4_10 : std_logic;
signal r4_12 : std_logic;
signal r4_13 : std_logic;
signal r4_5 : std_logic;
signal r4_6 : std_logic;
signal \ALU.a_3_ns_1_14_cascade_\ : std_logic;
signal r4_14 : std_logic;
signal r2_14 : std_logic;
signal r3_14 : std_logic;
signal r7_14 : std_logic;
signal \ALU.a_6_ns_1_14_cascade_\ : std_logic;
signal r6_14 : std_logic;
signal \ALU.r6_RNID4772Z0Z_14_cascade_\ : std_logic;
signal \ALU.r5_RNI54M52Z0Z_14\ : std_logic;
signal r0_14 : std_logic;
signal \aZ0Z_0\ : std_logic;
signal \aZ0Z_2\ : std_logic;
signal \ALU.a_3_ns_1_15_cascade_\ : std_logic;
signal \ALU.r5_RNI98M52Z0Z_15\ : std_logic;
signal \ALU.r0_12_11\ : std_logic;
signal r5_11 : std_logic;
signal r5_12 : std_logic;
signal r5_13 : std_logic;
signal r5_14 : std_logic;
signal \ALU.r0_12_15\ : std_logic;
signal r5_5 : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \ALU.r0_12_prm_8_13_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_8_13_s0\ : std_logic;
signal \ALU.r0_12_prm_7_13_s0\ : std_logic;
signal \ALU.r0_12_prm_6_13_s0\ : std_logic;
signal \ALU.r0_12_prm_5_13_s0\ : std_logic;
signal \ALU.r0_12_prm_3_13_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_13_s0\ : std_logic;
signal \ALU.r0_12_prm_3_13_s0\ : std_logic;
signal \ALU.r0_12_prm_2_13_s0\ : std_logic;
signal \bfn_6_16_0_\ : std_logic;
signal \ALU.r0_12_s0_13\ : std_logic;
signal \ALU.r0_12_13\ : std_logic;
signal r0_13 : std_logic;
signal \ALU.r5_RNIK81F5Z0Z_13\ : std_logic;
signal \ALU.r0_12_prm_5_13_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_13_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_13_s0_c_RNOZ0\ : std_logic;
signal \ALU.madd_334\ : std_logic;
signal \ALU.madd_333\ : std_logic;
signal \ALU.madd_87\ : std_logic;
signal \ALU.madd_110\ : std_logic;
signal \ALU.madd_115\ : std_logic;
signal \ALU.madd_124\ : std_logic;
signal \ALU.madd_124_cascade_\ : std_logic;
signal \ALU.madd_160\ : std_logic;
signal \ALU.r6_RNIE0JB2Z0Z_6\ : std_logic;
signal \ALU.r4_RNI68Q22Z0Z_6\ : std_logic;
signal \ALU.a3_b_1\ : std_logic;
signal \ALU.a3_b_1_cascade_\ : std_logic;
signal \ALU.madd_18_cascade_\ : std_logic;
signal \ALU.madd_43_cascade_\ : std_logic;
signal \ALU.a2_b_3\ : std_logic;
signal \ALU.madd_332\ : std_logic;
signal \ALU.madd_94\ : std_logic;
signal \ALU.madd_33\ : std_logic;
signal \ALU.madd_38\ : std_logic;
signal \ALU.a0_b_6\ : std_logic;
signal \ALU.madd_51\ : std_logic;
signal \ALU.madd_51_cascade_\ : std_logic;
signal \ALU.madd_43\ : std_logic;
signal \ALU.madd_331\ : std_logic;
signal \ALU.a1_b_4\ : std_logic;
signal \ALU.madd_73_0_cascade_\ : std_logic;
signal \ALU.a1_b_5\ : std_logic;
signal \ALU.a2_b_4\ : std_logic;
signal \ALU.a1_b_5_cascade_\ : std_logic;
signal \b_fastZ0Z_1\ : std_logic;
signal \b_2_repZ0Z2\ : std_logic;
signal \ALU.r4_RNIMTDQZ0Z_1_cascade_\ : std_logic;
signal \ALU.b_7_ns_1_1\ : std_logic;
signal \ALU.madd_46\ : std_logic;
signal \ALU.a5_b_1\ : std_logic;
signal \ALU.a5_b_1_cascade_\ : std_logic;
signal \ALU.madd_50\ : std_logic;
signal \ALU.madd_55\ : std_logic;
signal \ALU.madd_50_cascade_\ : std_logic;
signal \ALU.madd_73\ : std_logic;
signal \ALU.madd_83\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_2\ : std_logic;
signal \TXbuffer_18_15_ns_1_2\ : std_logic;
signal \clkdivZ0Z_1\ : std_logic;
signal \clkdivZ0Z_2\ : std_logic;
signal \clkdivZ0Z_3\ : std_logic;
signal \clkdivZ0Z_0\ : std_logic;
signal params5 : std_logic;
signal \ALU.madd_axb_3_cascade_\ : std_logic;
signal \ALU.madd_14\ : std_logic;
signal \ALU.madd_cry_0_ma\ : std_logic;
signal \ALU.madd_axb_0_l_ofx\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \ALU.madd_cry_0\ : std_logic;
signal \ALU.madd_cry_1\ : std_logic;
signal \ALU.madd_cry_2\ : std_logic;
signal \ALU.madd_cry_3\ : std_logic;
signal \ALU.madd_axb_5_l_fx\ : std_logic;
signal \ALU.madd_cry_4\ : std_logic;
signal \ALU.madd_axb_6_l_ofx\ : std_logic;
signal \ALU.madd_cry_5\ : std_logic;
signal \ALU.madd_cry_6\ : std_logic;
signal \ALU.madd_cry_7\ : std_logic;
signal \ALU.madd_165\ : std_logic;
signal \ALU.madd_axb_8_l_fx\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \ALU.madd_axb_9_l_ofx\ : std_logic;
signal \ALU.madd_cry_9_ma\ : std_logic;
signal \ALU.madd_cry_8\ : std_logic;
signal \ALU.madd_axb_10\ : std_logic;
signal \ALU.madd_cry_9_THRU_CO\ : std_logic;
signal \ALU.madd_cry_9\ : std_logic;
signal \ALU.g0_13\ : std_logic;
signal \ALU.madd_axb_11_l_fx\ : std_logic;
signal \ALU.madd_cry_10\ : std_logic;
signal \ALU.madd_cry_12_ma\ : std_logic;
signal \ALU.madd_axb_12_l_ofx\ : std_logic;
signal \ALU.mult_13\ : std_logic;
signal \ALU.madd_cry_11\ : std_logic;
signal \ALU.madd_axb_13_l_ofx\ : std_logic;
signal \ALU.madd_cry_13_ma\ : std_logic;
signal \ALU.madd_cry_12\ : std_logic;
signal \ALU.madd_cry_13\ : std_logic;
signal \ALU.madd_cry_13_THRU_CO\ : std_logic;
signal \ALU.a13_b_1\ : std_logic;
signal \ALU.madd_373_0\ : std_logic;
signal \ALU.madd_368_0\ : std_logic;
signal \ALU.a9_b_5\ : std_logic;
signal \ALU.madd_398_0\ : std_logic;
signal \ALU.r4_RNIJJH11Z0Z_0\ : std_logic;
signal \ALU.r0_RNIBROOZ0Z_0_cascade_\ : std_logic;
signal \a_fastZ0Z_1\ : std_logic;
signal \ALU.a_7_ns_1_0\ : std_logic;
signal r4_0 : std_logic;
signal \TXbuffer_18_3_ns_1_0_cascade_\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_0\ : std_logic;
signal \TXbuffer_18_10_ns_1_0_cascade_\ : std_logic;
signal r5_0 : std_logic;
signal \TXbuffer_RNO_0Z0Z_0\ : std_logic;
signal r3_9 : std_logic;
signal \TXbuffer_18_13_ns_1_1\ : std_logic;
signal \TXbuffer_18_10_ns_1_1_cascade_\ : std_logic;
signal \TXbuffer_18_15_ns_1_1\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_1\ : std_logic;
signal r1_10 : std_logic;
signal r5_10 : std_logic;
signal \TXbuffer_18_10_ns_1_2_cascade_\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_2\ : std_logic;
signal r7_6 : std_logic;
signal r7_7 : std_logic;
signal r7_8 : std_logic;
signal r7_9 : std_logic;
signal r7_2 : std_logic;
signal r7_3 : std_logic;
signal r7_4 : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \ALU.r0_12_prm_8_10_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_8_10_s0\ : std_logic;
signal \ALU.r0_12_prm_7_10_s0\ : std_logic;
signal \ALU.r0_12_prm_6_10_s0\ : std_logic;
signal \ALU.r0_12_prm_5_10_s0\ : std_logic;
signal \ALU.r0_12_prm_3_10_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_10_s0\ : std_logic;
signal \ALU.r0_12_prm_3_10_s0\ : std_logic;
signal \ALU.r0_12_prm_2_10_s0\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \ALU.mult_10\ : std_logic;
signal \ALU.r0_12_s0_10\ : std_logic;
signal \ALU.r0_12_10\ : std_logic;
signal r0_10 : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \ALU.r0_12_prm_8_14_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_8_14_s0\ : std_logic;
signal \ALU.r0_12_prm_7_14_s0\ : std_logic;
signal \ALU.r0_12_prm_6_14_s0\ : std_logic;
signal \ALU.r0_12_prm_5_14_s0\ : std_logic;
signal \ALU.r0_12_prm_3_14_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_14_s0\ : std_logic;
signal \ALU.r0_12_prm_3_14_s0\ : std_logic;
signal \ALU.r0_12_prm_2_14_s0\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \ALU.mult_14\ : std_logic;
signal \ALU.r0_12_s0_14\ : std_logic;
signal \ALU.r0_12_14\ : std_logic;
signal r1_14 : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \ALU.r0_12_prm_8_12_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_8_12_s0\ : std_logic;
signal \ALU.r0_12_prm_7_12_s0\ : std_logic;
signal \ALU.r0_12_prm_6_12_s0\ : std_logic;
signal \ALU.r0_12_prm_5_12_s0\ : std_logic;
signal \ALU.r0_12_prm_3_12_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_12_s0\ : std_logic;
signal \ALU.r0_12_prm_3_12_s0\ : std_logic;
signal \ALU.r0_12_prm_2_12_s0\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \ALU.mult_12\ : std_logic;
signal \ALU.r0_12_s0_12\ : std_logic;
signal \ALU.r0_12_12\ : std_logic;
signal r0_12 : std_logic;
signal \TXbuffer_RNO_1Z0Z_5\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_5\ : std_logic;
signal \TXbuffer_18_15_ns_1_5\ : std_logic;
signal \ALU.a2_b_1_cascade_\ : std_logic;
signal \ALU.a1_b_2\ : std_logic;
signal \ALU.a2_b_1\ : std_logic;
signal \ALU.a1_b_2_cascade_\ : std_logic;
signal \ALU.madd_29_0\ : std_logic;
signal \ALU.madd_18\ : std_logic;
signal \ALU.madd_34\ : std_logic;
signal \ALU.madd_39_cascade_\ : std_logic;
signal \ALU.madd_39\ : std_logic;
signal \ALU.madd_23_cascade_\ : std_logic;
signal \ALU.madd_28\ : std_logic;
signal \ALU.madd_axb_4_l_fx\ : std_logic;
signal \ALU.madd_8\ : std_logic;
signal \ALU.madd_19\ : std_logic;
signal \ALU.madd_66\ : std_logic;
signal \a_1_repZ0Z1\ : std_logic;
signal \ALU.r6_RNIASIB2Z0Z_5\ : std_logic;
signal \ALU.r4_RNI24Q22Z0Z_5\ : std_logic;
signal \ALU.a0_b_4\ : std_logic;
signal \ALU.un2_addsub_axb_2\ : std_logic;
signal \ALU.madd_56\ : std_logic;
signal \ALU.madd_45\ : std_logic;
signal \ALU.madd_cry_6_ma\ : std_logic;
signal r3_0 : std_logic;
signal \a_0_repZ0Z2\ : std_logic;
signal \ALU.r2_RNI18BOZ0Z_0\ : std_logic;
signal r2_0 : std_logic;
signal r3_1 : std_logic;
signal r2_1 : std_logic;
signal \ALU.r2_RNI4H0SZ0Z_1\ : std_logic;
signal \b_0_repZ0Z2\ : std_logic;
signal r7_1 : std_logic;
signal r6_1 : std_logic;
signal \ALU.r6_RNIC9P41Z0Z_1\ : std_logic;
signal \ALU.r6_RNIE5FT1Z0Z_2\ : std_logic;
signal \ALU.madd_13\ : std_logic;
signal \ALU.a2_b_0\ : std_logic;
signal \ALU.madd_3\ : std_logic;
signal \ALU.madd_4\ : std_logic;
signal \ALU.madd_3_cascade_\ : std_logic;
signal \ALU.a0_b_3\ : std_logic;
signal \ALU.a3_b_2\ : std_logic;
signal \ALU.rshift_3_ns_1_7_cascade_\ : std_logic;
signal \ALU.b_3_ns_1_7_cascade_\ : std_logic;
signal \ALU.r4_RNI82OE1Z0Z_7\ : std_logic;
signal r1_15 : std_logic;
signal r5_15 : std_logic;
signal \TXbuffer_18_10_ns_1_7_cascade_\ : std_logic;
signal \clkdivZ0Z_7\ : std_logic;
signal r0_15 : std_logic;
signal \clkdivZ0Z_6\ : std_logic;
signal \TXbuffer_18_3_ns_1_7_cascade_\ : std_logic;
signal r4_15 : std_logic;
signal \clkdivZ0Z_5\ : std_logic;
signal \TXbuffer_RNO_5Z0Z_7_cascade_\ : std_logic;
signal \TXbuffer_RNO_6Z0Z_7\ : std_logic;
signal \ALU.a_3_ns_1_1_cascade_\ : std_logic;
signal r0_7 : std_logic;
signal \ALU.a_3_ns_1_7_cascade_\ : std_logic;
signal \ALU.r4_RNI6BA92Z0Z_7\ : std_logic;
signal r1_8 : std_logic;
signal \ALU.a_3_ns_1_8_cascade_\ : std_logic;
signal \ALU.r4_RNIAFA92Z0Z_8\ : std_logic;
signal \ALU.a_3_ns_1_3\ : std_logic;
signal \ALU.a_3_ns_1_2_cascade_\ : std_logic;
signal \a_2_repZ0Z1\ : std_logic;
signal \ALU.a_3_ns_1_4_cascade_\ : std_logic;
signal \a_fastZ0Z_2\ : std_logic;
signal r1_9 : std_logic;
signal \a_fastZ0Z_0\ : std_logic;
signal \a_2_repZ0Z2\ : std_logic;
signal \ALU.a_3_ns_1_9_cascade_\ : std_logic;
signal \ALU.r4_RNIEJA92Z0Z_9\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \ALU.r0_12_prm_8_9_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_8_9_s0\ : std_logic;
signal \ALU.r0_12_prm_6_9_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_9_s0\ : std_logic;
signal \ALU.r0_12_prm_6_9_s0\ : std_logic;
signal \ALU.r0_12_prm_5_9_s0\ : std_logic;
signal \ALU.r0_12_prm_3_9_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_9_s0\ : std_logic;
signal \ALU.r0_12_prm_2_9_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_9_s0\ : std_logic;
signal \ALU.r0_12_prm_2_9_s0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \ALU.mult_9\ : std_logic;
signal \ALU.r0_12_s0_9\ : std_logic;
signal r0_9 : std_logic;
signal \ALU.r0_12_prm_8_11_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_12_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_2_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_2_13_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_1_14_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.rshift_10_ns_1_3\ : std_logic;
signal \ALU.r5_RNI465TIZ0Z_13_cascade_\ : std_logic;
signal \ALU.r5_RNIOL1S71Z0Z_10\ : std_logic;
signal \ALU.r0_12_prm_5_12_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_11_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_12_s0_c_RNOZ0\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \ALU.r0_12_prm_8_13_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNID2JJ9_0Z0Z_13\ : std_logic;
signal \ALU.r0_12_prm_8_13_s1\ : std_logic;
signal \ALU.r0_12_prm_6_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_13\ : std_logic;
signal \ALU.r0_12_prm_7_13_s1\ : std_logic;
signal \ALU.r0_12_prm_5_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNID2JJ9_1Z0Z_13\ : std_logic;
signal \ALU.r0_12_prm_6_13_s1\ : std_logic;
signal \ALU.r0_12_prm_4_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_13\ : std_logic;
signal \ALU.r0_12_prm_5_13_s1\ : std_logic;
signal \ALU.r0_12_prm_4_13_s1\ : std_logic;
signal \ALU.r0_12_prm_3_13_s1\ : std_logic;
signal \ALU.r0_12_prm_2_13_s1\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \ALU.r0_12_s1_13\ : std_logic;
signal \ALU.r0_12_s1_13_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_1_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.rshift_3_ns_1_2_cascade_\ : std_logic;
signal \ALU.r6_RNIFJ8D2Z0Z_3\ : std_logic;
signal \ALU.r4_RNIMQ992Z0Z_3\ : std_logic;
signal \ALU.r4_RNIDI992Z0Z_1\ : std_logic;
signal \ALU.r6_RNI7B8D2Z0Z_1\ : std_logic;
signal \ALU.a1_b_3\ : std_logic;
signal \ALU.madd_135_0\ : std_logic;
signal \ALU.lshift_3_ns_1_6\ : std_logic;
signal \ALU.lshift_3_ns_1_7\ : std_logic;
signal \ALU.un9_addsub_axb_3\ : std_logic;
signal \ALU.madd_490_5\ : std_logic;
signal \ALU.rshift_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_3_c_RNOZ0Z_3_cascade_\ : std_logic;
signal \ALU.r5_RNI67NNKZ0Z_10\ : std_logic;
signal \bZ0Z_1\ : std_logic;
signal \ALU.r6_RNI6TET1Z0Z_0\ : std_logic;
signal \ALU.r4_RNIC5NE1Z0Z_0\ : std_logic;
signal \ALU.r6_RNIBF8D2Z0Z_2\ : std_logic;
signal \ALU.r4_RNIHM992Z0Z_2\ : std_logic;
signal \ALU.r6_RNI403D2Z0Z_4\ : std_logic;
signal \ALU.r4_RNIQU992Z0Z_4\ : std_logic;
signal \aZ0Z_1\ : std_logic;
signal \ALU.un2_addsub_axb_4_cascade_\ : std_logic;
signal \ALU.rshift_10\ : std_logic;
signal \ALU.madd_76_0\ : std_logic;
signal \ALU.lshift_3_ns_1_11_cascade_\ : std_logic;
signal \ALU.un9_addsub_axb_4\ : std_logic;
signal \ALU.lshift_3_ns_1_9\ : std_logic;
signal r1_1 : std_logic;
signal \ALU.r0_RNIE5LHZ0Z_1\ : std_logic;
signal \ALU.b_3_ns_1_0\ : std_logic;
signal r0_4 : std_logic;
signal r1_4 : std_logic;
signal \ALU.b_3_ns_1_4_cascade_\ : std_logic;
signal \ALU.r4_RNISLNE1Z0Z_4\ : std_logic;
signal r0_2 : std_logic;
signal r1_2 : std_logic;
signal \ALU.b_3_ns_1_2_cascade_\ : std_logic;
signal \ALU.r4_RNIKDNE1Z0Z_2\ : std_logic;
signal \b_fastZ0Z_2\ : std_logic;
signal r1_3 : std_logic;
signal \b_fastZ0Z_0\ : std_logic;
signal \b_2_repZ0Z1\ : std_logic;
signal r4_3 : std_logic;
signal \ALU.b_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.r4_RNIOHNE1Z0Z_3\ : std_logic;
signal r5_6 : std_logic;
signal r5_7 : std_logic;
signal r5_8 : std_logic;
signal r5_9 : std_logic;
signal r5_1 : std_logic;
signal r5_2 : std_logic;
signal r5_3 : std_logic;
signal r5_4 : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \ALU.r4_RNIUES39Z0Z_1\ : std_logic;
signal \ALU.un2_addsub_cry_0\ : std_logic;
signal \ALU.r4_RNIUM9JCZ0Z_2\ : std_logic;
signal \ALU.b_i_2\ : std_logic;
signal \ALU.un2_addsub_cry_1\ : std_logic;
signal \ALU.r4_RNINFAJCZ0Z_3\ : std_logic;
signal \ALU.b_i_3\ : std_logic;
signal \ALU.un2_addsub_cry_2\ : std_logic;
signal \ALU.r4_RNI20C8CZ0Z_4\ : std_logic;
signal \ALU.b_i_4\ : std_logic;
signal \ALU.un2_addsub_cry_3\ : std_logic;
signal \ALU.r4_RNI8B628_1Z0Z_5\ : std_logic;
signal \ALU.un2_addsub_cry_4\ : std_logic;
signal \ALU.r4_RNI2BKQ8_1Z0Z_6\ : std_logic;
signal \ALU.un2_addsub_cry_5\ : std_logic;
signal \ALU.un2_addsub_cry_6\ : std_logic;
signal \ALU.un2_addsub_cry_7\ : std_logic;
signal \ALU.r4_RNIKUMQ8_1Z0Z_8\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \ALU.un2_addsub_cry_8\ : std_logic;
signal \ALU.r5_RNIUF9K8_2Z0Z_10\ : std_logic;
signal \ALU.un2_addsub_cry_9\ : std_logic;
signal \ALU.r5_RNIE0AK8_2Z0Z_11\ : std_logic;
signal \ALU.un2_addsub_cry_10\ : std_logic;
signal \ALU.r5_RNISP2L9_2Z0Z_12\ : std_logic;
signal \ALU.un2_addsub_cry_11\ : std_logic;
signal \ALU.r5_RNID2JJ9_2Z0Z_13\ : std_logic;
signal \ALU.un2_addsub_cry_12\ : std_logic;
signal \ALU.r2_RNINPPC9_2Z0Z_14\ : std_logic;
signal \ALU.un2_addsub_cry_13\ : std_logic;
signal \ALU.un2_addsub_cry_14\ : std_logic;
signal r4_7 : std_logic;
signal r4_8 : std_logic;
signal \ALU.r0_12_9\ : std_logic;
signal r4_9 : std_logic;
signal r4_1 : std_logic;
signal r4_2 : std_logic;
signal r4_4 : std_logic;
signal \ALU.r5_RNIVF7TIZ0Z_13\ : std_logic;
signal \ALU.lshift_15_ns_1_15_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_11_s1_c_RNOZ0Z_1\ : std_logic;
signal \ALU.r0_12_prm_2_11_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_1_10_s0_c_RNOZ0\ : std_logic;
signal \ALU.N_884_i\ : std_logic;
signal \ALU.r0_12_prm_8_12_s0_c_RNOZ0\ : std_logic;
signal \ALU.lshift_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.r4_RNI1RK3KZ0Z_9\ : std_logic;
signal \ALU.r4_RNIOK1781Z0Z_9_cascade_\ : std_logic;
signal \ALU.lshift_11\ : std_logic;
signal \ALU.r5_RNI27VE5Z0Z_10\ : std_logic;
signal \ALU.un2_addsub_cry_12_c_RNI74A7EZ0\ : std_logic;
signal \ALU.r0_12_prm_2_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.rshift_11\ : std_logic;
signal \ALU.r0_12_prm_8_10_s1_c_RNOZ0Z_1\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \ALU.r0_12_prm_8_10_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNIUF9K8_0Z0Z_10\ : std_logic;
signal \ALU.r0_12_prm_8_10_s1\ : std_logic;
signal \ALU.r0_12_prm_6_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_10\ : std_logic;
signal \ALU.r0_12_prm_7_10_s1\ : std_logic;
signal \ALU.r0_12_prm_5_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNIUF9K8_1Z0Z_10\ : std_logic;
signal \ALU.r0_12_prm_6_10_s1\ : std_logic;
signal \ALU.r0_12_prm_4_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_10\ : std_logic;
signal \ALU.r0_12_prm_5_10_s1\ : std_logic;
signal \ALU.r0_12_prm_4_10_s1\ : std_logic;
signal \ALU.r0_12_prm_2_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_10_s1\ : std_logic;
signal \ALU.r0_12_prm_2_10_s1\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \ALU.r0_12_s1_10\ : std_logic;
signal \ALU.r0_12_s1_10_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_1_13_s0_c_RNOZ0\ : std_logic;
signal \bfn_11_1_0_\ : std_logic;
signal \ALU.r0_12_prm_8_6_s1_c_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_7_6_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_6_s1\ : std_logic;
signal \ALU.r0_12_prm_6_6_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_6_s1\ : std_logic;
signal \ALU.r0_12_prm_5_6_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_6_s1\ : std_logic;
signal \ALU.r0_12_prm_4_6_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_6_s1\ : std_logic;
signal \ALU.r0_12_prm_4_6_s1\ : std_logic;
signal \ALU.r0_12_prm_2_6_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_6_s1\ : std_logic;
signal \ALU.r0_12_prm_2_6_s1\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \ALU.r0_12_s1_6\ : std_logic;
signal \ALU.lshift_6_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_6_s1_c_RNOZ0\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \ALU.r0_12_prm_7_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_0_s0\ : std_logic;
signal \ALU.r0_12_prm_6_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_0_s0\ : std_logic;
signal \ALU.r0_12_prm_5_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_0_s0\ : std_logic;
signal \ALU.r2_RNIKG5N5Z0Z_0\ : std_logic;
signal \ALU.r0_12_prm_5_0_s0\ : std_logic;
signal \ALU.r0_12_prm_3_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_4_0_s0\ : std_logic;
signal \ALU.r0_12_prm_3_0_s0\ : std_logic;
signal \ALU.r0_12_prm_1_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_2_0_s0\ : std_logic;
signal \ALU.r0_12_s0_0\ : std_logic;
signal \ALU.rshift_0\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal r1_0 : std_logic;
signal \ALU.lshift_3_ns_1_8_cascade_\ : std_logic;
signal \ALU.r4_RNILIPV9Z0Z_6_cascade_\ : std_logic;
signal \ALU.r4_RNI1G9PKZ0Z_6_cascade_\ : std_logic;
signal r0_1 : std_logic;
signal r0_3 : std_logic;
signal \ALU.r0_12_0\ : std_logic;
signal r0_0 : std_logic;
signal \ALU.r5_RNI9S2TIZ0Z_11_cascade_\ : std_logic;
signal \ALU.lshift_15_ns_1_13_cascade_\ : std_logic;
signal \ALU.un9_addsub_axb_2\ : std_logic;
signal \ALU.un14_log_0_i_11\ : std_logic;
signal \ALU.a6_b_0\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \ALU.r4_RNI90J9EZ0Z_1\ : std_logic;
signal \ALU.un9_addsub_cry_0\ : std_logic;
signal \ALU.r4_RNI468UDZ0Z_2\ : std_logic;
signal \ALU.un9_addsub_cry_1\ : std_logic;
signal \ALU.r4_RNIUU8UDZ0Z_3\ : std_logic;
signal \ALU.un9_addsub_cry_2\ : std_logic;
signal \ALU.r4_RNIQK1EDZ0Z_4\ : std_logic;
signal \ALU.un9_addsub_cry_3\ : std_logic;
signal \ALU.un9_addsub_cry_4\ : std_logic;
signal \ALU.un9_addsub_cry_5\ : std_logic;
signal \ALU.un9_addsub_cry_6\ : std_logic;
signal \ALU.un9_addsub_cry_7\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \ALU.un9_addsub_cry_8\ : std_logic;
signal \ALU.un9_addsub_cry_9\ : std_logic;
signal \ALU.b_11\ : std_logic;
signal \ALU.un9_addsub_cry_10\ : std_logic;
signal \ALU.un9_addsub_cry_11\ : std_logic;
signal \ALU.b_13\ : std_logic;
signal \ALU.un9_addsub_cry_12_c_RNISR30AZ0\ : std_logic;
signal \ALU.un9_addsub_cry_12\ : std_logic;
signal \ALU.un9_addsub_cry_13\ : std_logic;
signal \ALU.un9_addsub_cry_14\ : std_logic;
signal \ALU.r0_12_prm_6_10_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_13_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_2_12_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_1_9_s0_c_RNOZ0\ : std_logic;
signal \ALU.lshift_3_ns_1_13\ : std_logic;
signal \ALU.rshift_12\ : std_logic;
signal \ALU.un2_addsub_cry_9_c_RNIS67KDZ0\ : std_logic;
signal \ALU.r0_12_prm_2_10_s0_c_RNOZ0\ : std_logic;
signal \ALU.un2_addsub_cry_10_c_RNIS4T7DZ0\ : std_logic;
signal \ALU.r0_12_prm_2_11_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNIAP7U9Z0Z_10\ : std_logic;
signal \ALU.r5_RNIKU3HJZ0Z_10_cascade_\ : std_logic;
signal \ALU.r4_RNIQK1V71Z0Z_5_cascade_\ : std_logic;
signal \ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09\ : std_logic;
signal \ALU.r0_12_prm_1_11_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_2_14_s0_c_RNOZ0\ : std_logic;
signal \ALU.rshift_15\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \ALU.lshift_15\ : std_logic;
signal \ALU.r0_12_prm_8_15_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_15_s0_cy\ : std_logic;
signal \ALU.r2_RNI7AQC9_0Z0Z_15\ : std_logic;
signal \ALU.r0_12_prm_8_15_s0\ : std_logic;
signal \ALU.r0_12_prm_6_15_s0_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_15\ : std_logic;
signal \ALU.r0_12_prm_7_15_s0\ : std_logic;
signal \ALU.r0_12_prm_5_15_s0_c_RNOZ0\ : std_logic;
signal \ALU.r2_RNI7AQC9_1Z0Z_15\ : std_logic;
signal \ALU.r0_12_prm_6_15_s0\ : std_logic;
signal \ALU.r5_RNI5P1F5Z0Z_15\ : std_logic;
signal \ALU.a_i_15\ : std_logic;
signal \ALU.r0_12_prm_5_15_s0\ : std_logic;
signal \ALU.r0_12_prm_3_15_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_15_s0\ : std_logic;
signal \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9\ : std_logic;
signal \ALU.r0_12_prm_2_15_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_15_s0\ : std_logic;
signal \ALU.r0_12_prm_2_15_s0\ : std_logic;
signal \ALU.r0_12_prm_1_15_s0_c_RNOZ0\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \ALU.r0_12_s0_15\ : std_logic;
signal \ALU.r0_12_s0_15_THRU_CO\ : std_logic;
signal \ALU.r5_RNIB8HG5Z0Z_12\ : std_logic;
signal \ALU.lshift_13\ : std_logic;
signal \ALU.r0_12_prm_8_13_s1_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8\ : std_logic;
signal \ALU.r0_12_prm_1_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_1_12_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_1_6_s1_c_RNOZ0\ : std_logic;
signal \ALU.rshift_3_ns_1_4_cascade_\ : std_logic;
signal \bfn_12_2_0_\ : std_logic;
signal \ALU.r0_12_prm_7_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_0_s1\ : std_logic;
signal \ALU.r0_12_prm_6_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_0\ : std_logic;
signal \ALU.r0_12_prm_7_0_s1\ : std_logic;
signal \ALU.r0_12_prm_5_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_0_s1\ : std_logic;
signal \ALU.r0_12_prm_4_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.N_883_i\ : std_logic;
signal \ALU.r0_12_prm_5_0_s1\ : std_logic;
signal \ALU.r0_12_prm_3_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.mult_0\ : std_logic;
signal \ALU.r0_12_prm_4_0_s1\ : std_logic;
signal \ALU.r0_12_prm_3_0_s1\ : std_logic;
signal \ALU.r0_12_prm_1_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_axb_0\ : std_logic;
signal \ALU.r0_12_prm_2_0_s1\ : std_logic;
signal \ALU.r0_12_s1_0\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \ALU.r0_12_s1_0_THRU_CO\ : std_logic;
signal \ALU.rshift_15_ns_1_0\ : std_logic;
signal \ALU.r0_12_prm_2_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.rshift_15_ns_1_6\ : std_logic;
signal \ALU.rshift_3_ns_1_5\ : std_logic;
signal \ALU.r4_RNI9OH6AZ0Z_1_cascade_\ : std_logic;
signal \ALU.r5_RNIVQN52Z0Z_10\ : std_logic;
signal \ALU.r6_RNIP3372Z0Z_10\ : std_logic;
signal \a_1_repZ0Z2\ : std_logic;
signal \ALU.a10_b_4\ : std_logic;
signal \ALU.lshift_3_ns_1_5\ : std_logic;
signal \ALU.lshift_15_ns_1_9\ : std_logic;
signal \ALU.r4_RNIF01FKZ0Z_2_cascade_\ : std_logic;
signal \ALU.r4_RNI2H9PKZ0Z_6\ : std_logic;
signal \ALU.lshift_9_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_9_s0_c_RNOZ0\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \ALU.r0_12_prm_8_7_s0_c_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_8_7_s0\ : std_logic;
signal \ALU.r0_12_prm_6_7_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_7_s0\ : std_logic;
signal \ALU.r0_12_prm_6_7_s0\ : std_logic;
signal \ALU.r4_RNIFR136Z0Z_7\ : std_logic;
signal \ALU.r0_12_prm_5_7_s0\ : std_logic;
signal \ALU.r0_12_prm_3_7_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_7_s0\ : std_logic;
signal \ALU.r0_12_prm_3_7_s0\ : std_logic;
signal \ALU.r0_12_prm_2_7_s0\ : std_logic;
signal \ALU.r0_12_prm_1_7_s0_c_RNOZ0\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \ALU.mult_7\ : std_logic;
signal \ALU.r0_12_s0_7\ : std_logic;
signal r1_7 : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \ALU.r0_12_prm_8_5_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_7_5_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_5_s0\ : std_logic;
signal \ALU.r0_12_prm_6_5_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_5_s0\ : std_logic;
signal \ALU.r0_12_prm_5_5_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_5_s0\ : std_logic;
signal \ALU.r4_RNIM8HG5Z0Z_5\ : std_logic;
signal \ALU.r0_12_prm_5_5_s0\ : std_logic;
signal \ALU.r0_12_prm_3_5_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_5_s0\ : std_logic;
signal \ALU.r0_12_prm_2_5_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_5_s0\ : std_logic;
signal \ALU.r0_12_prm_2_5_s0\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \ALU.mult_5\ : std_logic;
signal \ALU.r0_12_s0_5\ : std_logic;
signal \ALU.r0_12_5\ : std_logic;
signal r1_5 : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \ALU.r0_12_prm_8_8_s0_cy\ : std_logic;
signal \ALU.r0_12_prm_8_8_s0\ : std_logic;
signal \ALU.r0_12_prm_6_8_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_8_s0\ : std_logic;
signal \ALU.r0_12_prm_6_8_s0\ : std_logic;
signal \ALU.r0_12_prm_5_8_s0\ : std_logic;
signal \ALU.r0_12_prm_3_8_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_8_s0\ : std_logic;
signal \ALU.r0_12_prm_3_8_s0\ : std_logic;
signal \ALU.r0_12_prm_2_8_s0\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \ALU.r0_12_s0_8\ : std_logic;
signal \ALU.r0_12_prm_1_8_s0_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9\ : std_logic;
signal \ALU.r0_12_prm_1_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNIQK1V71Z0Z_5\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \ALU.r0_12_prm_8_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.lshift_12\ : std_logic;
signal \ALU.r0_12_prm_8_12_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNISP2L9_0Z0Z_12\ : std_logic;
signal \ALU.r0_12_prm_8_12_s1\ : std_logic;
signal \ALU.un14_log_0_i_12\ : std_logic;
signal \ALU.r0_12_prm_7_12_s1\ : std_logic;
signal \ALU.r0_12_prm_5_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNISP2L9_1Z0Z_12\ : std_logic;
signal \ALU.r0_12_prm_6_12_s1\ : std_logic;
signal \ALU.r0_12_prm_4_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_12\ : std_logic;
signal \ALU.r0_12_prm_5_12_s1\ : std_logic;
signal \ALU.r0_12_prm_4_12_s1\ : std_logic;
signal \ALU.un2_addsub_cry_11_c_RNICP8AEZ0\ : std_logic;
signal \ALU.r0_12_prm_2_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_12_s1\ : std_logic;
signal \ALU.r0_12_prm_2_12_s1\ : std_logic;
signal \ALU.r0_12_prm_1_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_11_c_RNIAHI1AZ0\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \ALU.r0_12_s1_12\ : std_logic;
signal \ALU.r0_12_s1_12_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_5_15_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_15_s1_c_RNOZ0Z_1\ : std_logic;
signal \ALU.r0_12_prm_8_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNIAV175Z0Z_15\ : std_logic;
signal \ALU.r0_12_prm_2_0_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_2_c_RNOZ0Z_3\ : std_logic;
signal \ALU.r4_RNI1G9PKZ0Z_6\ : std_logic;
signal \ALU.N_845_1\ : std_logic;
signal \ALU.rshift_15_ns_1_2_cascade_\ : std_logic;
signal \ALU.r5_RNI8R2TIZ0Z_11\ : std_logic;
signal \ALU.bZ0Z_0\ : std_logic;
signal \ALU.r4_RNID26E8_0Z0Z_0\ : std_logic;
signal \ALU.rshift_6\ : std_logic;
signal \bfn_13_3_0_\ : std_logic;
signal \ALU.lshift_6\ : std_logic;
signal \ALU.r0_12_prm_8_6_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_6_s0_c_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_8_6_s0\ : std_logic;
signal \ALU.un14_log_0_i_6\ : std_logic;
signal \ALU.r0_12_prm_7_6_s0\ : std_logic;
signal \ALU.r4_RNI2BKQ8_0Z0Z_6\ : std_logic;
signal \ALU.r0_12_prm_6_6_s0\ : std_logic;
signal \ALU.r4_RNIUGHG5Z0Z_6\ : std_logic;
signal \ALU.a_i_6\ : std_logic;
signal \ALU.r0_12_prm_5_6_s0\ : std_logic;
signal \ALU.r0_12_prm_3_6_s0_sf\ : std_logic;
signal \ALU.r0_12_prm_4_6_s0\ : std_logic;
signal \ALU.un2_addsub_cry_5_c_RNIO30SDZ0\ : std_logic;
signal \ALU.r0_12_prm_2_6_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_6_s0\ : std_logic;
signal \ALU.r0_12_prm_2_6_s0\ : std_logic;
signal \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019\ : std_logic;
signal \ALU.r0_12_prm_1_6_s0_c_RNOZ0\ : std_logic;
signal \bfn_13_4_0_\ : std_logic;
signal \ALU.r0_12_s1_6_THRU_CO\ : std_logic;
signal \ALU.mult_6\ : std_logic;
signal \ALU.r0_12_s0_6\ : std_logic;
signal r1_6 : std_logic;
signal \bfn_13_5_0_\ : std_logic;
signal \ALU.r0_12_prm_8_4_c_THRU_CO\ : std_logic;
signal \ALU.a4_b_4\ : std_logic;
signal \ALU.r0_12_prm_7_4_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_4\ : std_logic;
signal \ALU.r0_12_prm_6_4_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_4\ : std_logic;
signal \ALU.r0_12_prm_7_4\ : std_logic;
signal \ALU.r0_12_prm_5_4_c_RNOZ0Z_0\ : std_logic;
signal \ALU.r0_12_prm_6_4\ : std_logic;
signal \ALU.a_i_4\ : std_logic;
signal \ALU.r0_12_prm_5_4\ : std_logic;
signal \ALU.mult_4\ : std_logic;
signal \ALU.r0_12_prm_4_4\ : std_logic;
signal \ALU.r0_12_prm_3_4\ : std_logic;
signal \ALU.r0_12_prm_2_4\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \ALU.r0_12_4\ : std_logic;
signal \ALU.r5_RNIKS4A9Z0Z_11\ : std_logic;
signal \ALU.r4_RNIVLAIAZ0Z_9\ : std_logic;
signal \ALU.r5_RNI0QK3KZ0Z_11_cascade_\ : std_logic;
signal \ALU.rshift_8\ : std_logic;
signal \ALU.un2_addsub_cry_3_c_RNI8MVBGZ0\ : std_logic;
signal \ALU.r0_12_prm_2_4_c_RNOZ0\ : std_logic;
signal \ALU.madd_axb_3\ : std_logic;
signal \ALU.madd_cry_2_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_3_4_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_2_7_s0_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNIODO6KZ0Z_5\ : std_logic;
signal \ALU.lshift_8_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_8_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_12_s1_c_RNOZ0Z_1\ : std_logic;
signal \ALU.r0_12_prm_7_8_s0_c_RNOZ0\ : std_logic;
signal \ALU.rshift_5\ : std_logic;
signal \ALU.r0_12_6\ : std_logic;
signal r6_6 : std_logic;
signal \ALU.r0_12_7\ : std_logic;
signal r6_7 : std_logic;
signal r6_8 : std_logic;
signal r6_2 : std_logic;
signal r6_3 : std_logic;
signal \ALU.r0_12_4_THRU_CO\ : std_logic;
signal r6_4 : std_logic;
signal \ALU.r4_RNIN3236Z0Z_8\ : std_logic;
signal \ALU.rshift_3_ns_1_1\ : std_logic;
signal \ALU.r0_12_prm_8_1_c_RNOZ0Z_3_cascade_\ : std_logic;
signal \ALU.rshift_15_ns_1_1_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_8_s1_c_RNOZ0Z_1\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \ALU.lshift_8\ : std_logic;
signal \ALU.r0_12_prm_8_8_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_8_s1_cy\ : std_logic;
signal \ALU.a8_b_8\ : std_logic;
signal \ALU.r0_12_prm_8_8_s1\ : std_logic;
signal \ALU.un14_log_0_i_8\ : std_logic;
signal \ALU.r0_12_prm_7_8_s1\ : std_logic;
signal \ALU.r0_12_prm_6_8_s1\ : std_logic;
signal \ALU.r0_12_prm_4_8_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_8\ : std_logic;
signal \ALU.r0_12_prm_5_8_s1\ : std_logic;
signal \ALU.r0_12_prm_4_8_s1\ : std_logic;
signal \ALU.r0_12_prm_2_8_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_8_s1\ : std_logic;
signal \ALU.r0_12_prm_2_8_s1\ : std_logic;
signal \ALU.un9_addsub_cry_7_c_RNINZ0Z3519\ : std_logic;
signal \ALU.r0_12_prm_1_8_s1_c_RNOZ0\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \ALU.madd_cry_6_THRU_CO\ : std_logic;
signal \ALU.madd_axb_7\ : std_logic;
signal \ALU.r0_12_s0_8_THRU_CO\ : std_logic;
signal \ALU.r0_12_s1_8\ : std_logic;
signal \ALU.r0_12_8\ : std_logic;
signal r0_8 : std_logic;
signal \ALU.un2_addsub_cry_7_c_RNI5ELEEZ0\ : std_logic;
signal \ALU.r0_12_prm_2_8_s0_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNITTMB9Z0Z_12\ : std_logic;
signal \ALU.r5_RNITTMB9Z0Z_12_cascade_\ : std_logic;
signal \ALU.r5_RNITG1F5Z0Z_14\ : std_logic;
signal \ALU.r0_12_prm_5_14_s0_c_RNOZ0\ : std_logic;
signal \ALU.rshift_13\ : std_logic;
signal \ALU.r0_12_prm_6_14_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_14_s0_c_RNOZ0\ : std_logic;
signal \ALU.a_15\ : std_logic;
signal \ALU.b_15\ : std_logic;
signal \ALU.r0_12_prm_7_15_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_13_s1_c_RNOZ0Z_1\ : std_logic;
signal \ALU.b_12\ : std_logic;
signal \ALU.r0_12_prm_6_12_s1_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNIPV8A9_0Z0Z_13\ : std_logic;
signal \ALU.rshift_2\ : std_logic;
signal \bfn_14_1_0_\ : std_logic;
signal \ALU.r0_12_prm_8_2_c_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_8_2\ : std_logic;
signal \ALU.r0_12_prm_7_2\ : std_logic;
signal \ALU.r0_12_prm_5_2_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_2\ : std_logic;
signal \ALU.r4_RNIL9636Z0Z_2\ : std_logic;
signal \ALU.a_i_2\ : std_logic;
signal \ALU.r0_12_prm_5_2\ : std_logic;
signal \ALU.r0_12_prm_4_2\ : std_logic;
signal \ALU.r0_12_prm_3_2\ : std_logic;
signal \ALU.r0_12_prm_2_2\ : std_logic;
signal \bfn_14_2_0_\ : std_logic;
signal \ALU.r0_12_2\ : std_logic;
signal \ALU.r0_12_2_THRU_CO\ : std_logic;
signal \ALU.lshift_2\ : std_logic;
signal \ALU.r0_12_prm_8_2_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_0_s0_c_RNOZ0\ : std_logic;
signal \ALU.a2_b_2\ : std_logic;
signal \ALU.r0_12_prm_7_2_c_RNOZ0\ : std_logic;
signal \ALU.lshift_0\ : std_logic;
signal \ALU.r4_RNIHENK8_1Z0Z_7\ : std_logic;
signal \ALU.b_i_0\ : std_logic;
signal \ALU.un2_addsub_axb_0_i\ : std_logic;
signal \ALU.un2_addsub_cry_1_c_RNI1H7SGZ0\ : std_logic;
signal \ALU.r0_12_prm_2_2_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_2_c_RNOZ0\ : std_logic;
signal \ALU.b_4\ : std_logic;
signal \ALU.r0_12_prm_5_4_c_RNOZ0\ : std_logic;
signal \ALU.rshift_3_ns_1_9_cascade_\ : std_logic;
signal \ALU.a_11\ : std_logic;
signal \ALU.r0_12_prm_5_8_s0_c_RNOZ0\ : std_logic;
signal \ALU.N_610_1_cascade_\ : std_logic;
signal \ALU.r4_RNIVFRGQ_0Z0Z_2_cascade_\ : std_logic;
signal \ALU.lshift_4\ : std_logic;
signal \ALU.r0_12_prm_6_6_s0_c_RNOZ0\ : std_logic;
signal \ALU.a_13\ : std_logic;
signal \ALU.a_12\ : std_logic;
signal \ALU.r4_RNI9H7SJZ0Z_6\ : std_logic;
signal \ALU.r5_RNI0QK3KZ0Z_11\ : std_logic;
signal \ALU.r0_12_prm_8_4_c_RNOZ0Z_2_cascade_\ : std_logic;
signal \ALU.rshift_4\ : std_logic;
signal \ALU.lshift_15_ns_1_8\ : std_logic;
signal \ALU.lshift_3_ns_1_4\ : std_logic;
signal \ALU.r4_RNI6PL1LZ0Z_2\ : std_logic;
signal \ALU.r4_RNI6PL1LZ0Z_2_cascade_\ : std_logic;
signal \ALU.r4_RNIVFRGQZ0Z_2\ : std_logic;
signal \ALU.r4_RNIVFRGQ_0Z0Z_2\ : std_logic;
signal \ALU.r0_12_prm_8_4_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNIODO6KZ0Z_7\ : std_logic;
signal \ALU.r0_12_prm_8_4_c_RNOZ0Z_3\ : std_logic;
signal \ALU.un9_addsub_cry_3_c_RNIV8DFIZ0\ : std_logic;
signal \ALU.r0_12_prm_1_4_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNI7NOB9Z0Z_13\ : std_logic;
signal \ALU.r5_RNIUE7TIZ0Z_13\ : std_logic;
signal \ALU.r4_RNIRL1V71Z0Z_7\ : std_logic;
signal \ALU.a6_b_6\ : std_logic;
signal \ALU.r0_12_prm_7_6_s0_c_RNOZ0\ : std_logic;
signal \ALU.rshift_1\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \ALU.lshift_1\ : std_logic;
signal \ALU.r0_12_prm_8_1_c_THRU_CO\ : std_logic;
signal \ALU.a1_b_1\ : std_logic;
signal \ALU.r0_12_prm_7_1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_1\ : std_logic;
signal \ALU.r0_12_prm_6_1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_1\ : std_logic;
signal \ALU.r0_12_prm_5_1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_1\ : std_logic;
signal \ALU.r4_RNID1636Z0Z_1\ : std_logic;
signal \ALU.a_i_1\ : std_logic;
signal \ALU.r0_12_prm_5_1\ : std_logic;
signal \ALU.r0_12_prm_3_1_c_RNOZ0\ : std_logic;
signal \ALU.mult_1\ : std_logic;
signal \ALU.r0_12_prm_4_1\ : std_logic;
signal \ALU.r0_12_prm_3_1\ : std_logic;
signal \ALU.r0_12_prm_2_1\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \ALU.r0_12_1\ : std_logic;
signal \ALU.r0_12_1_THRU_CO\ : std_logic;
signal \ALU.un9_addsub_cry_0_c_RNIG8GLJZ0\ : std_logic;
signal \ALU.r0_12_prm_1_1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_9_s0_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNIKUMQ8_0Z0Z_8\ : std_logic;
signal \ALU.r0_12_prm_6_8_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_10_s0_c_RNOZ0\ : std_logic;
signal \ALU.lshift_3_ns_1_10\ : std_logic;
signal \ALU.r4_RNI67NNKZ0Z_7_cascade_\ : std_logic;
signal \ALU.lshift_10\ : std_logic;
signal \ALU.N_610_1\ : std_logic;
signal \ALU.r4_RNIAHIIAZ0Z_2\ : std_logic;
signal \ALU.r4_RNI38O1GZ0Z_2\ : std_logic;
signal \ALU.r4_RNI38O1GZ0Z_2_cascade_\ : std_logic;
signal \ALU.r4_RNICN8R81Z0Z_7\ : std_logic;
signal \ALU.r0_12_prm_8_10_s1_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNI67NNKZ0Z_7\ : std_logic;
signal \ALU.r5_RNI355TIZ0Z_13\ : std_logic;
signal \ALU.r4_RNIO7CSJZ0Z_4\ : std_logic;
signal \ALU.lshift_15_ns_1_14_cascade_\ : std_logic;
signal \ALU.r4_RNILVIQFZ0Z_2\ : std_logic;
signal \ALU.r0_12_prm_8_9_s1_c_RNOZ0Z_1\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \ALU.r0_12_prm_8_9_s1_c_RNOZ0\ : std_logic;
signal \ALU.lshift_9\ : std_logic;
signal \ALU.r0_12_prm_8_9_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_9_s1_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNISU5D9_0Z0Z_9\ : std_logic;
signal \ALU.r0_12_prm_8_9_s1\ : std_logic;
signal \ALU.r0_12_prm_6_9_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_9_s1\ : std_logic;
signal \ALU.r4_RNISU5D9_1Z0Z_9\ : std_logic;
signal \ALU.r0_12_prm_5_9_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_9_s1\ : std_logic;
signal \ALU.a_i_9\ : std_logic;
signal \ALU.r0_12_prm_5_9_s1\ : std_logic;
signal \ALU.r0_12_prm_4_9_s1\ : std_logic;
signal \ALU.r0_12_prm_2_9_s1_c_RNOZ0\ : std_logic;
signal \ALU.un2_addsub_cry_8_c_RNINO51FZ0\ : std_logic;
signal \ALU.r0_12_prm_3_9_s1\ : std_logic;
signal \ALU.r0_12_prm_2_9_s1\ : std_logic;
signal \ALU.r0_12_prm_1_9_s1_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \ALU.r0_12_s1_9\ : std_logic;
signal \ALU.r0_12_s1_9_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_7_14_s0_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_2\ : std_logic;
signal \ALU.mult_2\ : std_logic;
signal \ALU.madd_cry_0_THRU_CO\ : std_logic;
signal \ALU.madd_axb_1\ : std_logic;
signal \ALU.r0_12_prm_3_2_c_RNOZ0\ : std_logic;
signal \ALU.a_4\ : std_logic;
signal \ALU.r4_RNI87HO5Z0Z_4\ : std_logic;
signal \ALU.b_2\ : std_logic;
signal \ALU.r0_12_prm_5_2_c_RNOZ0Z_0\ : std_logic;
signal \ALU.un9_addsub_cry_1_c_RNIKO6AJZ0\ : std_logic;
signal \ALU.r0_12_prm_1_2_c_RNOZ0\ : std_logic;
signal \ALU.b_6\ : std_logic;
signal \ALU.a_6\ : std_logic;
signal \ALU.r0_12_prm_5_6_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_7_s0_c_RNOZ0\ : std_logic;
signal \ALU.r5_RNILM5AEZ0Z_15\ : std_logic;
signal \ALU.r5_RNILV3HJZ0Z_12\ : std_logic;
signal \ALU.rshift_9\ : std_logic;
signal \ALU.r4_RNI9H7SJZ0Z_5\ : std_logic;
signal \ALU.lshift_7_cascade_\ : std_logic;
signal \ALU.r0_12_prm_8_7_s0_c_RNOZ0\ : std_logic;
signal \ALU.rshift_7\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \ALU.r0_12_prm_8_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.lshift_7\ : std_logic;
signal \ALU.r0_12_prm_8_7_s1_c_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_8_7_s1\ : std_logic;
signal \ALU.un14_log_0_i_7\ : std_logic;
signal \ALU.r0_12_prm_7_7_s1\ : std_logic;
signal \ALU.r0_12_prm_5_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNIHENK8_0Z0Z_7\ : std_logic;
signal \ALU.r0_12_prm_6_7_s1\ : std_logic;
signal \ALU.r0_12_prm_4_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_7\ : std_logic;
signal \ALU.r0_12_prm_5_7_s1\ : std_logic;
signal \ALU.r0_12_prm_4_7_s1\ : std_logic;
signal \ALU.un2_addsub_cry_6_c_RNIPJK8EZ0\ : std_logic;
signal \ALU.r0_12_prm_2_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_7_s1\ : std_logic;
signal \ALU.r0_12_prm_2_7_s1\ : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal \ALU.r0_12_s1_7\ : std_logic;
signal \ALU.r0_12_s1_7_THRU_CO\ : std_logic;
signal \ALU.r5_RNISMSV4Z0Z_15\ : std_logic;
signal \ALU.rshift_15_ns_1_3\ : std_logic;
signal \ALU.r5_RNI465TIZ0Z_13\ : std_logic;
signal \ALU.r4_RNIF01FKZ0Z_2\ : std_logic;
signal \ALU.b_7\ : std_logic;
signal \ALU.a_7\ : std_logic;
signal \ALU.r0_12_prm_6_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.b_3\ : std_logic;
signal \ALU.r0_12_prm_1_5_s0_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_9\ : std_logic;
signal \ALU.a_5\ : std_logic;
signal \ALU.b_5\ : std_logic;
signal \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8\ : std_logic;
signal \ALU.r0_12_prm_1_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_5_s1_c_RNOZ0Z_1\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \ALU.r0_12_prm_8_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_5_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_8_5_s1\ : std_logic;
signal \ALU.r0_12_prm_6_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_5\ : std_logic;
signal \ALU.r0_12_prm_7_5_s1\ : std_logic;
signal \ALU.r4_RNI8B628_0Z0Z_5\ : std_logic;
signal \ALU.r0_12_prm_5_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_6_5_s1\ : std_logic;
signal \ALU.r0_12_prm_4_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_5\ : std_logic;
signal \ALU.r0_12_prm_5_5_s1\ : std_logic;
signal \ALU.r0_12_prm_4_5_s1\ : std_logic;
signal \ALU.r0_12_prm_2_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.un2_addsub_cry_4_c_RNILPG3DZ0\ : std_logic;
signal \ALU.r0_12_prm_3_5_s1\ : std_logic;
signal \ALU.r0_12_prm_2_5_s1\ : std_logic;
signal \ALU.r0_12_prm_1_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \ALU.r0_12_s1_5\ : std_logic;
signal \ALU.r0_12_s1_5_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_5_8_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_10_s0_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_1_c_RNOZ0Z_0\ : std_logic;
signal \ALU.rshift_14\ : std_logic;
signal \ALU.N_622_1\ : std_logic;
signal \ALU.r0_12_prm_8_1_c_RNOZ0\ : std_logic;
signal \ALU.b_8\ : std_logic;
signal \ALU.a_8\ : std_logic;
signal \ALU.r0_12_prm_7_8_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_9_s0_c_RNOZ0\ : std_logic;
signal \ALU.un1_yindexZ0Z_1\ : std_logic;
signal \ALU.un1_yindexZ0Z_2\ : std_logic;
signal \ALU.un1_yindexZ0Z_3\ : std_logic;
signal \ALU.un1_yindexZ0Z_4\ : std_logic;
signal \ALU.un1_yindexZ0Z_5\ : std_logic;
signal \ALU.un1_yindexZ0Z_6\ : std_logic;
signal \ALU.un1_yindexZ0Z_7\ : std_logic;
signal \ALU.b_9\ : std_logic;
signal \ALU.r4_RNISU5D9_2Z0Z_9\ : std_logic;
signal \ALU.a5_b_5\ : std_logic;
signal \ALU.r0_12_prm_7_5_s1_c_RNOZ0\ : std_logic;
signal \ALU.b_14\ : std_logic;
signal \ALU.a_14\ : std_logic;
signal \ALU.r0_12_prm_7_7_s1_c_RNOZ0\ : std_logic;
signal \ALU.b_1\ : std_logic;
signal \ALU.un14_log_0_i_1\ : std_logic;
signal \ALU.a7_b_7\ : std_logic;
signal \ALU.r0_12_prm_7_7_s0_c_RNOZ0\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \ALU.r0_12_prm_8_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.lshift_14\ : std_logic;
signal \ALU.r0_12_prm_8_14_s1_cy\ : std_logic;
signal \ALU.r0_12_prm_7_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.r2_RNINPPC9_0Z0Z_14\ : std_logic;
signal \ALU.r0_12_prm_8_14_s1\ : std_logic;
signal \ALU.r0_12_prm_6_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.un14_log_0_i_14\ : std_logic;
signal \ALU.r0_12_prm_7_14_s1\ : std_logic;
signal \ALU.r0_12_prm_5_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.r2_RNINPPC9_1Z0Z_14\ : std_logic;
signal \ALU.r0_12_prm_6_14_s1\ : std_logic;
signal \ALU.r0_12_prm_4_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.a_i_14\ : std_logic;
signal \ALU.r0_12_prm_5_14_s1\ : std_logic;
signal \ALU.r0_12_prm_4_14_s1\ : std_logic;
signal \ALU.un2_addsub_cry_13_c_RNIR5I0EZ0\ : std_logic;
signal \ALU.r0_12_prm_2_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_14_s1\ : std_logic;
signal \ALU.r0_12_prm_2_14_s1\ : std_logic;
signal \ALU.r0_12_prm_1_14_s1_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \ALU.r0_12_s1_14\ : std_logic;
signal \ALU.r0_12_s1_14_THRU_CO\ : std_logic;
signal \ALU.aZ0Z_0\ : std_logic;
signal \ALU.a_1\ : std_logic;
signal \ALU.a_2\ : std_logic;
signal \ALU.rshift_3_ns_1_0_cascade_\ : std_logic;
signal \ALU.r4_RNII2A0LZ0Z_2\ : std_logic;
signal \ALU.lshift_5\ : std_logic;
signal \ALU.r0_12_prm_8_5_s0_c_RNOZ0\ : std_logic;
signal \ALU.r4_RNI0C236Z0Z_9\ : std_logic;
signal \ALU.rshift_3\ : std_logic;
signal \bfn_16_5_0_\ : std_logic;
signal \ALU.r0_12_prm_8_3_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_8_3_c_THRU_CO\ : std_logic;
signal \ALU.r0_12_prm_7_3_c_RNOZ0\ : std_logic;
signal \ALU.a3_b_3\ : std_logic;
signal \ALU.r0_12_prm_8_3\ : std_logic;
signal \ALU.un14_log_0_i_3\ : std_logic;
signal \ALU.r0_12_prm_6_3_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_7_3\ : std_logic;
signal \ALU.r0_12_prm_5_3_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_5_3_c_RNOZ0Z_0\ : std_logic;
signal \ALU.r0_12_prm_6_3\ : std_logic;
signal \ALU.r4_RNIUH636Z0Z_3\ : std_logic;
signal \ALU.a_3\ : std_logic;
signal \ALU.a_i_3\ : std_logic;
signal \ALU.r0_12_prm_5_3\ : std_logic;
signal \ALU.r0_12_prm_4_3\ : std_logic;
signal \ALU.r0_12_prm_3_3\ : std_logic;
signal \ALU.r0_12_prm_2_3\ : std_logic;
signal \ALU.r0_12_prm_1_3_c_RNOZ0\ : std_logic;
signal \ALU.un9_addsub_cry_2_c_RNIOR8AJZ0\ : std_logic;
signal \bfn_16_6_0_\ : std_logic;
signal \ALU.r0_12_3\ : std_logic;
signal \ALU.r0_12_3_THRU_CO\ : std_logic;
signal \ALU.un2_addsub_cry_2_c_RNI3K9SGZ0\ : std_logic;
signal \ALU.r0_12_prm_2_3_c_RNOZ0\ : std_logic;
signal \ALU.r0_12_prm_3_3_c_RNOZ0\ : std_logic;
signal \ALU.madd_axb_2\ : std_logic;
signal \ALU.madd_cry_1_THRU_CO\ : std_logic;
signal \ALU.mult_3\ : std_logic;
signal \TXbuffer_RNO_1Z0Z_7\ : std_logic;
signal \TXbuffer_RNO_0Z0Z_7\ : std_logic;
signal \clkdivZ0Z_4\ : std_logic;
signal \TXbuffer_18_15_ns_1_7\ : std_logic;
signal \yZ0Z_2\ : std_logic;
signal \ALU.un1_yindexZ0Z_8\ : std_logic;
signal \yZ0Z_0\ : std_logic;
signal \yZ0Z_1\ : std_logic;
signal \TXbufferZ0Z_7\ : std_logic;
signal \INVFTDI.TXshift_7C_net\ : std_logic;
signal \TXbufferZ0Z_1\ : std_logic;
signal \TXbufferZ0Z_2\ : std_logic;
signal \FTDI.TXshiftZ0Z_2\ : std_logic;
signal \INVFTDI.TXshift_1C_net\ : std_logic;
signal \TXbufferZ0Z_4\ : std_logic;
signal \FTDI.TXshiftZ0Z_4\ : std_logic;
signal \TXbufferZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_7\ : std_logic;
signal \TXbufferZ0Z_6\ : std_logic;
signal \FTDI.TXshiftZ0Z_6\ : std_logic;
signal \TXbufferZ0Z_5\ : std_logic;
signal \FTDI.TXshiftZ0Z_5\ : std_logic;
signal \INVFTDI.TXshift_4C_net\ : std_logic;
signal \ALU.b_10\ : std_logic;
signal \ALU.a_10\ : std_logic;
signal \ALU.r0_12_prm_7_10_s0_c_RNOZ0\ : std_logic;
signal \paramsZ0Z_3\ : std_logic;
signal \paramsZ0Z_2\ : std_logic;
signal \ALU.r4_RNII2A0LZ0Z_1\ : std_logic;
signal \ALU.lshift_3\ : std_logic;
signal \ALU.lshift63Z0Z_2\ : std_logic;
signal \ALU.r5_RNIAG9A9Z0Z_15\ : std_logic;
signal \ALU.r0_12_prm_8_14_s1_c_RNOZ0Z_1\ : std_logic;
signal op_i_0 : std_logic;
signal \ALU.un2_addsub_cry_0_c_RNIJPSHDZ0\ : std_logic;
signal \ALU.r0_12_prm_2_1_c_RNOZ0\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal op_1_cry_1 : std_logic;
signal op_1_cry_2 : std_logic;
signal op_1_cry_3 : std_logic;
signal \CLK_c_g\ : std_logic;
signal params5_g : std_logic;
signal \FTDI.N_208_0_cascade_\ : std_logic;
signal \FTDI.N_185_0_cascade_\ : std_logic;
signal \FTDI.N_207_0\ : std_logic;
signal \INVFTDI.TXstate_1C_net\ : std_logic;
signal \opZ0Z_0\ : std_logic;
signal \opZ0Z_3\ : std_logic;
signal \opZ0Z_1\ : std_logic;
signal \ALU.un1_op_1Z0Z_1_cascade_\ : std_logic;
signal \opZ0Z_4\ : std_logic;
signal \ALU.un1_op_1_0\ : std_logic;
signal \paramsZ0Z_1\ : std_logic;
signal \paramsZ0Z_0\ : std_logic;
signal \opZ0Z_2\ : std_logic;
signal \ALU.a_9\ : std_logic;
signal \ALU.r0_12_prm_4_9_s1_c_RNOZ0\ : std_logic;
signal \FTDI.TXstate_cnst_0_0_2_cascade_\ : std_logic;
signal \INVFTDI.TXstate_2C_net\ : std_logic;
signal \TXstartZ0\ : std_logic;
signal \FTDI.TXshiftZ0Z_1\ : std_logic;
signal \TXbufferZ0Z_0\ : std_logic;
signal \INVFTDI.TXshift_0C_net\ : std_logic;
signal \FTDI.un1_TXstate_0_sqmuxa_0_i\ : std_logic;
signal \bfn_18_6_0_\ : std_logic;
signal \FTDI.un3_TX_axb_3\ : std_logic;
signal \FTDI.un3_TX_cry_2\ : std_logic;
signal \FTDI.TXshiftZ0Z_0\ : std_logic;
signal \FTDI.un3_TX_cry_3\ : std_logic;
signal \FTDI_TX_0_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \FTDI.un3_TX_0_i\ : std_logic;
signal \FTDI.N_185_0\ : std_logic;
signal \INVFTDI.TXstate_0C_net\ : std_logic;
signal \FTDI.TXstateZ1Z_1\ : std_logic;
signal \FTDI.N_186_0\ : std_logic;
signal \FTDI.TXstate_e_1_3\ : std_logic;
signal \FTDI.N_186_0_cascade_\ : std_logic;
signal \FTDI.un3_TX_0\ : std_logic;
signal \INVFTDI.TXstate_3C_net\ : std_logic;
signal \FTDI.TXstateZ1Z_0\ : std_logic;
signal \FTDI.TXstateZ0Z_3\ : std_logic;
signal \FTDI.baudAccZ0Z_2\ : std_logic;
signal \FTDI.TXstate_e_1_0\ : std_logic;
signal \FTDI.TXready\ : std_logic;
signal \FTDI.baudAccZ0Z_0\ : std_logic;
signal \FTDI.baudAccZ0Z_1\ : std_logic;
signal \INVFTDI.baudAcc_0C_net\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \GPIO3_wire\ : std_logic;
signal \GPIO11_wire\ : std_logic;
signal \GPIO9_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    TX <= \TX_wire\;
    GPIO3 <= \GPIO3_wire\;
    GPIO11 <= \GPIO11_wire\;
    GPIO9 <= \GPIO9_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__57005\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57007\,
            DIN => \N__57006\,
            DOUT => \N__57005\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__57007\,
            PADOUT => \N__57006\,
            PADIN => \N__57005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TX_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56996\,
            DIN => \N__56995\,
            DOUT => \N__56994\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__56996\,
            PADOUT => \N__56995\,
            PADIN => \N__56994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__56524\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56987\,
            DIN => \N__56986\,
            DOUT => \N__56985\,
            PACKAGEPIN => \GPIO3_wire\
        );

    \GPIO3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__56987\,
            PADOUT => \N__56986\,
            PADIN => \N__56985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO11_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56978\,
            DIN => \N__56977\,
            DOUT => \N__56976\,
            PACKAGEPIN => \GPIO11_wire\
        );

    \GPIO11_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__56978\,
            PADOUT => \N__56977\,
            PADIN => \N__56976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO9_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56969\,
            DIN => \N__56968\,
            DOUT => \N__56967\,
            PACKAGEPIN => \GPIO9_wire\
        );

    \GPIO9_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__56969\,
            PADOUT => \N__56968\,
            PADIN => \N__56967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__56397\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__14264\ : InMux
    port map (
            O => \N__56950\,
            I => \N__56942\
        );

    \I__14263\ : InMux
    port map (
            O => \N__56949\,
            I => \N__56937\
        );

    \I__14262\ : InMux
    port map (
            O => \N__56948\,
            I => \N__56937\
        );

    \I__14261\ : InMux
    port map (
            O => \N__56947\,
            I => \N__56932\
        );

    \I__14260\ : InMux
    port map (
            O => \N__56946\,
            I => \N__56932\
        );

    \I__14259\ : InMux
    port map (
            O => \N__56945\,
            I => \N__56929\
        );

    \I__14258\ : LocalMux
    port map (
            O => \N__56942\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__14257\ : LocalMux
    port map (
            O => \N__56937\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__14256\ : LocalMux
    port map (
            O => \N__56932\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__14255\ : LocalMux
    port map (
            O => \N__56929\,
            I => \FTDI.TXstateZ1Z_1\
        );

    \I__14254\ : InMux
    port map (
            O => \N__56920\,
            I => \N__56917\
        );

    \I__14253\ : LocalMux
    port map (
            O => \N__56917\,
            I => \FTDI.N_186_0\
        );

    \I__14252\ : InMux
    port map (
            O => \N__56914\,
            I => \N__56911\
        );

    \I__14251\ : LocalMux
    port map (
            O => \N__56911\,
            I => \FTDI.TXstate_e_1_3\
        );

    \I__14250\ : CascadeMux
    port map (
            O => \N__56908\,
            I => \FTDI.N_186_0_cascade_\
        );

    \I__14249\ : InMux
    port map (
            O => \N__56905\,
            I => \N__56901\
        );

    \I__14248\ : CascadeMux
    port map (
            O => \N__56904\,
            I => \N__56897\
        );

    \I__14247\ : LocalMux
    port map (
            O => \N__56901\,
            I => \N__56891\
        );

    \I__14246\ : InMux
    port map (
            O => \N__56900\,
            I => \N__56888\
        );

    \I__14245\ : InMux
    port map (
            O => \N__56897\,
            I => \N__56885\
        );

    \I__14244\ : InMux
    port map (
            O => \N__56896\,
            I => \N__56882\
        );

    \I__14243\ : InMux
    port map (
            O => \N__56895\,
            I => \N__56877\
        );

    \I__14242\ : InMux
    port map (
            O => \N__56894\,
            I => \N__56877\
        );

    \I__14241\ : Odrv4
    port map (
            O => \N__56891\,
            I => \FTDI.un3_TX_0\
        );

    \I__14240\ : LocalMux
    port map (
            O => \N__56888\,
            I => \FTDI.un3_TX_0\
        );

    \I__14239\ : LocalMux
    port map (
            O => \N__56885\,
            I => \FTDI.un3_TX_0\
        );

    \I__14238\ : LocalMux
    port map (
            O => \N__56882\,
            I => \FTDI.un3_TX_0\
        );

    \I__14237\ : LocalMux
    port map (
            O => \N__56877\,
            I => \FTDI.un3_TX_0\
        );

    \I__14236\ : InMux
    port map (
            O => \N__56866\,
            I => \N__56858\
        );

    \I__14235\ : InMux
    port map (
            O => \N__56865\,
            I => \N__56851\
        );

    \I__14234\ : InMux
    port map (
            O => \N__56864\,
            I => \N__56851\
        );

    \I__14233\ : InMux
    port map (
            O => \N__56863\,
            I => \N__56851\
        );

    \I__14232\ : InMux
    port map (
            O => \N__56862\,
            I => \N__56846\
        );

    \I__14231\ : InMux
    port map (
            O => \N__56861\,
            I => \N__56846\
        );

    \I__14230\ : LocalMux
    port map (
            O => \N__56858\,
            I => \FTDI.TXstateZ1Z_0\
        );

    \I__14229\ : LocalMux
    port map (
            O => \N__56851\,
            I => \FTDI.TXstateZ1Z_0\
        );

    \I__14228\ : LocalMux
    port map (
            O => \N__56846\,
            I => \FTDI.TXstateZ1Z_0\
        );

    \I__14227\ : InMux
    port map (
            O => \N__56839\,
            I => \N__56826\
        );

    \I__14226\ : InMux
    port map (
            O => \N__56838\,
            I => \N__56826\
        );

    \I__14225\ : InMux
    port map (
            O => \N__56837\,
            I => \N__56817\
        );

    \I__14224\ : InMux
    port map (
            O => \N__56836\,
            I => \N__56817\
        );

    \I__14223\ : InMux
    port map (
            O => \N__56835\,
            I => \N__56817\
        );

    \I__14222\ : InMux
    port map (
            O => \N__56834\,
            I => \N__56817\
        );

    \I__14221\ : InMux
    port map (
            O => \N__56833\,
            I => \N__56811\
        );

    \I__14220\ : InMux
    port map (
            O => \N__56832\,
            I => \N__56811\
        );

    \I__14219\ : InMux
    port map (
            O => \N__56831\,
            I => \N__56807\
        );

    \I__14218\ : LocalMux
    port map (
            O => \N__56826\,
            I => \N__56804\
        );

    \I__14217\ : LocalMux
    port map (
            O => \N__56817\,
            I => \N__56801\
        );

    \I__14216\ : CascadeMux
    port map (
            O => \N__56816\,
            I => \N__56792\
        );

    \I__14215\ : LocalMux
    port map (
            O => \N__56811\,
            I => \N__56789\
        );

    \I__14214\ : InMux
    port map (
            O => \N__56810\,
            I => \N__56786\
        );

    \I__14213\ : LocalMux
    port map (
            O => \N__56807\,
            I => \N__56781\
        );

    \I__14212\ : Span4Mux_v
    port map (
            O => \N__56804\,
            I => \N__56781\
        );

    \I__14211\ : Span4Mux_h
    port map (
            O => \N__56801\,
            I => \N__56778\
        );

    \I__14210\ : InMux
    port map (
            O => \N__56800\,
            I => \N__56773\
        );

    \I__14209\ : InMux
    port map (
            O => \N__56799\,
            I => \N__56773\
        );

    \I__14208\ : InMux
    port map (
            O => \N__56798\,
            I => \N__56768\
        );

    \I__14207\ : InMux
    port map (
            O => \N__56797\,
            I => \N__56768\
        );

    \I__14206\ : InMux
    port map (
            O => \N__56796\,
            I => \N__56763\
        );

    \I__14205\ : InMux
    port map (
            O => \N__56795\,
            I => \N__56763\
        );

    \I__14204\ : InMux
    port map (
            O => \N__56792\,
            I => \N__56760\
        );

    \I__14203\ : Odrv4
    port map (
            O => \N__56789\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14202\ : LocalMux
    port map (
            O => \N__56786\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14201\ : Odrv4
    port map (
            O => \N__56781\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14200\ : Odrv4
    port map (
            O => \N__56778\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14199\ : LocalMux
    port map (
            O => \N__56773\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14198\ : LocalMux
    port map (
            O => \N__56768\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14197\ : LocalMux
    port map (
            O => \N__56763\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14196\ : LocalMux
    port map (
            O => \N__56760\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__14195\ : InMux
    port map (
            O => \N__56743\,
            I => \N__56732\
        );

    \I__14194\ : InMux
    port map (
            O => \N__56742\,
            I => \N__56732\
        );

    \I__14193\ : InMux
    port map (
            O => \N__56741\,
            I => \N__56727\
        );

    \I__14192\ : InMux
    port map (
            O => \N__56740\,
            I => \N__56727\
        );

    \I__14191\ : InMux
    port map (
            O => \N__56739\,
            I => \N__56720\
        );

    \I__14190\ : InMux
    port map (
            O => \N__56738\,
            I => \N__56720\
        );

    \I__14189\ : InMux
    port map (
            O => \N__56737\,
            I => \N__56720\
        );

    \I__14188\ : LocalMux
    port map (
            O => \N__56732\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__56727\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__14186\ : LocalMux
    port map (
            O => \N__56720\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__14185\ : CascadeMux
    port map (
            O => \N__56713\,
            I => \N__56710\
        );

    \I__14184\ : InMux
    port map (
            O => \N__56710\,
            I => \N__56707\
        );

    \I__14183\ : LocalMux
    port map (
            O => \N__56707\,
            I => \FTDI.TXstate_e_1_0\
        );

    \I__14182\ : InMux
    port map (
            O => \N__56704\,
            I => \N__56696\
        );

    \I__14181\ : InMux
    port map (
            O => \N__56703\,
            I => \N__56696\
        );

    \I__14180\ : CascadeMux
    port map (
            O => \N__56702\,
            I => \N__56692\
        );

    \I__14179\ : InMux
    port map (
            O => \N__56701\,
            I => \N__56689\
        );

    \I__14178\ : LocalMux
    port map (
            O => \N__56696\,
            I => \N__56686\
        );

    \I__14177\ : InMux
    port map (
            O => \N__56695\,
            I => \N__56681\
        );

    \I__14176\ : InMux
    port map (
            O => \N__56692\,
            I => \N__56681\
        );

    \I__14175\ : LocalMux
    port map (
            O => \N__56689\,
            I => \FTDI.TXready\
        );

    \I__14174\ : Odrv4
    port map (
            O => \N__56686\,
            I => \FTDI.TXready\
        );

    \I__14173\ : LocalMux
    port map (
            O => \N__56681\,
            I => \FTDI.TXready\
        );

    \I__14172\ : CascadeMux
    port map (
            O => \N__56674\,
            I => \N__56670\
        );

    \I__14171\ : InMux
    port map (
            O => \N__56673\,
            I => \N__56666\
        );

    \I__14170\ : InMux
    port map (
            O => \N__56670\,
            I => \N__56661\
        );

    \I__14169\ : InMux
    port map (
            O => \N__56669\,
            I => \N__56661\
        );

    \I__14168\ : LocalMux
    port map (
            O => \N__56666\,
            I => \FTDI.baudAccZ0Z_0\
        );

    \I__14167\ : LocalMux
    port map (
            O => \N__56661\,
            I => \FTDI.baudAccZ0Z_0\
        );

    \I__14166\ : InMux
    port map (
            O => \N__56656\,
            I => \N__56652\
        );

    \I__14165\ : InMux
    port map (
            O => \N__56655\,
            I => \N__56649\
        );

    \I__14164\ : LocalMux
    port map (
            O => \N__56652\,
            I => \FTDI.baudAccZ0Z_1\
        );

    \I__14163\ : LocalMux
    port map (
            O => \N__56649\,
            I => \FTDI.baudAccZ0Z_1\
        );

    \I__14162\ : CascadeMux
    port map (
            O => \N__56644\,
            I => \FTDI.TXstate_cnst_0_0_2_cascade_\
        );

    \I__14161\ : InMux
    port map (
            O => \N__56641\,
            I => \N__56635\
        );

    \I__14160\ : InMux
    port map (
            O => \N__56640\,
            I => \N__56635\
        );

    \I__14159\ : LocalMux
    port map (
            O => \N__56635\,
            I => \N__56632\
        );

    \I__14158\ : Span4Mux_v
    port map (
            O => \N__56632\,
            I => \N__56629\
        );

    \I__14157\ : Span4Mux_v
    port map (
            O => \N__56629\,
            I => \N__56626\
        );

    \I__14156\ : Sp12to4
    port map (
            O => \N__56626\,
            I => \N__56623\
        );

    \I__14155\ : Span12Mux_h
    port map (
            O => \N__56623\,
            I => \N__56620\
        );

    \I__14154\ : Odrv12
    port map (
            O => \N__56620\,
            I => \TXstartZ0\
        );

    \I__14153\ : InMux
    port map (
            O => \N__56617\,
            I => \N__56614\
        );

    \I__14152\ : LocalMux
    port map (
            O => \N__56614\,
            I => \FTDI.TXshiftZ0Z_1\
        );

    \I__14151\ : InMux
    port map (
            O => \N__56611\,
            I => \N__56608\
        );

    \I__14150\ : LocalMux
    port map (
            O => \N__56608\,
            I => \N__56605\
        );

    \I__14149\ : Span4Mux_v
    port map (
            O => \N__56605\,
            I => \N__56602\
        );

    \I__14148\ : Sp12to4
    port map (
            O => \N__56602\,
            I => \N__56599\
        );

    \I__14147\ : Span12Mux_h
    port map (
            O => \N__56599\,
            I => \N__56596\
        );

    \I__14146\ : Odrv12
    port map (
            O => \N__56596\,
            I => \TXbufferZ0Z_0\
        );

    \I__14145\ : CEMux
    port map (
            O => \N__56593\,
            I => \N__56590\
        );

    \I__14144\ : LocalMux
    port map (
            O => \N__56590\,
            I => \N__56587\
        );

    \I__14143\ : Span4Mux_v
    port map (
            O => \N__56587\,
            I => \N__56583\
        );

    \I__14142\ : CEMux
    port map (
            O => \N__56586\,
            I => \N__56580\
        );

    \I__14141\ : Span4Mux_v
    port map (
            O => \N__56583\,
            I => \N__56573\
        );

    \I__14140\ : LocalMux
    port map (
            O => \N__56580\,
            I => \N__56573\
        );

    \I__14139\ : CEMux
    port map (
            O => \N__56579\,
            I => \N__56570\
        );

    \I__14138\ : CEMux
    port map (
            O => \N__56578\,
            I => \N__56567\
        );

    \I__14137\ : Span4Mux_v
    port map (
            O => \N__56573\,
            I => \N__56564\
        );

    \I__14136\ : LocalMux
    port map (
            O => \N__56570\,
            I => \N__56561\
        );

    \I__14135\ : LocalMux
    port map (
            O => \N__56567\,
            I => \N__56558\
        );

    \I__14134\ : Span4Mux_v
    port map (
            O => \N__56564\,
            I => \N__56555\
        );

    \I__14133\ : Span4Mux_v
    port map (
            O => \N__56561\,
            I => \N__56550\
        );

    \I__14132\ : Span4Mux_h
    port map (
            O => \N__56558\,
            I => \N__56550\
        );

    \I__14131\ : Odrv4
    port map (
            O => \N__56555\,
            I => \FTDI.un1_TXstate_0_sqmuxa_0_i\
        );

    \I__14130\ : Odrv4
    port map (
            O => \N__56550\,
            I => \FTDI.un1_TXstate_0_sqmuxa_0_i\
        );

    \I__14129\ : InMux
    port map (
            O => \N__56545\,
            I => \N__56542\
        );

    \I__14128\ : LocalMux
    port map (
            O => \N__56542\,
            I => \FTDI.un3_TX_axb_3\
        );

    \I__14127\ : InMux
    port map (
            O => \N__56539\,
            I => \N__56536\
        );

    \I__14126\ : LocalMux
    port map (
            O => \N__56536\,
            I => \N__56533\
        );

    \I__14125\ : Span4Mux_v
    port map (
            O => \N__56533\,
            I => \N__56530\
        );

    \I__14124\ : Odrv4
    port map (
            O => \N__56530\,
            I => \FTDI.TXshiftZ0Z_0\
        );

    \I__14123\ : InMux
    port map (
            O => \N__56527\,
            I => \FTDI.un3_TX_cry_3\
        );

    \I__14122\ : IoInMux
    port map (
            O => \N__56524\,
            I => \N__56521\
        );

    \I__14121\ : LocalMux
    port map (
            O => \N__56521\,
            I => \N__56518\
        );

    \I__14120\ : Span12Mux_s5_v
    port map (
            O => \N__56518\,
            I => \N__56515\
        );

    \I__14119\ : Odrv12
    port map (
            O => \N__56515\,
            I => \FTDI_TX_0_i\
        );

    \I__14118\ : CascadeMux
    port map (
            O => \N__56512\,
            I => \N__56509\
        );

    \I__14117\ : InMux
    port map (
            O => \N__56509\,
            I => \N__56501\
        );

    \I__14116\ : CascadeMux
    port map (
            O => \N__56508\,
            I => \N__56498\
        );

    \I__14115\ : CascadeMux
    port map (
            O => \N__56507\,
            I => \N__56495\
        );

    \I__14114\ : CascadeMux
    port map (
            O => \N__56506\,
            I => \N__56492\
        );

    \I__14113\ : InMux
    port map (
            O => \N__56505\,
            I => \N__56489\
        );

    \I__14112\ : CascadeMux
    port map (
            O => \N__56504\,
            I => \N__56485\
        );

    \I__14111\ : LocalMux
    port map (
            O => \N__56501\,
            I => \N__56482\
        );

    \I__14110\ : InMux
    port map (
            O => \N__56498\,
            I => \N__56478\
        );

    \I__14109\ : InMux
    port map (
            O => \N__56495\,
            I => \N__56472\
        );

    \I__14108\ : InMux
    port map (
            O => \N__56492\,
            I => \N__56469\
        );

    \I__14107\ : LocalMux
    port map (
            O => \N__56489\,
            I => \N__56466\
        );

    \I__14106\ : InMux
    port map (
            O => \N__56488\,
            I => \N__56463\
        );

    \I__14105\ : InMux
    port map (
            O => \N__56485\,
            I => \N__56460\
        );

    \I__14104\ : Span4Mux_s1_v
    port map (
            O => \N__56482\,
            I => \N__56457\
        );

    \I__14103\ : CascadeMux
    port map (
            O => \N__56481\,
            I => \N__56454\
        );

    \I__14102\ : LocalMux
    port map (
            O => \N__56478\,
            I => \N__56451\
        );

    \I__14101\ : CascadeMux
    port map (
            O => \N__56477\,
            I => \N__56448\
        );

    \I__14100\ : CascadeMux
    port map (
            O => \N__56476\,
            I => \N__56445\
        );

    \I__14099\ : CascadeMux
    port map (
            O => \N__56475\,
            I => \N__56442\
        );

    \I__14098\ : LocalMux
    port map (
            O => \N__56472\,
            I => \N__56437\
        );

    \I__14097\ : LocalMux
    port map (
            O => \N__56469\,
            I => \N__56437\
        );

    \I__14096\ : Span4Mux_v
    port map (
            O => \N__56466\,
            I => \N__56434\
        );

    \I__14095\ : LocalMux
    port map (
            O => \N__56463\,
            I => \N__56431\
        );

    \I__14094\ : LocalMux
    port map (
            O => \N__56460\,
            I => \N__56426\
        );

    \I__14093\ : Span4Mux_h
    port map (
            O => \N__56457\,
            I => \N__56426\
        );

    \I__14092\ : InMux
    port map (
            O => \N__56454\,
            I => \N__56423\
        );

    \I__14091\ : Span4Mux_v
    port map (
            O => \N__56451\,
            I => \N__56420\
        );

    \I__14090\ : InMux
    port map (
            O => \N__56448\,
            I => \N__56417\
        );

    \I__14089\ : InMux
    port map (
            O => \N__56445\,
            I => \N__56414\
        );

    \I__14088\ : InMux
    port map (
            O => \N__56442\,
            I => \N__56410\
        );

    \I__14087\ : Span4Mux_v
    port map (
            O => \N__56437\,
            I => \N__56399\
        );

    \I__14086\ : Span4Mux_h
    port map (
            O => \N__56434\,
            I => \N__56399\
        );

    \I__14085\ : Span4Mux_v
    port map (
            O => \N__56431\,
            I => \N__56399\
        );

    \I__14084\ : Span4Mux_v
    port map (
            O => \N__56426\,
            I => \N__56399\
        );

    \I__14083\ : LocalMux
    port map (
            O => \N__56423\,
            I => \N__56399\
        );

    \I__14082\ : Span4Mux_v
    port map (
            O => \N__56420\,
            I => \N__56394\
        );

    \I__14081\ : LocalMux
    port map (
            O => \N__56417\,
            I => \N__56389\
        );

    \I__14080\ : LocalMux
    port map (
            O => \N__56414\,
            I => \N__56389\
        );

    \I__14079\ : CascadeMux
    port map (
            O => \N__56413\,
            I => \N__56386\
        );

    \I__14078\ : LocalMux
    port map (
            O => \N__56410\,
            I => \N__56381\
        );

    \I__14077\ : Span4Mux_v
    port map (
            O => \N__56399\,
            I => \N__56381\
        );

    \I__14076\ : InMux
    port map (
            O => \N__56398\,
            I => \N__56378\
        );

    \I__14075\ : IoInMux
    port map (
            O => \N__56397\,
            I => \N__56375\
        );

    \I__14074\ : Span4Mux_v
    port map (
            O => \N__56394\,
            I => \N__56372\
        );

    \I__14073\ : Span4Mux_v
    port map (
            O => \N__56389\,
            I => \N__56369\
        );

    \I__14072\ : InMux
    port map (
            O => \N__56386\,
            I => \N__56366\
        );

    \I__14071\ : Span4Mux_h
    port map (
            O => \N__56381\,
            I => \N__56363\
        );

    \I__14070\ : LocalMux
    port map (
            O => \N__56378\,
            I => \N__56360\
        );

    \I__14069\ : LocalMux
    port map (
            O => \N__56375\,
            I => \N__56357\
        );

    \I__14068\ : Sp12to4
    port map (
            O => \N__56372\,
            I => \N__56354\
        );

    \I__14067\ : Span4Mux_h
    port map (
            O => \N__56369\,
            I => \N__56351\
        );

    \I__14066\ : LocalMux
    port map (
            O => \N__56366\,
            I => \N__56348\
        );

    \I__14065\ : Span4Mux_h
    port map (
            O => \N__56363\,
            I => \N__56343\
        );

    \I__14064\ : Span4Mux_v
    port map (
            O => \N__56360\,
            I => \N__56343\
        );

    \I__14063\ : Span12Mux_s10_v
    port map (
            O => \N__56357\,
            I => \N__56334\
        );

    \I__14062\ : Span12Mux_h
    port map (
            O => \N__56354\,
            I => \N__56334\
        );

    \I__14061\ : Sp12to4
    port map (
            O => \N__56351\,
            I => \N__56334\
        );

    \I__14060\ : Sp12to4
    port map (
            O => \N__56348\,
            I => \N__56334\
        );

    \I__14059\ : Sp12to4
    port map (
            O => \N__56343\,
            I => \N__56331\
        );

    \I__14058\ : Span12Mux_v
    port map (
            O => \N__56334\,
            I => \N__56326\
        );

    \I__14057\ : Span12Mux_s5_h
    port map (
            O => \N__56331\,
            I => \N__56326\
        );

    \I__14056\ : Odrv12
    port map (
            O => \N__56326\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14055\ : InMux
    port map (
            O => \N__56323\,
            I => \N__56319\
        );

    \I__14054\ : InMux
    port map (
            O => \N__56322\,
            I => \N__56316\
        );

    \I__14053\ : LocalMux
    port map (
            O => \N__56319\,
            I => \FTDI.un3_TX_0_i\
        );

    \I__14052\ : LocalMux
    port map (
            O => \N__56316\,
            I => \FTDI.un3_TX_0_i\
        );

    \I__14051\ : InMux
    port map (
            O => \N__56311\,
            I => \N__56308\
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__56308\,
            I => \FTDI.N_185_0\
        );

    \I__14049\ : ClkMux
    port map (
            O => \N__56305\,
            I => \N__56065\
        );

    \I__14048\ : ClkMux
    port map (
            O => \N__56304\,
            I => \N__56065\
        );

    \I__14047\ : ClkMux
    port map (
            O => \N__56303\,
            I => \N__56065\
        );

    \I__14046\ : ClkMux
    port map (
            O => \N__56302\,
            I => \N__56065\
        );

    \I__14045\ : ClkMux
    port map (
            O => \N__56301\,
            I => \N__56065\
        );

    \I__14044\ : ClkMux
    port map (
            O => \N__56300\,
            I => \N__56065\
        );

    \I__14043\ : ClkMux
    port map (
            O => \N__56299\,
            I => \N__56065\
        );

    \I__14042\ : ClkMux
    port map (
            O => \N__56298\,
            I => \N__56065\
        );

    \I__14041\ : ClkMux
    port map (
            O => \N__56297\,
            I => \N__56065\
        );

    \I__14040\ : ClkMux
    port map (
            O => \N__56296\,
            I => \N__56065\
        );

    \I__14039\ : ClkMux
    port map (
            O => \N__56295\,
            I => \N__56065\
        );

    \I__14038\ : ClkMux
    port map (
            O => \N__56294\,
            I => \N__56065\
        );

    \I__14037\ : ClkMux
    port map (
            O => \N__56293\,
            I => \N__56065\
        );

    \I__14036\ : ClkMux
    port map (
            O => \N__56292\,
            I => \N__56065\
        );

    \I__14035\ : ClkMux
    port map (
            O => \N__56291\,
            I => \N__56065\
        );

    \I__14034\ : ClkMux
    port map (
            O => \N__56290\,
            I => \N__56065\
        );

    \I__14033\ : ClkMux
    port map (
            O => \N__56289\,
            I => \N__56065\
        );

    \I__14032\ : ClkMux
    port map (
            O => \N__56288\,
            I => \N__56065\
        );

    \I__14031\ : ClkMux
    port map (
            O => \N__56287\,
            I => \N__56065\
        );

    \I__14030\ : ClkMux
    port map (
            O => \N__56286\,
            I => \N__56065\
        );

    \I__14029\ : ClkMux
    port map (
            O => \N__56285\,
            I => \N__56065\
        );

    \I__14028\ : ClkMux
    port map (
            O => \N__56284\,
            I => \N__56065\
        );

    \I__14027\ : ClkMux
    port map (
            O => \N__56283\,
            I => \N__56065\
        );

    \I__14026\ : ClkMux
    port map (
            O => \N__56282\,
            I => \N__56065\
        );

    \I__14025\ : ClkMux
    port map (
            O => \N__56281\,
            I => \N__56065\
        );

    \I__14024\ : ClkMux
    port map (
            O => \N__56280\,
            I => \N__56065\
        );

    \I__14023\ : ClkMux
    port map (
            O => \N__56279\,
            I => \N__56065\
        );

    \I__14022\ : ClkMux
    port map (
            O => \N__56278\,
            I => \N__56065\
        );

    \I__14021\ : ClkMux
    port map (
            O => \N__56277\,
            I => \N__56065\
        );

    \I__14020\ : ClkMux
    port map (
            O => \N__56276\,
            I => \N__56065\
        );

    \I__14019\ : ClkMux
    port map (
            O => \N__56275\,
            I => \N__56065\
        );

    \I__14018\ : ClkMux
    port map (
            O => \N__56274\,
            I => \N__56065\
        );

    \I__14017\ : ClkMux
    port map (
            O => \N__56273\,
            I => \N__56065\
        );

    \I__14016\ : ClkMux
    port map (
            O => \N__56272\,
            I => \N__56065\
        );

    \I__14015\ : ClkMux
    port map (
            O => \N__56271\,
            I => \N__56065\
        );

    \I__14014\ : ClkMux
    port map (
            O => \N__56270\,
            I => \N__56065\
        );

    \I__14013\ : ClkMux
    port map (
            O => \N__56269\,
            I => \N__56065\
        );

    \I__14012\ : ClkMux
    port map (
            O => \N__56268\,
            I => \N__56065\
        );

    \I__14011\ : ClkMux
    port map (
            O => \N__56267\,
            I => \N__56065\
        );

    \I__14010\ : ClkMux
    port map (
            O => \N__56266\,
            I => \N__56065\
        );

    \I__14009\ : ClkMux
    port map (
            O => \N__56265\,
            I => \N__56065\
        );

    \I__14008\ : ClkMux
    port map (
            O => \N__56264\,
            I => \N__56065\
        );

    \I__14007\ : ClkMux
    port map (
            O => \N__56263\,
            I => \N__56065\
        );

    \I__14006\ : ClkMux
    port map (
            O => \N__56262\,
            I => \N__56065\
        );

    \I__14005\ : ClkMux
    port map (
            O => \N__56261\,
            I => \N__56065\
        );

    \I__14004\ : ClkMux
    port map (
            O => \N__56260\,
            I => \N__56065\
        );

    \I__14003\ : ClkMux
    port map (
            O => \N__56259\,
            I => \N__56065\
        );

    \I__14002\ : ClkMux
    port map (
            O => \N__56258\,
            I => \N__56065\
        );

    \I__14001\ : ClkMux
    port map (
            O => \N__56257\,
            I => \N__56065\
        );

    \I__14000\ : ClkMux
    port map (
            O => \N__56256\,
            I => \N__56065\
        );

    \I__13999\ : ClkMux
    port map (
            O => \N__56255\,
            I => \N__56065\
        );

    \I__13998\ : ClkMux
    port map (
            O => \N__56254\,
            I => \N__56065\
        );

    \I__13997\ : ClkMux
    port map (
            O => \N__56253\,
            I => \N__56065\
        );

    \I__13996\ : ClkMux
    port map (
            O => \N__56252\,
            I => \N__56065\
        );

    \I__13995\ : ClkMux
    port map (
            O => \N__56251\,
            I => \N__56065\
        );

    \I__13994\ : ClkMux
    port map (
            O => \N__56250\,
            I => \N__56065\
        );

    \I__13993\ : ClkMux
    port map (
            O => \N__56249\,
            I => \N__56065\
        );

    \I__13992\ : ClkMux
    port map (
            O => \N__56248\,
            I => \N__56065\
        );

    \I__13991\ : ClkMux
    port map (
            O => \N__56247\,
            I => \N__56065\
        );

    \I__13990\ : ClkMux
    port map (
            O => \N__56246\,
            I => \N__56065\
        );

    \I__13989\ : ClkMux
    port map (
            O => \N__56245\,
            I => \N__56065\
        );

    \I__13988\ : ClkMux
    port map (
            O => \N__56244\,
            I => \N__56065\
        );

    \I__13987\ : ClkMux
    port map (
            O => \N__56243\,
            I => \N__56065\
        );

    \I__13986\ : ClkMux
    port map (
            O => \N__56242\,
            I => \N__56065\
        );

    \I__13985\ : ClkMux
    port map (
            O => \N__56241\,
            I => \N__56065\
        );

    \I__13984\ : ClkMux
    port map (
            O => \N__56240\,
            I => \N__56065\
        );

    \I__13983\ : ClkMux
    port map (
            O => \N__56239\,
            I => \N__56065\
        );

    \I__13982\ : ClkMux
    port map (
            O => \N__56238\,
            I => \N__56065\
        );

    \I__13981\ : ClkMux
    port map (
            O => \N__56237\,
            I => \N__56065\
        );

    \I__13980\ : ClkMux
    port map (
            O => \N__56236\,
            I => \N__56065\
        );

    \I__13979\ : ClkMux
    port map (
            O => \N__56235\,
            I => \N__56065\
        );

    \I__13978\ : ClkMux
    port map (
            O => \N__56234\,
            I => \N__56065\
        );

    \I__13977\ : ClkMux
    port map (
            O => \N__56233\,
            I => \N__56065\
        );

    \I__13976\ : ClkMux
    port map (
            O => \N__56232\,
            I => \N__56065\
        );

    \I__13975\ : ClkMux
    port map (
            O => \N__56231\,
            I => \N__56065\
        );

    \I__13974\ : ClkMux
    port map (
            O => \N__56230\,
            I => \N__56065\
        );

    \I__13973\ : ClkMux
    port map (
            O => \N__56229\,
            I => \N__56065\
        );

    \I__13972\ : ClkMux
    port map (
            O => \N__56228\,
            I => \N__56065\
        );

    \I__13971\ : ClkMux
    port map (
            O => \N__56227\,
            I => \N__56065\
        );

    \I__13970\ : ClkMux
    port map (
            O => \N__56226\,
            I => \N__56065\
        );

    \I__13969\ : GlobalMux
    port map (
            O => \N__56065\,
            I => \N__56062\
        );

    \I__13968\ : gio2CtrlBuf
    port map (
            O => \N__56062\,
            I => \CLK_c_g\
        );

    \I__13967\ : CEMux
    port map (
            O => \N__56059\,
            I => \N__55987\
        );

    \I__13966\ : CEMux
    port map (
            O => \N__56058\,
            I => \N__55987\
        );

    \I__13965\ : CEMux
    port map (
            O => \N__56057\,
            I => \N__55987\
        );

    \I__13964\ : CEMux
    port map (
            O => \N__56056\,
            I => \N__55987\
        );

    \I__13963\ : CEMux
    port map (
            O => \N__56055\,
            I => \N__55987\
        );

    \I__13962\ : CEMux
    port map (
            O => \N__56054\,
            I => \N__55987\
        );

    \I__13961\ : CEMux
    port map (
            O => \N__56053\,
            I => \N__55987\
        );

    \I__13960\ : CEMux
    port map (
            O => \N__56052\,
            I => \N__55987\
        );

    \I__13959\ : CEMux
    port map (
            O => \N__56051\,
            I => \N__55987\
        );

    \I__13958\ : CEMux
    port map (
            O => \N__56050\,
            I => \N__55987\
        );

    \I__13957\ : CEMux
    port map (
            O => \N__56049\,
            I => \N__55987\
        );

    \I__13956\ : CEMux
    port map (
            O => \N__56048\,
            I => \N__55987\
        );

    \I__13955\ : CEMux
    port map (
            O => \N__56047\,
            I => \N__55987\
        );

    \I__13954\ : CEMux
    port map (
            O => \N__56046\,
            I => \N__55987\
        );

    \I__13953\ : CEMux
    port map (
            O => \N__56045\,
            I => \N__55987\
        );

    \I__13952\ : CEMux
    port map (
            O => \N__56044\,
            I => \N__55987\
        );

    \I__13951\ : CEMux
    port map (
            O => \N__56043\,
            I => \N__55987\
        );

    \I__13950\ : CEMux
    port map (
            O => \N__56042\,
            I => \N__55987\
        );

    \I__13949\ : CEMux
    port map (
            O => \N__56041\,
            I => \N__55987\
        );

    \I__13948\ : CEMux
    port map (
            O => \N__56040\,
            I => \N__55987\
        );

    \I__13947\ : CEMux
    port map (
            O => \N__56039\,
            I => \N__55987\
        );

    \I__13946\ : CEMux
    port map (
            O => \N__56038\,
            I => \N__55987\
        );

    \I__13945\ : CEMux
    port map (
            O => \N__56037\,
            I => \N__55987\
        );

    \I__13944\ : CEMux
    port map (
            O => \N__56036\,
            I => \N__55987\
        );

    \I__13943\ : GlobalMux
    port map (
            O => \N__55987\,
            I => \N__55984\
        );

    \I__13942\ : gio2CtrlBuf
    port map (
            O => \N__55984\,
            I => params5_g
        );

    \I__13941\ : CascadeMux
    port map (
            O => \N__55981\,
            I => \FTDI.N_208_0_cascade_\
        );

    \I__13940\ : CascadeMux
    port map (
            O => \N__55978\,
            I => \FTDI.N_185_0_cascade_\
        );

    \I__13939\ : InMux
    port map (
            O => \N__55975\,
            I => \N__55972\
        );

    \I__13938\ : LocalMux
    port map (
            O => \N__55972\,
            I => \FTDI.N_207_0\
        );

    \I__13937\ : InMux
    port map (
            O => \N__55969\,
            I => \N__55965\
        );

    \I__13936\ : InMux
    port map (
            O => \N__55968\,
            I => \N__55962\
        );

    \I__13935\ : LocalMux
    port map (
            O => \N__55965\,
            I => \N__55952\
        );

    \I__13934\ : LocalMux
    port map (
            O => \N__55962\,
            I => \N__55947\
        );

    \I__13933\ : CascadeMux
    port map (
            O => \N__55961\,
            I => \N__55943\
        );

    \I__13932\ : InMux
    port map (
            O => \N__55960\,
            I => \N__55934\
        );

    \I__13931\ : InMux
    port map (
            O => \N__55959\,
            I => \N__55934\
        );

    \I__13930\ : InMux
    port map (
            O => \N__55958\,
            I => \N__55924\
        );

    \I__13929\ : InMux
    port map (
            O => \N__55957\,
            I => \N__55921\
        );

    \I__13928\ : CascadeMux
    port map (
            O => \N__55956\,
            I => \N__55916\
        );

    \I__13927\ : CascadeMux
    port map (
            O => \N__55955\,
            I => \N__55913\
        );

    \I__13926\ : Span4Mux_h
    port map (
            O => \N__55952\,
            I => \N__55910\
        );

    \I__13925\ : InMux
    port map (
            O => \N__55951\,
            I => \N__55905\
        );

    \I__13924\ : InMux
    port map (
            O => \N__55950\,
            I => \N__55905\
        );

    \I__13923\ : Span4Mux_h
    port map (
            O => \N__55947\,
            I => \N__55896\
        );

    \I__13922\ : InMux
    port map (
            O => \N__55946\,
            I => \N__55893\
        );

    \I__13921\ : InMux
    port map (
            O => \N__55943\,
            I => \N__55888\
        );

    \I__13920\ : InMux
    port map (
            O => \N__55942\,
            I => \N__55888\
        );

    \I__13919\ : InMux
    port map (
            O => \N__55941\,
            I => \N__55885\
        );

    \I__13918\ : InMux
    port map (
            O => \N__55940\,
            I => \N__55882\
        );

    \I__13917\ : InMux
    port map (
            O => \N__55939\,
            I => \N__55879\
        );

    \I__13916\ : LocalMux
    port map (
            O => \N__55934\,
            I => \N__55876\
        );

    \I__13915\ : InMux
    port map (
            O => \N__55933\,
            I => \N__55871\
        );

    \I__13914\ : InMux
    port map (
            O => \N__55932\,
            I => \N__55871\
        );

    \I__13913\ : InMux
    port map (
            O => \N__55931\,
            I => \N__55862\
        );

    \I__13912\ : InMux
    port map (
            O => \N__55930\,
            I => \N__55862\
        );

    \I__13911\ : InMux
    port map (
            O => \N__55929\,
            I => \N__55862\
        );

    \I__13910\ : InMux
    port map (
            O => \N__55928\,
            I => \N__55862\
        );

    \I__13909\ : InMux
    port map (
            O => \N__55927\,
            I => \N__55858\
        );

    \I__13908\ : LocalMux
    port map (
            O => \N__55924\,
            I => \N__55853\
        );

    \I__13907\ : LocalMux
    port map (
            O => \N__55921\,
            I => \N__55853\
        );

    \I__13906\ : InMux
    port map (
            O => \N__55920\,
            I => \N__55848\
        );

    \I__13905\ : InMux
    port map (
            O => \N__55919\,
            I => \N__55848\
        );

    \I__13904\ : InMux
    port map (
            O => \N__55916\,
            I => \N__55842\
        );

    \I__13903\ : InMux
    port map (
            O => \N__55913\,
            I => \N__55842\
        );

    \I__13902\ : Span4Mux_h
    port map (
            O => \N__55910\,
            I => \N__55834\
        );

    \I__13901\ : LocalMux
    port map (
            O => \N__55905\,
            I => \N__55834\
        );

    \I__13900\ : InMux
    port map (
            O => \N__55904\,
            I => \N__55831\
        );

    \I__13899\ : InMux
    port map (
            O => \N__55903\,
            I => \N__55826\
        );

    \I__13898\ : InMux
    port map (
            O => \N__55902\,
            I => \N__55826\
        );

    \I__13897\ : InMux
    port map (
            O => \N__55901\,
            I => \N__55819\
        );

    \I__13896\ : InMux
    port map (
            O => \N__55900\,
            I => \N__55819\
        );

    \I__13895\ : InMux
    port map (
            O => \N__55899\,
            I => \N__55819\
        );

    \I__13894\ : Span4Mux_h
    port map (
            O => \N__55896\,
            I => \N__55814\
        );

    \I__13893\ : LocalMux
    port map (
            O => \N__55893\,
            I => \N__55809\
        );

    \I__13892\ : LocalMux
    port map (
            O => \N__55888\,
            I => \N__55809\
        );

    \I__13891\ : LocalMux
    port map (
            O => \N__55885\,
            I => \N__55802\
        );

    \I__13890\ : LocalMux
    port map (
            O => \N__55882\,
            I => \N__55787\
        );

    \I__13889\ : LocalMux
    port map (
            O => \N__55879\,
            I => \N__55787\
        );

    \I__13888\ : Span4Mux_v
    port map (
            O => \N__55876\,
            I => \N__55787\
        );

    \I__13887\ : LocalMux
    port map (
            O => \N__55871\,
            I => \N__55787\
        );

    \I__13886\ : LocalMux
    port map (
            O => \N__55862\,
            I => \N__55787\
        );

    \I__13885\ : InMux
    port map (
            O => \N__55861\,
            I => \N__55784\
        );

    \I__13884\ : LocalMux
    port map (
            O => \N__55858\,
            I => \N__55777\
        );

    \I__13883\ : Span4Mux_v
    port map (
            O => \N__55853\,
            I => \N__55777\
        );

    \I__13882\ : LocalMux
    port map (
            O => \N__55848\,
            I => \N__55777\
        );

    \I__13881\ : CascadeMux
    port map (
            O => \N__55847\,
            I => \N__55773\
        );

    \I__13880\ : LocalMux
    port map (
            O => \N__55842\,
            I => \N__55769\
        );

    \I__13879\ : InMux
    port map (
            O => \N__55841\,
            I => \N__55766\
        );

    \I__13878\ : InMux
    port map (
            O => \N__55840\,
            I => \N__55763\
        );

    \I__13877\ : CascadeMux
    port map (
            O => \N__55839\,
            I => \N__55760\
        );

    \I__13876\ : Span4Mux_h
    port map (
            O => \N__55834\,
            I => \N__55754\
        );

    \I__13875\ : LocalMux
    port map (
            O => \N__55831\,
            I => \N__55754\
        );

    \I__13874\ : LocalMux
    port map (
            O => \N__55826\,
            I => \N__55749\
        );

    \I__13873\ : LocalMux
    port map (
            O => \N__55819\,
            I => \N__55749\
        );

    \I__13872\ : InMux
    port map (
            O => \N__55818\,
            I => \N__55744\
        );

    \I__13871\ : InMux
    port map (
            O => \N__55817\,
            I => \N__55744\
        );

    \I__13870\ : Span4Mux_v
    port map (
            O => \N__55814\,
            I => \N__55741\
        );

    \I__13869\ : Span4Mux_h
    port map (
            O => \N__55809\,
            I => \N__55738\
        );

    \I__13868\ : InMux
    port map (
            O => \N__55808\,
            I => \N__55731\
        );

    \I__13867\ : InMux
    port map (
            O => \N__55807\,
            I => \N__55731\
        );

    \I__13866\ : InMux
    port map (
            O => \N__55806\,
            I => \N__55724\
        );

    \I__13865\ : InMux
    port map (
            O => \N__55805\,
            I => \N__55724\
        );

    \I__13864\ : Span4Mux_h
    port map (
            O => \N__55802\,
            I => \N__55719\
        );

    \I__13863\ : InMux
    port map (
            O => \N__55801\,
            I => \N__55716\
        );

    \I__13862\ : InMux
    port map (
            O => \N__55800\,
            I => \N__55709\
        );

    \I__13861\ : InMux
    port map (
            O => \N__55799\,
            I => \N__55709\
        );

    \I__13860\ : InMux
    port map (
            O => \N__55798\,
            I => \N__55709\
        );

    \I__13859\ : Span4Mux_v
    port map (
            O => \N__55787\,
            I => \N__55706\
        );

    \I__13858\ : LocalMux
    port map (
            O => \N__55784\,
            I => \N__55701\
        );

    \I__13857\ : Span4Mux_v
    port map (
            O => \N__55777\,
            I => \N__55701\
        );

    \I__13856\ : InMux
    port map (
            O => \N__55776\,
            I => \N__55694\
        );

    \I__13855\ : InMux
    port map (
            O => \N__55773\,
            I => \N__55694\
        );

    \I__13854\ : InMux
    port map (
            O => \N__55772\,
            I => \N__55694\
        );

    \I__13853\ : Span4Mux_h
    port map (
            O => \N__55769\,
            I => \N__55690\
        );

    \I__13852\ : LocalMux
    port map (
            O => \N__55766\,
            I => \N__55685\
        );

    \I__13851\ : LocalMux
    port map (
            O => \N__55763\,
            I => \N__55685\
        );

    \I__13850\ : InMux
    port map (
            O => \N__55760\,
            I => \N__55682\
        );

    \I__13849\ : InMux
    port map (
            O => \N__55759\,
            I => \N__55679\
        );

    \I__13848\ : Span4Mux_h
    port map (
            O => \N__55754\,
            I => \N__55676\
        );

    \I__13847\ : Span4Mux_v
    port map (
            O => \N__55749\,
            I => \N__55671\
        );

    \I__13846\ : LocalMux
    port map (
            O => \N__55744\,
            I => \N__55671\
        );

    \I__13845\ : Span4Mux_h
    port map (
            O => \N__55741\,
            I => \N__55666\
        );

    \I__13844\ : Span4Mux_v
    port map (
            O => \N__55738\,
            I => \N__55666\
        );

    \I__13843\ : InMux
    port map (
            O => \N__55737\,
            I => \N__55663\
        );

    \I__13842\ : InMux
    port map (
            O => \N__55736\,
            I => \N__55660\
        );

    \I__13841\ : LocalMux
    port map (
            O => \N__55731\,
            I => \N__55656\
        );

    \I__13840\ : InMux
    port map (
            O => \N__55730\,
            I => \N__55653\
        );

    \I__13839\ : InMux
    port map (
            O => \N__55729\,
            I => \N__55650\
        );

    \I__13838\ : LocalMux
    port map (
            O => \N__55724\,
            I => \N__55647\
        );

    \I__13837\ : InMux
    port map (
            O => \N__55723\,
            I => \N__55642\
        );

    \I__13836\ : InMux
    port map (
            O => \N__55722\,
            I => \N__55642\
        );

    \I__13835\ : Span4Mux_h
    port map (
            O => \N__55719\,
            I => \N__55631\
        );

    \I__13834\ : LocalMux
    port map (
            O => \N__55716\,
            I => \N__55631\
        );

    \I__13833\ : LocalMux
    port map (
            O => \N__55709\,
            I => \N__55631\
        );

    \I__13832\ : Span4Mux_h
    port map (
            O => \N__55706\,
            I => \N__55631\
        );

    \I__13831\ : Sp12to4
    port map (
            O => \N__55701\,
            I => \N__55626\
        );

    \I__13830\ : LocalMux
    port map (
            O => \N__55694\,
            I => \N__55626\
        );

    \I__13829\ : InMux
    port map (
            O => \N__55693\,
            I => \N__55623\
        );

    \I__13828\ : Span4Mux_h
    port map (
            O => \N__55690\,
            I => \N__55618\
        );

    \I__13827\ : Span4Mux_h
    port map (
            O => \N__55685\,
            I => \N__55618\
        );

    \I__13826\ : LocalMux
    port map (
            O => \N__55682\,
            I => \N__55609\
        );

    \I__13825\ : LocalMux
    port map (
            O => \N__55679\,
            I => \N__55609\
        );

    \I__13824\ : Span4Mux_v
    port map (
            O => \N__55676\,
            I => \N__55609\
        );

    \I__13823\ : Span4Mux_h
    port map (
            O => \N__55671\,
            I => \N__55609\
        );

    \I__13822\ : Span4Mux_v
    port map (
            O => \N__55666\,
            I => \N__55604\
        );

    \I__13821\ : LocalMux
    port map (
            O => \N__55663\,
            I => \N__55604\
        );

    \I__13820\ : LocalMux
    port map (
            O => \N__55660\,
            I => \N__55601\
        );

    \I__13819\ : InMux
    port map (
            O => \N__55659\,
            I => \N__55598\
        );

    \I__13818\ : Span4Mux_h
    port map (
            O => \N__55656\,
            I => \N__55589\
        );

    \I__13817\ : LocalMux
    port map (
            O => \N__55653\,
            I => \N__55589\
        );

    \I__13816\ : LocalMux
    port map (
            O => \N__55650\,
            I => \N__55589\
        );

    \I__13815\ : Span4Mux_h
    port map (
            O => \N__55647\,
            I => \N__55589\
        );

    \I__13814\ : LocalMux
    port map (
            O => \N__55642\,
            I => \N__55586\
        );

    \I__13813\ : InMux
    port map (
            O => \N__55641\,
            I => \N__55582\
        );

    \I__13812\ : InMux
    port map (
            O => \N__55640\,
            I => \N__55579\
        );

    \I__13811\ : Sp12to4
    port map (
            O => \N__55631\,
            I => \N__55574\
        );

    \I__13810\ : Span12Mux_h
    port map (
            O => \N__55626\,
            I => \N__55574\
        );

    \I__13809\ : LocalMux
    port map (
            O => \N__55623\,
            I => \N__55567\
        );

    \I__13808\ : Span4Mux_h
    port map (
            O => \N__55618\,
            I => \N__55567\
        );

    \I__13807\ : Span4Mux_v
    port map (
            O => \N__55609\,
            I => \N__55567\
        );

    \I__13806\ : Span4Mux_h
    port map (
            O => \N__55604\,
            I => \N__55564\
        );

    \I__13805\ : Span4Mux_h
    port map (
            O => \N__55601\,
            I => \N__55555\
        );

    \I__13804\ : LocalMux
    port map (
            O => \N__55598\,
            I => \N__55555\
        );

    \I__13803\ : Span4Mux_v
    port map (
            O => \N__55589\,
            I => \N__55555\
        );

    \I__13802\ : Span4Mux_s2_v
    port map (
            O => \N__55586\,
            I => \N__55555\
        );

    \I__13801\ : InMux
    port map (
            O => \N__55585\,
            I => \N__55552\
        );

    \I__13800\ : LocalMux
    port map (
            O => \N__55582\,
            I => \opZ0Z_0\
        );

    \I__13799\ : LocalMux
    port map (
            O => \N__55579\,
            I => \opZ0Z_0\
        );

    \I__13798\ : Odrv12
    port map (
            O => \N__55574\,
            I => \opZ0Z_0\
        );

    \I__13797\ : Odrv4
    port map (
            O => \N__55567\,
            I => \opZ0Z_0\
        );

    \I__13796\ : Odrv4
    port map (
            O => \N__55564\,
            I => \opZ0Z_0\
        );

    \I__13795\ : Odrv4
    port map (
            O => \N__55555\,
            I => \opZ0Z_0\
        );

    \I__13794\ : LocalMux
    port map (
            O => \N__55552\,
            I => \opZ0Z_0\
        );

    \I__13793\ : CascadeMux
    port map (
            O => \N__55537\,
            I => \N__55530\
        );

    \I__13792\ : CascadeMux
    port map (
            O => \N__55536\,
            I => \N__55524\
        );

    \I__13791\ : InMux
    port map (
            O => \N__55535\,
            I => \N__55518\
        );

    \I__13790\ : CascadeMux
    port map (
            O => \N__55534\,
            I => \N__55514\
        );

    \I__13789\ : InMux
    port map (
            O => \N__55533\,
            I => \N__55510\
        );

    \I__13788\ : InMux
    port map (
            O => \N__55530\,
            I => \N__55507\
        );

    \I__13787\ : InMux
    port map (
            O => \N__55529\,
            I => \N__55503\
        );

    \I__13786\ : InMux
    port map (
            O => \N__55528\,
            I => \N__55500\
        );

    \I__13785\ : InMux
    port map (
            O => \N__55527\,
            I => \N__55497\
        );

    \I__13784\ : InMux
    port map (
            O => \N__55524\,
            I => \N__55492\
        );

    \I__13783\ : InMux
    port map (
            O => \N__55523\,
            I => \N__55492\
        );

    \I__13782\ : CascadeMux
    port map (
            O => \N__55522\,
            I => \N__55485\
        );

    \I__13781\ : InMux
    port map (
            O => \N__55521\,
            I => \N__55482\
        );

    \I__13780\ : LocalMux
    port map (
            O => \N__55518\,
            I => \N__55477\
        );

    \I__13779\ : InMux
    port map (
            O => \N__55517\,
            I => \N__55473\
        );

    \I__13778\ : InMux
    port map (
            O => \N__55514\,
            I => \N__55468\
        );

    \I__13777\ : InMux
    port map (
            O => \N__55513\,
            I => \N__55468\
        );

    \I__13776\ : LocalMux
    port map (
            O => \N__55510\,
            I => \N__55465\
        );

    \I__13775\ : LocalMux
    port map (
            O => \N__55507\,
            I => \N__55462\
        );

    \I__13774\ : InMux
    port map (
            O => \N__55506\,
            I => \N__55459\
        );

    \I__13773\ : LocalMux
    port map (
            O => \N__55503\,
            I => \N__55449\
        );

    \I__13772\ : LocalMux
    port map (
            O => \N__55500\,
            I => \N__55449\
        );

    \I__13771\ : LocalMux
    port map (
            O => \N__55497\,
            I => \N__55449\
        );

    \I__13770\ : LocalMux
    port map (
            O => \N__55492\,
            I => \N__55449\
        );

    \I__13769\ : InMux
    port map (
            O => \N__55491\,
            I => \N__55441\
        );

    \I__13768\ : InMux
    port map (
            O => \N__55490\,
            I => \N__55441\
        );

    \I__13767\ : InMux
    port map (
            O => \N__55489\,
            I => \N__55438\
        );

    \I__13766\ : InMux
    port map (
            O => \N__55488\,
            I => \N__55435\
        );

    \I__13765\ : InMux
    port map (
            O => \N__55485\,
            I => \N__55431\
        );

    \I__13764\ : LocalMux
    port map (
            O => \N__55482\,
            I => \N__55428\
        );

    \I__13763\ : InMux
    port map (
            O => \N__55481\,
            I => \N__55423\
        );

    \I__13762\ : InMux
    port map (
            O => \N__55480\,
            I => \N__55423\
        );

    \I__13761\ : Span4Mux_h
    port map (
            O => \N__55477\,
            I => \N__55420\
        );

    \I__13760\ : InMux
    port map (
            O => \N__55476\,
            I => \N__55417\
        );

    \I__13759\ : LocalMux
    port map (
            O => \N__55473\,
            I => \N__55414\
        );

    \I__13758\ : LocalMux
    port map (
            O => \N__55468\,
            I => \N__55411\
        );

    \I__13757\ : Span4Mux_v
    port map (
            O => \N__55465\,
            I => \N__55404\
        );

    \I__13756\ : Span4Mux_h
    port map (
            O => \N__55462\,
            I => \N__55404\
        );

    \I__13755\ : LocalMux
    port map (
            O => \N__55459\,
            I => \N__55404\
        );

    \I__13754\ : InMux
    port map (
            O => \N__55458\,
            I => \N__55401\
        );

    \I__13753\ : Span4Mux_v
    port map (
            O => \N__55449\,
            I => \N__55396\
        );

    \I__13752\ : InMux
    port map (
            O => \N__55448\,
            I => \N__55393\
        );

    \I__13751\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55388\
        );

    \I__13750\ : InMux
    port map (
            O => \N__55446\,
            I => \N__55388\
        );

    \I__13749\ : LocalMux
    port map (
            O => \N__55441\,
            I => \N__55383\
        );

    \I__13748\ : LocalMux
    port map (
            O => \N__55438\,
            I => \N__55383\
        );

    \I__13747\ : LocalMux
    port map (
            O => \N__55435\,
            I => \N__55378\
        );

    \I__13746\ : InMux
    port map (
            O => \N__55434\,
            I => \N__55375\
        );

    \I__13745\ : LocalMux
    port map (
            O => \N__55431\,
            I => \N__55366\
        );

    \I__13744\ : Span4Mux_h
    port map (
            O => \N__55428\,
            I => \N__55366\
        );

    \I__13743\ : LocalMux
    port map (
            O => \N__55423\,
            I => \N__55366\
        );

    \I__13742\ : Span4Mux_v
    port map (
            O => \N__55420\,
            I => \N__55366\
        );

    \I__13741\ : LocalMux
    port map (
            O => \N__55417\,
            I => \N__55359\
        );

    \I__13740\ : Span4Mux_v
    port map (
            O => \N__55414\,
            I => \N__55359\
        );

    \I__13739\ : Span4Mux_v
    port map (
            O => \N__55411\,
            I => \N__55359\
        );

    \I__13738\ : Span4Mux_h
    port map (
            O => \N__55404\,
            I => \N__55356\
        );

    \I__13737\ : LocalMux
    port map (
            O => \N__55401\,
            I => \N__55353\
        );

    \I__13736\ : InMux
    port map (
            O => \N__55400\,
            I => \N__55348\
        );

    \I__13735\ : InMux
    port map (
            O => \N__55399\,
            I => \N__55348\
        );

    \I__13734\ : Span4Mux_h
    port map (
            O => \N__55396\,
            I => \N__55345\
        );

    \I__13733\ : LocalMux
    port map (
            O => \N__55393\,
            I => \N__55342\
        );

    \I__13732\ : LocalMux
    port map (
            O => \N__55388\,
            I => \N__55337\
        );

    \I__13731\ : Span4Mux_s2_v
    port map (
            O => \N__55383\,
            I => \N__55337\
        );

    \I__13730\ : InMux
    port map (
            O => \N__55382\,
            I => \N__55334\
        );

    \I__13729\ : InMux
    port map (
            O => \N__55381\,
            I => \N__55331\
        );

    \I__13728\ : Span12Mux_h
    port map (
            O => \N__55378\,
            I => \N__55328\
        );

    \I__13727\ : LocalMux
    port map (
            O => \N__55375\,
            I => \N__55325\
        );

    \I__13726\ : Span4Mux_v
    port map (
            O => \N__55366\,
            I => \N__55322\
        );

    \I__13725\ : Span4Mux_h
    port map (
            O => \N__55359\,
            I => \N__55319\
        );

    \I__13724\ : Span4Mux_v
    port map (
            O => \N__55356\,
            I => \N__55316\
        );

    \I__13723\ : Span12Mux_s6_v
    port map (
            O => \N__55353\,
            I => \N__55311\
        );

    \I__13722\ : LocalMux
    port map (
            O => \N__55348\,
            I => \N__55311\
        );

    \I__13721\ : Span4Mux_h
    port map (
            O => \N__55345\,
            I => \N__55306\
        );

    \I__13720\ : Span4Mux_h
    port map (
            O => \N__55342\,
            I => \N__55306\
        );

    \I__13719\ : Span4Mux_h
    port map (
            O => \N__55337\,
            I => \N__55303\
        );

    \I__13718\ : LocalMux
    port map (
            O => \N__55334\,
            I => \opZ0Z_3\
        );

    \I__13717\ : LocalMux
    port map (
            O => \N__55331\,
            I => \opZ0Z_3\
        );

    \I__13716\ : Odrv12
    port map (
            O => \N__55328\,
            I => \opZ0Z_3\
        );

    \I__13715\ : Odrv4
    port map (
            O => \N__55325\,
            I => \opZ0Z_3\
        );

    \I__13714\ : Odrv4
    port map (
            O => \N__55322\,
            I => \opZ0Z_3\
        );

    \I__13713\ : Odrv4
    port map (
            O => \N__55319\,
            I => \opZ0Z_3\
        );

    \I__13712\ : Odrv4
    port map (
            O => \N__55316\,
            I => \opZ0Z_3\
        );

    \I__13711\ : Odrv12
    port map (
            O => \N__55311\,
            I => \opZ0Z_3\
        );

    \I__13710\ : Odrv4
    port map (
            O => \N__55306\,
            I => \opZ0Z_3\
        );

    \I__13709\ : Odrv4
    port map (
            O => \N__55303\,
            I => \opZ0Z_3\
        );

    \I__13708\ : InMux
    port map (
            O => \N__55282\,
            I => \N__55276\
        );

    \I__13707\ : InMux
    port map (
            O => \N__55281\,
            I => \N__55273\
        );

    \I__13706\ : InMux
    port map (
            O => \N__55280\,
            I => \N__55269\
        );

    \I__13705\ : InMux
    port map (
            O => \N__55279\,
            I => \N__55265\
        );

    \I__13704\ : LocalMux
    port map (
            O => \N__55276\,
            I => \N__55256\
        );

    \I__13703\ : LocalMux
    port map (
            O => \N__55273\,
            I => \N__55253\
        );

    \I__13702\ : InMux
    port map (
            O => \N__55272\,
            I => \N__55250\
        );

    \I__13701\ : LocalMux
    port map (
            O => \N__55269\,
            I => \N__55247\
        );

    \I__13700\ : InMux
    port map (
            O => \N__55268\,
            I => \N__55244\
        );

    \I__13699\ : LocalMux
    port map (
            O => \N__55265\,
            I => \N__55241\
        );

    \I__13698\ : InMux
    port map (
            O => \N__55264\,
            I => \N__55238\
        );

    \I__13697\ : InMux
    port map (
            O => \N__55263\,
            I => \N__55235\
        );

    \I__13696\ : InMux
    port map (
            O => \N__55262\,
            I => \N__55231\
        );

    \I__13695\ : InMux
    port map (
            O => \N__55261\,
            I => \N__55227\
        );

    \I__13694\ : InMux
    port map (
            O => \N__55260\,
            I => \N__55224\
        );

    \I__13693\ : CascadeMux
    port map (
            O => \N__55259\,
            I => \N__55217\
        );

    \I__13692\ : Span4Mux_v
    port map (
            O => \N__55256\,
            I => \N__55205\
        );

    \I__13691\ : Span4Mux_h
    port map (
            O => \N__55253\,
            I => \N__55205\
        );

    \I__13690\ : LocalMux
    port map (
            O => \N__55250\,
            I => \N__55205\
        );

    \I__13689\ : Span4Mux_v
    port map (
            O => \N__55247\,
            I => \N__55205\
        );

    \I__13688\ : LocalMux
    port map (
            O => \N__55244\,
            I => \N__55205\
        );

    \I__13687\ : Span4Mux_v
    port map (
            O => \N__55241\,
            I => \N__55202\
        );

    \I__13686\ : LocalMux
    port map (
            O => \N__55238\,
            I => \N__55199\
        );

    \I__13685\ : LocalMux
    port map (
            O => \N__55235\,
            I => \N__55196\
        );

    \I__13684\ : InMux
    port map (
            O => \N__55234\,
            I => \N__55193\
        );

    \I__13683\ : LocalMux
    port map (
            O => \N__55231\,
            I => \N__55189\
        );

    \I__13682\ : InMux
    port map (
            O => \N__55230\,
            I => \N__55186\
        );

    \I__13681\ : LocalMux
    port map (
            O => \N__55227\,
            I => \N__55182\
        );

    \I__13680\ : LocalMux
    port map (
            O => \N__55224\,
            I => \N__55179\
        );

    \I__13679\ : InMux
    port map (
            O => \N__55223\,
            I => \N__55176\
        );

    \I__13678\ : InMux
    port map (
            O => \N__55222\,
            I => \N__55173\
        );

    \I__13677\ : InMux
    port map (
            O => \N__55221\,
            I => \N__55169\
        );

    \I__13676\ : InMux
    port map (
            O => \N__55220\,
            I => \N__55163\
        );

    \I__13675\ : InMux
    port map (
            O => \N__55217\,
            I => \N__55159\
        );

    \I__13674\ : InMux
    port map (
            O => \N__55216\,
            I => \N__55156\
        );

    \I__13673\ : Span4Mux_v
    port map (
            O => \N__55205\,
            I => \N__55153\
        );

    \I__13672\ : Span4Mux_h
    port map (
            O => \N__55202\,
            I => \N__55150\
        );

    \I__13671\ : Span4Mux_h
    port map (
            O => \N__55199\,
            I => \N__55143\
        );

    \I__13670\ : Span4Mux_h
    port map (
            O => \N__55196\,
            I => \N__55143\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__55193\,
            I => \N__55143\
        );

    \I__13668\ : InMux
    port map (
            O => \N__55192\,
            I => \N__55139\
        );

    \I__13667\ : Span4Mux_v
    port map (
            O => \N__55189\,
            I => \N__55133\
        );

    \I__13666\ : LocalMux
    port map (
            O => \N__55186\,
            I => \N__55133\
        );

    \I__13665\ : InMux
    port map (
            O => \N__55185\,
            I => \N__55130\
        );

    \I__13664\ : Span4Mux_v
    port map (
            O => \N__55182\,
            I => \N__55123\
        );

    \I__13663\ : Span4Mux_h
    port map (
            O => \N__55179\,
            I => \N__55123\
        );

    \I__13662\ : LocalMux
    port map (
            O => \N__55176\,
            I => \N__55123\
        );

    \I__13661\ : LocalMux
    port map (
            O => \N__55173\,
            I => \N__55120\
        );

    \I__13660\ : InMux
    port map (
            O => \N__55172\,
            I => \N__55117\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__55169\,
            I => \N__55114\
        );

    \I__13658\ : InMux
    port map (
            O => \N__55168\,
            I => \N__55111\
        );

    \I__13657\ : InMux
    port map (
            O => \N__55167\,
            I => \N__55108\
        );

    \I__13656\ : InMux
    port map (
            O => \N__55166\,
            I => \N__55105\
        );

    \I__13655\ : LocalMux
    port map (
            O => \N__55163\,
            I => \N__55102\
        );

    \I__13654\ : InMux
    port map (
            O => \N__55162\,
            I => \N__55099\
        );

    \I__13653\ : LocalMux
    port map (
            O => \N__55159\,
            I => \N__55095\
        );

    \I__13652\ : LocalMux
    port map (
            O => \N__55156\,
            I => \N__55092\
        );

    \I__13651\ : Span4Mux_h
    port map (
            O => \N__55153\,
            I => \N__55085\
        );

    \I__13650\ : Span4Mux_h
    port map (
            O => \N__55150\,
            I => \N__55085\
        );

    \I__13649\ : Span4Mux_v
    port map (
            O => \N__55143\,
            I => \N__55085\
        );

    \I__13648\ : InMux
    port map (
            O => \N__55142\,
            I => \N__55082\
        );

    \I__13647\ : LocalMux
    port map (
            O => \N__55139\,
            I => \N__55079\
        );

    \I__13646\ : InMux
    port map (
            O => \N__55138\,
            I => \N__55076\
        );

    \I__13645\ : Span4Mux_v
    port map (
            O => \N__55133\,
            I => \N__55073\
        );

    \I__13644\ : LocalMux
    port map (
            O => \N__55130\,
            I => \N__55068\
        );

    \I__13643\ : Span4Mux_v
    port map (
            O => \N__55123\,
            I => \N__55065\
        );

    \I__13642\ : Span4Mux_h
    port map (
            O => \N__55120\,
            I => \N__55062\
        );

    \I__13641\ : LocalMux
    port map (
            O => \N__55117\,
            I => \N__55057\
        );

    \I__13640\ : Span4Mux_h
    port map (
            O => \N__55114\,
            I => \N__55057\
        );

    \I__13639\ : LocalMux
    port map (
            O => \N__55111\,
            I => \N__55048\
        );

    \I__13638\ : LocalMux
    port map (
            O => \N__55108\,
            I => \N__55048\
        );

    \I__13637\ : LocalMux
    port map (
            O => \N__55105\,
            I => \N__55048\
        );

    \I__13636\ : Sp12to4
    port map (
            O => \N__55102\,
            I => \N__55048\
        );

    \I__13635\ : LocalMux
    port map (
            O => \N__55099\,
            I => \N__55045\
        );

    \I__13634\ : InMux
    port map (
            O => \N__55098\,
            I => \N__55042\
        );

    \I__13633\ : Span12Mux_s4_h
    port map (
            O => \N__55095\,
            I => \N__55035\
        );

    \I__13632\ : Span12Mux_v
    port map (
            O => \N__55092\,
            I => \N__55035\
        );

    \I__13631\ : Sp12to4
    port map (
            O => \N__55085\,
            I => \N__55035\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__55082\,
            I => \N__55030\
        );

    \I__13629\ : Span4Mux_h
    port map (
            O => \N__55079\,
            I => \N__55030\
        );

    \I__13628\ : LocalMux
    port map (
            O => \N__55076\,
            I => \N__55027\
        );

    \I__13627\ : Span4Mux_h
    port map (
            O => \N__55073\,
            I => \N__55024\
        );

    \I__13626\ : InMux
    port map (
            O => \N__55072\,
            I => \N__55021\
        );

    \I__13625\ : InMux
    port map (
            O => \N__55071\,
            I => \N__55018\
        );

    \I__13624\ : Span4Mux_h
    port map (
            O => \N__55068\,
            I => \N__55015\
        );

    \I__13623\ : Span4Mux_v
    port map (
            O => \N__55065\,
            I => \N__55008\
        );

    \I__13622\ : Span4Mux_v
    port map (
            O => \N__55062\,
            I => \N__55008\
        );

    \I__13621\ : Span4Mux_v
    port map (
            O => \N__55057\,
            I => \N__55008\
        );

    \I__13620\ : Span12Mux_v
    port map (
            O => \N__55048\,
            I => \N__55003\
        );

    \I__13619\ : Span12Mux_s6_h
    port map (
            O => \N__55045\,
            I => \N__55003\
        );

    \I__13618\ : LocalMux
    port map (
            O => \N__55042\,
            I => \N__54998\
        );

    \I__13617\ : Span12Mux_h
    port map (
            O => \N__55035\,
            I => \N__54998\
        );

    \I__13616\ : Span4Mux_v
    port map (
            O => \N__55030\,
            I => \N__54991\
        );

    \I__13615\ : Span4Mux_h
    port map (
            O => \N__55027\,
            I => \N__54991\
        );

    \I__13614\ : Span4Mux_h
    port map (
            O => \N__55024\,
            I => \N__54991\
        );

    \I__13613\ : LocalMux
    port map (
            O => \N__55021\,
            I => \opZ0Z_1\
        );

    \I__13612\ : LocalMux
    port map (
            O => \N__55018\,
            I => \opZ0Z_1\
        );

    \I__13611\ : Odrv4
    port map (
            O => \N__55015\,
            I => \opZ0Z_1\
        );

    \I__13610\ : Odrv4
    port map (
            O => \N__55008\,
            I => \opZ0Z_1\
        );

    \I__13609\ : Odrv12
    port map (
            O => \N__55003\,
            I => \opZ0Z_1\
        );

    \I__13608\ : Odrv12
    port map (
            O => \N__54998\,
            I => \opZ0Z_1\
        );

    \I__13607\ : Odrv4
    port map (
            O => \N__54991\,
            I => \opZ0Z_1\
        );

    \I__13606\ : CascadeMux
    port map (
            O => \N__54976\,
            I => \ALU.un1_op_1Z0Z_1_cascade_\
        );

    \I__13605\ : InMux
    port map (
            O => \N__54973\,
            I => \N__54969\
        );

    \I__13604\ : InMux
    port map (
            O => \N__54972\,
            I => \N__54966\
        );

    \I__13603\ : LocalMux
    port map (
            O => \N__54969\,
            I => \opZ0Z_4\
        );

    \I__13602\ : LocalMux
    port map (
            O => \N__54966\,
            I => \opZ0Z_4\
        );

    \I__13601\ : InMux
    port map (
            O => \N__54961\,
            I => \N__54940\
        );

    \I__13600\ : InMux
    port map (
            O => \N__54960\,
            I => \N__54940\
        );

    \I__13599\ : InMux
    port map (
            O => \N__54959\,
            I => \N__54940\
        );

    \I__13598\ : InMux
    port map (
            O => \N__54958\,
            I => \N__54940\
        );

    \I__13597\ : InMux
    port map (
            O => \N__54957\,
            I => \N__54940\
        );

    \I__13596\ : InMux
    port map (
            O => \N__54956\,
            I => \N__54940\
        );

    \I__13595\ : InMux
    port map (
            O => \N__54955\,
            I => \N__54940\
        );

    \I__13594\ : LocalMux
    port map (
            O => \N__54940\,
            I => \N__54937\
        );

    \I__13593\ : Span4Mux_h
    port map (
            O => \N__54937\,
            I => \N__54933\
        );

    \I__13592\ : InMux
    port map (
            O => \N__54936\,
            I => \N__54930\
        );

    \I__13591\ : Odrv4
    port map (
            O => \N__54933\,
            I => \ALU.un1_op_1_0\
        );

    \I__13590\ : LocalMux
    port map (
            O => \N__54930\,
            I => \ALU.un1_op_1_0\
        );

    \I__13589\ : InMux
    port map (
            O => \N__54925\,
            I => \N__54916\
        );

    \I__13588\ : CascadeMux
    port map (
            O => \N__54924\,
            I => \N__54911\
        );

    \I__13587\ : CascadeMux
    port map (
            O => \N__54923\,
            I => \N__54908\
        );

    \I__13586\ : InMux
    port map (
            O => \N__54922\,
            I => \N__54902\
        );

    \I__13585\ : CascadeMux
    port map (
            O => \N__54921\,
            I => \N__54895\
        );

    \I__13584\ : CascadeMux
    port map (
            O => \N__54920\,
            I => \N__54891\
        );

    \I__13583\ : InMux
    port map (
            O => \N__54919\,
            I => \N__54881\
        );

    \I__13582\ : LocalMux
    port map (
            O => \N__54916\,
            I => \N__54878\
        );

    \I__13581\ : InMux
    port map (
            O => \N__54915\,
            I => \N__54871\
        );

    \I__13580\ : InMux
    port map (
            O => \N__54914\,
            I => \N__54871\
        );

    \I__13579\ : InMux
    port map (
            O => \N__54911\,
            I => \N__54871\
        );

    \I__13578\ : InMux
    port map (
            O => \N__54908\,
            I => \N__54864\
        );

    \I__13577\ : InMux
    port map (
            O => \N__54907\,
            I => \N__54864\
        );

    \I__13576\ : InMux
    port map (
            O => \N__54906\,
            I => \N__54864\
        );

    \I__13575\ : InMux
    port map (
            O => \N__54905\,
            I => \N__54861\
        );

    \I__13574\ : LocalMux
    port map (
            O => \N__54902\,
            I => \N__54855\
        );

    \I__13573\ : InMux
    port map (
            O => \N__54901\,
            I => \N__54850\
        );

    \I__13572\ : InMux
    port map (
            O => \N__54900\,
            I => \N__54850\
        );

    \I__13571\ : InMux
    port map (
            O => \N__54899\,
            I => \N__54843\
        );

    \I__13570\ : InMux
    port map (
            O => \N__54898\,
            I => \N__54843\
        );

    \I__13569\ : InMux
    port map (
            O => \N__54895\,
            I => \N__54843\
        );

    \I__13568\ : InMux
    port map (
            O => \N__54894\,
            I => \N__54838\
        );

    \I__13567\ : InMux
    port map (
            O => \N__54891\,
            I => \N__54838\
        );

    \I__13566\ : InMux
    port map (
            O => \N__54890\,
            I => \N__54830\
        );

    \I__13565\ : CascadeMux
    port map (
            O => \N__54889\,
            I => \N__54824\
        );

    \I__13564\ : CascadeMux
    port map (
            O => \N__54888\,
            I => \N__54818\
        );

    \I__13563\ : CascadeMux
    port map (
            O => \N__54887\,
            I => \N__54814\
        );

    \I__13562\ : CascadeMux
    port map (
            O => \N__54886\,
            I => \N__54807\
        );

    \I__13561\ : CascadeMux
    port map (
            O => \N__54885\,
            I => \N__54797\
        );

    \I__13560\ : CascadeMux
    port map (
            O => \N__54884\,
            I => \N__54792\
        );

    \I__13559\ : LocalMux
    port map (
            O => \N__54881\,
            I => \N__54770\
        );

    \I__13558\ : Span4Mux_h
    port map (
            O => \N__54878\,
            I => \N__54770\
        );

    \I__13557\ : LocalMux
    port map (
            O => \N__54871\,
            I => \N__54770\
        );

    \I__13556\ : LocalMux
    port map (
            O => \N__54864\,
            I => \N__54765\
        );

    \I__13555\ : LocalMux
    port map (
            O => \N__54861\,
            I => \N__54765\
        );

    \I__13554\ : InMux
    port map (
            O => \N__54860\,
            I => \N__54760\
        );

    \I__13553\ : InMux
    port map (
            O => \N__54859\,
            I => \N__54760\
        );

    \I__13552\ : InMux
    port map (
            O => \N__54858\,
            I => \N__54757\
        );

    \I__13551\ : Span4Mux_v
    port map (
            O => \N__54855\,
            I => \N__54754\
        );

    \I__13550\ : LocalMux
    port map (
            O => \N__54850\,
            I => \N__54749\
        );

    \I__13549\ : LocalMux
    port map (
            O => \N__54843\,
            I => \N__54749\
        );

    \I__13548\ : LocalMux
    port map (
            O => \N__54838\,
            I => \N__54746\
        );

    \I__13547\ : InMux
    port map (
            O => \N__54837\,
            I => \N__54739\
        );

    \I__13546\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54739\
        );

    \I__13545\ : InMux
    port map (
            O => \N__54835\,
            I => \N__54739\
        );

    \I__13544\ : InMux
    port map (
            O => \N__54834\,
            I => \N__54734\
        );

    \I__13543\ : InMux
    port map (
            O => \N__54833\,
            I => \N__54734\
        );

    \I__13542\ : LocalMux
    port map (
            O => \N__54830\,
            I => \N__54731\
        );

    \I__13541\ : InMux
    port map (
            O => \N__54829\,
            I => \N__54728\
        );

    \I__13540\ : InMux
    port map (
            O => \N__54828\,
            I => \N__54725\
        );

    \I__13539\ : InMux
    port map (
            O => \N__54827\,
            I => \N__54720\
        );

    \I__13538\ : InMux
    port map (
            O => \N__54824\,
            I => \N__54720\
        );

    \I__13537\ : CascadeMux
    port map (
            O => \N__54823\,
            I => \N__54715\
        );

    \I__13536\ : InMux
    port map (
            O => \N__54822\,
            I => \N__54708\
        );

    \I__13535\ : InMux
    port map (
            O => \N__54821\,
            I => \N__54708\
        );

    \I__13534\ : InMux
    port map (
            O => \N__54818\,
            I => \N__54708\
        );

    \I__13533\ : InMux
    port map (
            O => \N__54817\,
            I => \N__54703\
        );

    \I__13532\ : InMux
    port map (
            O => \N__54814\,
            I => \N__54703\
        );

    \I__13531\ : CascadeMux
    port map (
            O => \N__54813\,
            I => \N__54698\
        );

    \I__13530\ : InMux
    port map (
            O => \N__54812\,
            I => \N__54694\
        );

    \I__13529\ : InMux
    port map (
            O => \N__54811\,
            I => \N__54691\
        );

    \I__13528\ : InMux
    port map (
            O => \N__54810\,
            I => \N__54686\
        );

    \I__13527\ : InMux
    port map (
            O => \N__54807\,
            I => \N__54686\
        );

    \I__13526\ : InMux
    port map (
            O => \N__54806\,
            I => \N__54681\
        );

    \I__13525\ : InMux
    port map (
            O => \N__54805\,
            I => \N__54681\
        );

    \I__13524\ : InMux
    port map (
            O => \N__54804\,
            I => \N__54672\
        );

    \I__13523\ : InMux
    port map (
            O => \N__54803\,
            I => \N__54672\
        );

    \I__13522\ : InMux
    port map (
            O => \N__54802\,
            I => \N__54672\
        );

    \I__13521\ : InMux
    port map (
            O => \N__54801\,
            I => \N__54672\
        );

    \I__13520\ : CascadeMux
    port map (
            O => \N__54800\,
            I => \N__54669\
        );

    \I__13519\ : InMux
    port map (
            O => \N__54797\,
            I => \N__54664\
        );

    \I__13518\ : InMux
    port map (
            O => \N__54796\,
            I => \N__54664\
        );

    \I__13517\ : InMux
    port map (
            O => \N__54795\,
            I => \N__54659\
        );

    \I__13516\ : InMux
    port map (
            O => \N__54792\,
            I => \N__54659\
        );

    \I__13515\ : CascadeMux
    port map (
            O => \N__54791\,
            I => \N__54655\
        );

    \I__13514\ : CascadeMux
    port map (
            O => \N__54790\,
            I => \N__54652\
        );

    \I__13513\ : CascadeMux
    port map (
            O => \N__54789\,
            I => \N__54648\
        );

    \I__13512\ : CascadeMux
    port map (
            O => \N__54788\,
            I => \N__54645\
        );

    \I__13511\ : CascadeMux
    port map (
            O => \N__54787\,
            I => \N__54642\
        );

    \I__13510\ : InMux
    port map (
            O => \N__54786\,
            I => \N__54633\
        );

    \I__13509\ : InMux
    port map (
            O => \N__54785\,
            I => \N__54633\
        );

    \I__13508\ : CascadeMux
    port map (
            O => \N__54784\,
            I => \N__54622\
        );

    \I__13507\ : InMux
    port map (
            O => \N__54783\,
            I => \N__54619\
        );

    \I__13506\ : InMux
    port map (
            O => \N__54782\,
            I => \N__54612\
        );

    \I__13505\ : CascadeMux
    port map (
            O => \N__54781\,
            I => \N__54608\
        );

    \I__13504\ : CascadeMux
    port map (
            O => \N__54780\,
            I => \N__54600\
        );

    \I__13503\ : CascadeMux
    port map (
            O => \N__54779\,
            I => \N__54597\
        );

    \I__13502\ : CascadeMux
    port map (
            O => \N__54778\,
            I => \N__54587\
        );

    \I__13501\ : CascadeMux
    port map (
            O => \N__54777\,
            I => \N__54577\
        );

    \I__13500\ : Span4Mux_v
    port map (
            O => \N__54770\,
            I => \N__54568\
        );

    \I__13499\ : Span4Mux_v
    port map (
            O => \N__54765\,
            I => \N__54568\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__54760\,
            I => \N__54568\
        );

    \I__13497\ : LocalMux
    port map (
            O => \N__54757\,
            I => \N__54568\
        );

    \I__13496\ : Span4Mux_h
    port map (
            O => \N__54754\,
            I => \N__54563\
        );

    \I__13495\ : Span4Mux_v
    port map (
            O => \N__54749\,
            I => \N__54563\
        );

    \I__13494\ : Span4Mux_s3_v
    port map (
            O => \N__54746\,
            I => \N__54558\
        );

    \I__13493\ : LocalMux
    port map (
            O => \N__54739\,
            I => \N__54558\
        );

    \I__13492\ : LocalMux
    port map (
            O => \N__54734\,
            I => \N__54547\
        );

    \I__13491\ : Span4Mux_v
    port map (
            O => \N__54731\,
            I => \N__54547\
        );

    \I__13490\ : LocalMux
    port map (
            O => \N__54728\,
            I => \N__54540\
        );

    \I__13489\ : LocalMux
    port map (
            O => \N__54725\,
            I => \N__54540\
        );

    \I__13488\ : LocalMux
    port map (
            O => \N__54720\,
            I => \N__54540\
        );

    \I__13487\ : InMux
    port map (
            O => \N__54719\,
            I => \N__54533\
        );

    \I__13486\ : InMux
    port map (
            O => \N__54718\,
            I => \N__54533\
        );

    \I__13485\ : InMux
    port map (
            O => \N__54715\,
            I => \N__54533\
        );

    \I__13484\ : LocalMux
    port map (
            O => \N__54708\,
            I => \N__54528\
        );

    \I__13483\ : LocalMux
    port map (
            O => \N__54703\,
            I => \N__54528\
        );

    \I__13482\ : InMux
    port map (
            O => \N__54702\,
            I => \N__54521\
        );

    \I__13481\ : InMux
    port map (
            O => \N__54701\,
            I => \N__54521\
        );

    \I__13480\ : InMux
    port map (
            O => \N__54698\,
            I => \N__54521\
        );

    \I__13479\ : CascadeMux
    port map (
            O => \N__54697\,
            I => \N__54517\
        );

    \I__13478\ : LocalMux
    port map (
            O => \N__54694\,
            I => \N__54512\
        );

    \I__13477\ : LocalMux
    port map (
            O => \N__54691\,
            I => \N__54512\
        );

    \I__13476\ : LocalMux
    port map (
            O => \N__54686\,
            I => \N__54509\
        );

    \I__13475\ : LocalMux
    port map (
            O => \N__54681\,
            I => \N__54504\
        );

    \I__13474\ : LocalMux
    port map (
            O => \N__54672\,
            I => \N__54504\
        );

    \I__13473\ : InMux
    port map (
            O => \N__54669\,
            I => \N__54501\
        );

    \I__13472\ : LocalMux
    port map (
            O => \N__54664\,
            I => \N__54496\
        );

    \I__13471\ : LocalMux
    port map (
            O => \N__54659\,
            I => \N__54496\
        );

    \I__13470\ : InMux
    port map (
            O => \N__54658\,
            I => \N__54489\
        );

    \I__13469\ : InMux
    port map (
            O => \N__54655\,
            I => \N__54489\
        );

    \I__13468\ : InMux
    port map (
            O => \N__54652\,
            I => \N__54489\
        );

    \I__13467\ : InMux
    port map (
            O => \N__54651\,
            I => \N__54484\
        );

    \I__13466\ : InMux
    port map (
            O => \N__54648\,
            I => \N__54484\
        );

    \I__13465\ : InMux
    port map (
            O => \N__54645\,
            I => \N__54479\
        );

    \I__13464\ : InMux
    port map (
            O => \N__54642\,
            I => \N__54479\
        );

    \I__13463\ : InMux
    port map (
            O => \N__54641\,
            I => \N__54475\
        );

    \I__13462\ : InMux
    port map (
            O => \N__54640\,
            I => \N__54470\
        );

    \I__13461\ : InMux
    port map (
            O => \N__54639\,
            I => \N__54470\
        );

    \I__13460\ : CascadeMux
    port map (
            O => \N__54638\,
            I => \N__54467\
        );

    \I__13459\ : LocalMux
    port map (
            O => \N__54633\,
            I => \N__54464\
        );

    \I__13458\ : InMux
    port map (
            O => \N__54632\,
            I => \N__54461\
        );

    \I__13457\ : InMux
    port map (
            O => \N__54631\,
            I => \N__54448\
        );

    \I__13456\ : InMux
    port map (
            O => \N__54630\,
            I => \N__54448\
        );

    \I__13455\ : InMux
    port map (
            O => \N__54629\,
            I => \N__54448\
        );

    \I__13454\ : InMux
    port map (
            O => \N__54628\,
            I => \N__54448\
        );

    \I__13453\ : InMux
    port map (
            O => \N__54627\,
            I => \N__54448\
        );

    \I__13452\ : InMux
    port map (
            O => \N__54626\,
            I => \N__54448\
        );

    \I__13451\ : InMux
    port map (
            O => \N__54625\,
            I => \N__54442\
        );

    \I__13450\ : InMux
    port map (
            O => \N__54622\,
            I => \N__54442\
        );

    \I__13449\ : LocalMux
    port map (
            O => \N__54619\,
            I => \N__54439\
        );

    \I__13448\ : InMux
    port map (
            O => \N__54618\,
            I => \N__54432\
        );

    \I__13447\ : InMux
    port map (
            O => \N__54617\,
            I => \N__54432\
        );

    \I__13446\ : InMux
    port map (
            O => \N__54616\,
            I => \N__54432\
        );

    \I__13445\ : InMux
    port map (
            O => \N__54615\,
            I => \N__54429\
        );

    \I__13444\ : LocalMux
    port map (
            O => \N__54612\,
            I => \N__54426\
        );

    \I__13443\ : InMux
    port map (
            O => \N__54611\,
            I => \N__54423\
        );

    \I__13442\ : InMux
    port map (
            O => \N__54608\,
            I => \N__54420\
        );

    \I__13441\ : CascadeMux
    port map (
            O => \N__54607\,
            I => \N__54417\
        );

    \I__13440\ : InMux
    port map (
            O => \N__54606\,
            I => \N__54414\
        );

    \I__13439\ : InMux
    port map (
            O => \N__54605\,
            I => \N__54409\
        );

    \I__13438\ : InMux
    port map (
            O => \N__54604\,
            I => \N__54409\
        );

    \I__13437\ : InMux
    port map (
            O => \N__54603\,
            I => \N__54406\
        );

    \I__13436\ : InMux
    port map (
            O => \N__54600\,
            I => \N__54403\
        );

    \I__13435\ : InMux
    port map (
            O => \N__54597\,
            I => \N__54396\
        );

    \I__13434\ : InMux
    port map (
            O => \N__54596\,
            I => \N__54396\
        );

    \I__13433\ : InMux
    port map (
            O => \N__54595\,
            I => \N__54396\
        );

    \I__13432\ : InMux
    port map (
            O => \N__54594\,
            I => \N__54393\
        );

    \I__13431\ : InMux
    port map (
            O => \N__54593\,
            I => \N__54384\
        );

    \I__13430\ : InMux
    port map (
            O => \N__54592\,
            I => \N__54384\
        );

    \I__13429\ : InMux
    port map (
            O => \N__54591\,
            I => \N__54384\
        );

    \I__13428\ : InMux
    port map (
            O => \N__54590\,
            I => \N__54384\
        );

    \I__13427\ : InMux
    port map (
            O => \N__54587\,
            I => \N__54376\
        );

    \I__13426\ : InMux
    port map (
            O => \N__54586\,
            I => \N__54376\
        );

    \I__13425\ : InMux
    port map (
            O => \N__54585\,
            I => \N__54376\
        );

    \I__13424\ : InMux
    port map (
            O => \N__54584\,
            I => \N__54373\
        );

    \I__13423\ : InMux
    port map (
            O => \N__54583\,
            I => \N__54370\
        );

    \I__13422\ : InMux
    port map (
            O => \N__54582\,
            I => \N__54365\
        );

    \I__13421\ : InMux
    port map (
            O => \N__54581\,
            I => \N__54365\
        );

    \I__13420\ : InMux
    port map (
            O => \N__54580\,
            I => \N__54362\
        );

    \I__13419\ : InMux
    port map (
            O => \N__54577\,
            I => \N__54359\
        );

    \I__13418\ : Span4Mux_h
    port map (
            O => \N__54568\,
            I => \N__54352\
        );

    \I__13417\ : Span4Mux_h
    port map (
            O => \N__54563\,
            I => \N__54352\
        );

    \I__13416\ : Span4Mux_v
    port map (
            O => \N__54558\,
            I => \N__54352\
        );

    \I__13415\ : CascadeMux
    port map (
            O => \N__54557\,
            I => \N__54349\
        );

    \I__13414\ : InMux
    port map (
            O => \N__54556\,
            I => \N__54346\
        );

    \I__13413\ : InMux
    port map (
            O => \N__54555\,
            I => \N__54343\
        );

    \I__13412\ : InMux
    port map (
            O => \N__54554\,
            I => \N__54338\
        );

    \I__13411\ : InMux
    port map (
            O => \N__54553\,
            I => \N__54338\
        );

    \I__13410\ : InMux
    port map (
            O => \N__54552\,
            I => \N__54335\
        );

    \I__13409\ : Span4Mux_v
    port map (
            O => \N__54547\,
            I => \N__54328\
        );

    \I__13408\ : Span4Mux_v
    port map (
            O => \N__54540\,
            I => \N__54328\
        );

    \I__13407\ : LocalMux
    port map (
            O => \N__54533\,
            I => \N__54328\
        );

    \I__13406\ : Span4Mux_h
    port map (
            O => \N__54528\,
            I => \N__54325\
        );

    \I__13405\ : LocalMux
    port map (
            O => \N__54521\,
            I => \N__54322\
        );

    \I__13404\ : InMux
    port map (
            O => \N__54520\,
            I => \N__54319\
        );

    \I__13403\ : InMux
    port map (
            O => \N__54517\,
            I => \N__54316\
        );

    \I__13402\ : Span4Mux_h
    port map (
            O => \N__54512\,
            I => \N__54301\
        );

    \I__13401\ : Span4Mux_s2_v
    port map (
            O => \N__54509\,
            I => \N__54301\
        );

    \I__13400\ : Span4Mux_s2_v
    port map (
            O => \N__54504\,
            I => \N__54301\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__54501\,
            I => \N__54301\
        );

    \I__13398\ : Span4Mux_v
    port map (
            O => \N__54496\,
            I => \N__54301\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__54489\,
            I => \N__54301\
        );

    \I__13396\ : LocalMux
    port map (
            O => \N__54484\,
            I => \N__54301\
        );

    \I__13395\ : LocalMux
    port map (
            O => \N__54479\,
            I => \N__54298\
        );

    \I__13394\ : CascadeMux
    port map (
            O => \N__54478\,
            I => \N__54295\
        );

    \I__13393\ : LocalMux
    port map (
            O => \N__54475\,
            I => \N__54290\
        );

    \I__13392\ : LocalMux
    port map (
            O => \N__54470\,
            I => \N__54290\
        );

    \I__13391\ : InMux
    port map (
            O => \N__54467\,
            I => \N__54287\
        );

    \I__13390\ : Span4Mux_s2_v
    port map (
            O => \N__54464\,
            I => \N__54280\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__54461\,
            I => \N__54280\
        );

    \I__13388\ : LocalMux
    port map (
            O => \N__54448\,
            I => \N__54280\
        );

    \I__13387\ : InMux
    port map (
            O => \N__54447\,
            I => \N__54277\
        );

    \I__13386\ : LocalMux
    port map (
            O => \N__54442\,
            I => \N__54274\
        );

    \I__13385\ : Span4Mux_s2_v
    port map (
            O => \N__54439\,
            I => \N__54269\
        );

    \I__13384\ : LocalMux
    port map (
            O => \N__54432\,
            I => \N__54269\
        );

    \I__13383\ : LocalMux
    port map (
            O => \N__54429\,
            I => \N__54260\
        );

    \I__13382\ : Span4Mux_h
    port map (
            O => \N__54426\,
            I => \N__54260\
        );

    \I__13381\ : LocalMux
    port map (
            O => \N__54423\,
            I => \N__54260\
        );

    \I__13380\ : LocalMux
    port map (
            O => \N__54420\,
            I => \N__54260\
        );

    \I__13379\ : InMux
    port map (
            O => \N__54417\,
            I => \N__54257\
        );

    \I__13378\ : LocalMux
    port map (
            O => \N__54414\,
            I => \N__54250\
        );

    \I__13377\ : LocalMux
    port map (
            O => \N__54409\,
            I => \N__54250\
        );

    \I__13376\ : LocalMux
    port map (
            O => \N__54406\,
            I => \N__54250\
        );

    \I__13375\ : LocalMux
    port map (
            O => \N__54403\,
            I => \N__54247\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__54396\,
            I => \N__54244\
        );

    \I__13373\ : LocalMux
    port map (
            O => \N__54393\,
            I => \N__54239\
        );

    \I__13372\ : LocalMux
    port map (
            O => \N__54384\,
            I => \N__54239\
        );

    \I__13371\ : InMux
    port map (
            O => \N__54383\,
            I => \N__54236\
        );

    \I__13370\ : LocalMux
    port map (
            O => \N__54376\,
            I => \N__54233\
        );

    \I__13369\ : LocalMux
    port map (
            O => \N__54373\,
            I => \N__54230\
        );

    \I__13368\ : LocalMux
    port map (
            O => \N__54370\,
            I => \N__54219\
        );

    \I__13367\ : LocalMux
    port map (
            O => \N__54365\,
            I => \N__54219\
        );

    \I__13366\ : LocalMux
    port map (
            O => \N__54362\,
            I => \N__54219\
        );

    \I__13365\ : LocalMux
    port map (
            O => \N__54359\,
            I => \N__54219\
        );

    \I__13364\ : Span4Mux_v
    port map (
            O => \N__54352\,
            I => \N__54219\
        );

    \I__13363\ : InMux
    port map (
            O => \N__54349\,
            I => \N__54216\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__54346\,
            I => \N__54212\
        );

    \I__13361\ : LocalMux
    port map (
            O => \N__54343\,
            I => \N__54209\
        );

    \I__13360\ : LocalMux
    port map (
            O => \N__54338\,
            I => \N__54204\
        );

    \I__13359\ : LocalMux
    port map (
            O => \N__54335\,
            I => \N__54204\
        );

    \I__13358\ : Span4Mux_h
    port map (
            O => \N__54328\,
            I => \N__54193\
        );

    \I__13357\ : Span4Mux_v
    port map (
            O => \N__54325\,
            I => \N__54193\
        );

    \I__13356\ : Span4Mux_v
    port map (
            O => \N__54322\,
            I => \N__54193\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__54319\,
            I => \N__54193\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__54316\,
            I => \N__54193\
        );

    \I__13353\ : Span4Mux_h
    port map (
            O => \N__54301\,
            I => \N__54188\
        );

    \I__13352\ : Span4Mux_s2_v
    port map (
            O => \N__54298\,
            I => \N__54188\
        );

    \I__13351\ : InMux
    port map (
            O => \N__54295\,
            I => \N__54185\
        );

    \I__13350\ : Span4Mux_v
    port map (
            O => \N__54290\,
            I => \N__54178\
        );

    \I__13349\ : LocalMux
    port map (
            O => \N__54287\,
            I => \N__54178\
        );

    \I__13348\ : Span4Mux_v
    port map (
            O => \N__54280\,
            I => \N__54178\
        );

    \I__13347\ : LocalMux
    port map (
            O => \N__54277\,
            I => \N__54167\
        );

    \I__13346\ : Span4Mux_h
    port map (
            O => \N__54274\,
            I => \N__54167\
        );

    \I__13345\ : Span4Mux_v
    port map (
            O => \N__54269\,
            I => \N__54167\
        );

    \I__13344\ : Span4Mux_v
    port map (
            O => \N__54260\,
            I => \N__54167\
        );

    \I__13343\ : LocalMux
    port map (
            O => \N__54257\,
            I => \N__54167\
        );

    \I__13342\ : Span4Mux_v
    port map (
            O => \N__54250\,
            I => \N__54164\
        );

    \I__13341\ : Span4Mux_h
    port map (
            O => \N__54247\,
            I => \N__54155\
        );

    \I__13340\ : Span4Mux_h
    port map (
            O => \N__54244\,
            I => \N__54155\
        );

    \I__13339\ : Span4Mux_v
    port map (
            O => \N__54239\,
            I => \N__54155\
        );

    \I__13338\ : LocalMux
    port map (
            O => \N__54236\,
            I => \N__54155\
        );

    \I__13337\ : Span4Mux_v
    port map (
            O => \N__54233\,
            I => \N__54152\
        );

    \I__13336\ : Span4Mux_h
    port map (
            O => \N__54230\,
            I => \N__54145\
        );

    \I__13335\ : Span4Mux_v
    port map (
            O => \N__54219\,
            I => \N__54145\
        );

    \I__13334\ : LocalMux
    port map (
            O => \N__54216\,
            I => \N__54145\
        );

    \I__13333\ : CascadeMux
    port map (
            O => \N__54215\,
            I => \N__54142\
        );

    \I__13332\ : Span4Mux_s0_v
    port map (
            O => \N__54212\,
            I => \N__54133\
        );

    \I__13331\ : Span4Mux_h
    port map (
            O => \N__54209\,
            I => \N__54133\
        );

    \I__13330\ : Span4Mux_h
    port map (
            O => \N__54204\,
            I => \N__54133\
        );

    \I__13329\ : Span4Mux_h
    port map (
            O => \N__54193\,
            I => \N__54133\
        );

    \I__13328\ : Span4Mux_h
    port map (
            O => \N__54188\,
            I => \N__54130\
        );

    \I__13327\ : LocalMux
    port map (
            O => \N__54185\,
            I => \N__54125\
        );

    \I__13326\ : Span4Mux_h
    port map (
            O => \N__54178\,
            I => \N__54120\
        );

    \I__13325\ : Span4Mux_v
    port map (
            O => \N__54167\,
            I => \N__54120\
        );

    \I__13324\ : Span4Mux_h
    port map (
            O => \N__54164\,
            I => \N__54111\
        );

    \I__13323\ : Span4Mux_v
    port map (
            O => \N__54155\,
            I => \N__54111\
        );

    \I__13322\ : Span4Mux_h
    port map (
            O => \N__54152\,
            I => \N__54111\
        );

    \I__13321\ : Span4Mux_h
    port map (
            O => \N__54145\,
            I => \N__54111\
        );

    \I__13320\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54108\
        );

    \I__13319\ : Sp12to4
    port map (
            O => \N__54133\,
            I => \N__54105\
        );

    \I__13318\ : Span4Mux_v
    port map (
            O => \N__54130\,
            I => \N__54102\
        );

    \I__13317\ : InMux
    port map (
            O => \N__54129\,
            I => \N__54099\
        );

    \I__13316\ : InMux
    port map (
            O => \N__54128\,
            I => \N__54096\
        );

    \I__13315\ : Span4Mux_v
    port map (
            O => \N__54125\,
            I => \N__54091\
        );

    \I__13314\ : Span4Mux_h
    port map (
            O => \N__54120\,
            I => \N__54091\
        );

    \I__13313\ : Span4Mux_v
    port map (
            O => \N__54111\,
            I => \N__54086\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__54108\,
            I => \N__54086\
        );

    \I__13311\ : Span12Mux_s6_v
    port map (
            O => \N__54105\,
            I => \N__54081\
        );

    \I__13310\ : Sp12to4
    port map (
            O => \N__54102\,
            I => \N__54081\
        );

    \I__13309\ : LocalMux
    port map (
            O => \N__54099\,
            I => \paramsZ0Z_1\
        );

    \I__13308\ : LocalMux
    port map (
            O => \N__54096\,
            I => \paramsZ0Z_1\
        );

    \I__13307\ : Odrv4
    port map (
            O => \N__54091\,
            I => \paramsZ0Z_1\
        );

    \I__13306\ : Odrv4
    port map (
            O => \N__54086\,
            I => \paramsZ0Z_1\
        );

    \I__13305\ : Odrv12
    port map (
            O => \N__54081\,
            I => \paramsZ0Z_1\
        );

    \I__13304\ : CascadeMux
    port map (
            O => \N__54070\,
            I => \N__54066\
        );

    \I__13303\ : CascadeMux
    port map (
            O => \N__54069\,
            I => \N__54063\
        );

    \I__13302\ : InMux
    port map (
            O => \N__54066\,
            I => \N__54042\
        );

    \I__13301\ : InMux
    port map (
            O => \N__54063\,
            I => \N__54042\
        );

    \I__13300\ : InMux
    port map (
            O => \N__54062\,
            I => \N__54033\
        );

    \I__13299\ : CascadeMux
    port map (
            O => \N__54061\,
            I => \N__54029\
        );

    \I__13298\ : InMux
    port map (
            O => \N__54060\,
            I => \N__54017\
        );

    \I__13297\ : InMux
    port map (
            O => \N__54059\,
            I => \N__54014\
        );

    \I__13296\ : InMux
    port map (
            O => \N__54058\,
            I => \N__54009\
        );

    \I__13295\ : InMux
    port map (
            O => \N__54057\,
            I => \N__54009\
        );

    \I__13294\ : InMux
    port map (
            O => \N__54056\,
            I => \N__54006\
        );

    \I__13293\ : InMux
    port map (
            O => \N__54055\,
            I => \N__54003\
        );

    \I__13292\ : InMux
    port map (
            O => \N__54054\,
            I => \N__53987\
        );

    \I__13291\ : InMux
    port map (
            O => \N__54053\,
            I => \N__53987\
        );

    \I__13290\ : InMux
    port map (
            O => \N__54052\,
            I => \N__53987\
        );

    \I__13289\ : InMux
    port map (
            O => \N__54051\,
            I => \N__53987\
        );

    \I__13288\ : InMux
    port map (
            O => \N__54050\,
            I => \N__53980\
        );

    \I__13287\ : InMux
    port map (
            O => \N__54049\,
            I => \N__53980\
        );

    \I__13286\ : CascadeMux
    port map (
            O => \N__54048\,
            I => \N__53977\
        );

    \I__13285\ : CascadeMux
    port map (
            O => \N__54047\,
            I => \N__53952\
        );

    \I__13284\ : LocalMux
    port map (
            O => \N__54042\,
            I => \N__53942\
        );

    \I__13283\ : InMux
    port map (
            O => \N__54041\,
            I => \N__53939\
        );

    \I__13282\ : InMux
    port map (
            O => \N__54040\,
            I => \N__53930\
        );

    \I__13281\ : InMux
    port map (
            O => \N__54039\,
            I => \N__53930\
        );

    \I__13280\ : InMux
    port map (
            O => \N__54038\,
            I => \N__53930\
        );

    \I__13279\ : InMux
    port map (
            O => \N__54037\,
            I => \N__53930\
        );

    \I__13278\ : InMux
    port map (
            O => \N__54036\,
            I => \N__53920\
        );

    \I__13277\ : LocalMux
    port map (
            O => \N__54033\,
            I => \N__53917\
        );

    \I__13276\ : InMux
    port map (
            O => \N__54032\,
            I => \N__53914\
        );

    \I__13275\ : InMux
    port map (
            O => \N__54029\,
            I => \N__53908\
        );

    \I__13274\ : InMux
    port map (
            O => \N__54028\,
            I => \N__53901\
        );

    \I__13273\ : InMux
    port map (
            O => \N__54027\,
            I => \N__53901\
        );

    \I__13272\ : InMux
    port map (
            O => \N__54026\,
            I => \N__53901\
        );

    \I__13271\ : InMux
    port map (
            O => \N__54025\,
            I => \N__53890\
        );

    \I__13270\ : InMux
    port map (
            O => \N__54024\,
            I => \N__53887\
        );

    \I__13269\ : InMux
    port map (
            O => \N__54023\,
            I => \N__53880\
        );

    \I__13268\ : InMux
    port map (
            O => \N__54022\,
            I => \N__53880\
        );

    \I__13267\ : InMux
    port map (
            O => \N__54021\,
            I => \N__53875\
        );

    \I__13266\ : InMux
    port map (
            O => \N__54020\,
            I => \N__53875\
        );

    \I__13265\ : LocalMux
    port map (
            O => \N__54017\,
            I => \N__53864\
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__54014\,
            I => \N__53864\
        );

    \I__13263\ : LocalMux
    port map (
            O => \N__54009\,
            I => \N__53864\
        );

    \I__13262\ : LocalMux
    port map (
            O => \N__54006\,
            I => \N__53861\
        );

    \I__13261\ : LocalMux
    port map (
            O => \N__54003\,
            I => \N__53858\
        );

    \I__13260\ : InMux
    port map (
            O => \N__54002\,
            I => \N__53853\
        );

    \I__13259\ : InMux
    port map (
            O => \N__54001\,
            I => \N__53848\
        );

    \I__13258\ : InMux
    port map (
            O => \N__54000\,
            I => \N__53848\
        );

    \I__13257\ : InMux
    port map (
            O => \N__53999\,
            I => \N__53843\
        );

    \I__13256\ : InMux
    port map (
            O => \N__53998\,
            I => \N__53843\
        );

    \I__13255\ : InMux
    port map (
            O => \N__53997\,
            I => \N__53838\
        );

    \I__13254\ : InMux
    port map (
            O => \N__53996\,
            I => \N__53838\
        );

    \I__13253\ : LocalMux
    port map (
            O => \N__53987\,
            I => \N__53835\
        );

    \I__13252\ : InMux
    port map (
            O => \N__53986\,
            I => \N__53832\
        );

    \I__13251\ : InMux
    port map (
            O => \N__53985\,
            I => \N__53829\
        );

    \I__13250\ : LocalMux
    port map (
            O => \N__53980\,
            I => \N__53826\
        );

    \I__13249\ : InMux
    port map (
            O => \N__53977\,
            I => \N__53823\
        );

    \I__13248\ : InMux
    port map (
            O => \N__53976\,
            I => \N__53816\
        );

    \I__13247\ : InMux
    port map (
            O => \N__53975\,
            I => \N__53816\
        );

    \I__13246\ : InMux
    port map (
            O => \N__53974\,
            I => \N__53816\
        );

    \I__13245\ : InMux
    port map (
            O => \N__53973\,
            I => \N__53813\
        );

    \I__13244\ : InMux
    port map (
            O => \N__53972\,
            I => \N__53808\
        );

    \I__13243\ : InMux
    port map (
            O => \N__53971\,
            I => \N__53799\
        );

    \I__13242\ : InMux
    port map (
            O => \N__53970\,
            I => \N__53799\
        );

    \I__13241\ : InMux
    port map (
            O => \N__53969\,
            I => \N__53792\
        );

    \I__13240\ : InMux
    port map (
            O => \N__53968\,
            I => \N__53792\
        );

    \I__13239\ : InMux
    port map (
            O => \N__53967\,
            I => \N__53792\
        );

    \I__13238\ : InMux
    port map (
            O => \N__53966\,
            I => \N__53783\
        );

    \I__13237\ : InMux
    port map (
            O => \N__53965\,
            I => \N__53783\
        );

    \I__13236\ : InMux
    port map (
            O => \N__53964\,
            I => \N__53783\
        );

    \I__13235\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53783\
        );

    \I__13234\ : InMux
    port map (
            O => \N__53962\,
            I => \N__53771\
        );

    \I__13233\ : InMux
    port map (
            O => \N__53961\,
            I => \N__53771\
        );

    \I__13232\ : InMux
    port map (
            O => \N__53960\,
            I => \N__53771\
        );

    \I__13231\ : InMux
    port map (
            O => \N__53959\,
            I => \N__53766\
        );

    \I__13230\ : InMux
    port map (
            O => \N__53958\,
            I => \N__53766\
        );

    \I__13229\ : InMux
    port map (
            O => \N__53957\,
            I => \N__53763\
        );

    \I__13228\ : InMux
    port map (
            O => \N__53956\,
            I => \N__53760\
        );

    \I__13227\ : InMux
    port map (
            O => \N__53955\,
            I => \N__53754\
        );

    \I__13226\ : InMux
    port map (
            O => \N__53952\,
            I => \N__53748\
        );

    \I__13225\ : InMux
    port map (
            O => \N__53951\,
            I => \N__53748\
        );

    \I__13224\ : InMux
    port map (
            O => \N__53950\,
            I => \N__53743\
        );

    \I__13223\ : InMux
    port map (
            O => \N__53949\,
            I => \N__53743\
        );

    \I__13222\ : InMux
    port map (
            O => \N__53948\,
            I => \N__53735\
        );

    \I__13221\ : InMux
    port map (
            O => \N__53947\,
            I => \N__53735\
        );

    \I__13220\ : InMux
    port map (
            O => \N__53946\,
            I => \N__53735\
        );

    \I__13219\ : InMux
    port map (
            O => \N__53945\,
            I => \N__53732\
        );

    \I__13218\ : Span4Mux_s2_v
    port map (
            O => \N__53942\,
            I => \N__53725\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__53939\,
            I => \N__53725\
        );

    \I__13216\ : LocalMux
    port map (
            O => \N__53930\,
            I => \N__53725\
        );

    \I__13215\ : InMux
    port map (
            O => \N__53929\,
            I => \N__53718\
        );

    \I__13214\ : InMux
    port map (
            O => \N__53928\,
            I => \N__53718\
        );

    \I__13213\ : InMux
    port map (
            O => \N__53927\,
            I => \N__53718\
        );

    \I__13212\ : InMux
    port map (
            O => \N__53926\,
            I => \N__53709\
        );

    \I__13211\ : InMux
    port map (
            O => \N__53925\,
            I => \N__53709\
        );

    \I__13210\ : InMux
    port map (
            O => \N__53924\,
            I => \N__53709\
        );

    \I__13209\ : InMux
    port map (
            O => \N__53923\,
            I => \N__53709\
        );

    \I__13208\ : LocalMux
    port map (
            O => \N__53920\,
            I => \N__53702\
        );

    \I__13207\ : Span4Mux_v
    port map (
            O => \N__53917\,
            I => \N__53702\
        );

    \I__13206\ : LocalMux
    port map (
            O => \N__53914\,
            I => \N__53702\
        );

    \I__13205\ : InMux
    port map (
            O => \N__53913\,
            I => \N__53695\
        );

    \I__13204\ : InMux
    port map (
            O => \N__53912\,
            I => \N__53695\
        );

    \I__13203\ : InMux
    port map (
            O => \N__53911\,
            I => \N__53695\
        );

    \I__13202\ : LocalMux
    port map (
            O => \N__53908\,
            I => \N__53690\
        );

    \I__13201\ : LocalMux
    port map (
            O => \N__53901\,
            I => \N__53690\
        );

    \I__13200\ : InMux
    port map (
            O => \N__53900\,
            I => \N__53687\
        );

    \I__13199\ : CascadeMux
    port map (
            O => \N__53899\,
            I => \N__53682\
        );

    \I__13198\ : InMux
    port map (
            O => \N__53898\,
            I => \N__53677\
        );

    \I__13197\ : InMux
    port map (
            O => \N__53897\,
            I => \N__53672\
        );

    \I__13196\ : InMux
    port map (
            O => \N__53896\,
            I => \N__53669\
        );

    \I__13195\ : InMux
    port map (
            O => \N__53895\,
            I => \N__53662\
        );

    \I__13194\ : InMux
    port map (
            O => \N__53894\,
            I => \N__53662\
        );

    \I__13193\ : InMux
    port map (
            O => \N__53893\,
            I => \N__53662\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__53890\,
            I => \N__53657\
        );

    \I__13191\ : LocalMux
    port map (
            O => \N__53887\,
            I => \N__53657\
        );

    \I__13190\ : InMux
    port map (
            O => \N__53886\,
            I => \N__53652\
        );

    \I__13189\ : InMux
    port map (
            O => \N__53885\,
            I => \N__53652\
        );

    \I__13188\ : LocalMux
    port map (
            O => \N__53880\,
            I => \N__53647\
        );

    \I__13187\ : LocalMux
    port map (
            O => \N__53875\,
            I => \N__53647\
        );

    \I__13186\ : InMux
    port map (
            O => \N__53874\,
            I => \N__53641\
        );

    \I__13185\ : InMux
    port map (
            O => \N__53873\,
            I => \N__53636\
        );

    \I__13184\ : InMux
    port map (
            O => \N__53872\,
            I => \N__53636\
        );

    \I__13183\ : InMux
    port map (
            O => \N__53871\,
            I => \N__53633\
        );

    \I__13182\ : Span4Mux_v
    port map (
            O => \N__53864\,
            I => \N__53630\
        );

    \I__13181\ : Span4Mux_s3_v
    port map (
            O => \N__53861\,
            I => \N__53625\
        );

    \I__13180\ : Span4Mux_h
    port map (
            O => \N__53858\,
            I => \N__53625\
        );

    \I__13179\ : InMux
    port map (
            O => \N__53857\,
            I => \N__53620\
        );

    \I__13178\ : InMux
    port map (
            O => \N__53856\,
            I => \N__53620\
        );

    \I__13177\ : LocalMux
    port map (
            O => \N__53853\,
            I => \N__53613\
        );

    \I__13176\ : LocalMux
    port map (
            O => \N__53848\,
            I => \N__53613\
        );

    \I__13175\ : LocalMux
    port map (
            O => \N__53843\,
            I => \N__53613\
        );

    \I__13174\ : LocalMux
    port map (
            O => \N__53838\,
            I => \N__53610\
        );

    \I__13173\ : Span4Mux_h
    port map (
            O => \N__53835\,
            I => \N__53607\
        );

    \I__13172\ : LocalMux
    port map (
            O => \N__53832\,
            I => \N__53594\
        );

    \I__13171\ : LocalMux
    port map (
            O => \N__53829\,
            I => \N__53594\
        );

    \I__13170\ : Span4Mux_h
    port map (
            O => \N__53826\,
            I => \N__53594\
        );

    \I__13169\ : LocalMux
    port map (
            O => \N__53823\,
            I => \N__53594\
        );

    \I__13168\ : LocalMux
    port map (
            O => \N__53816\,
            I => \N__53594\
        );

    \I__13167\ : LocalMux
    port map (
            O => \N__53813\,
            I => \N__53594\
        );

    \I__13166\ : CascadeMux
    port map (
            O => \N__53812\,
            I => \N__53591\
        );

    \I__13165\ : InMux
    port map (
            O => \N__53811\,
            I => \N__53587\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__53808\,
            I => \N__53584\
        );

    \I__13163\ : InMux
    port map (
            O => \N__53807\,
            I => \N__53579\
        );

    \I__13162\ : InMux
    port map (
            O => \N__53806\,
            I => \N__53579\
        );

    \I__13161\ : InMux
    port map (
            O => \N__53805\,
            I => \N__53576\
        );

    \I__13160\ : InMux
    port map (
            O => \N__53804\,
            I => \N__53573\
        );

    \I__13159\ : LocalMux
    port map (
            O => \N__53799\,
            I => \N__53570\
        );

    \I__13158\ : LocalMux
    port map (
            O => \N__53792\,
            I => \N__53565\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__53783\,
            I => \N__53565\
        );

    \I__13156\ : InMux
    port map (
            O => \N__53782\,
            I => \N__53562\
        );

    \I__13155\ : InMux
    port map (
            O => \N__53781\,
            I => \N__53559\
        );

    \I__13154\ : InMux
    port map (
            O => \N__53780\,
            I => \N__53552\
        );

    \I__13153\ : InMux
    port map (
            O => \N__53779\,
            I => \N__53552\
        );

    \I__13152\ : InMux
    port map (
            O => \N__53778\,
            I => \N__53552\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__53771\,
            I => \N__53543\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__53766\,
            I => \N__53543\
        );

    \I__13149\ : LocalMux
    port map (
            O => \N__53763\,
            I => \N__53543\
        );

    \I__13148\ : LocalMux
    port map (
            O => \N__53760\,
            I => \N__53543\
        );

    \I__13147\ : InMux
    port map (
            O => \N__53759\,
            I => \N__53540\
        );

    \I__13146\ : InMux
    port map (
            O => \N__53758\,
            I => \N__53535\
        );

    \I__13145\ : InMux
    port map (
            O => \N__53757\,
            I => \N__53535\
        );

    \I__13144\ : LocalMux
    port map (
            O => \N__53754\,
            I => \N__53532\
        );

    \I__13143\ : InMux
    port map (
            O => \N__53753\,
            I => \N__53529\
        );

    \I__13142\ : LocalMux
    port map (
            O => \N__53748\,
            I => \N__53526\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__53743\,
            I => \N__53523\
        );

    \I__13140\ : InMux
    port map (
            O => \N__53742\,
            I => \N__53520\
        );

    \I__13139\ : LocalMux
    port map (
            O => \N__53735\,
            I => \N__53517\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__53732\,
            I => \N__53513\
        );

    \I__13137\ : Span4Mux_v
    port map (
            O => \N__53725\,
            I => \N__53510\
        );

    \I__13136\ : LocalMux
    port map (
            O => \N__53718\,
            I => \N__53505\
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__53709\,
            I => \N__53505\
        );

    \I__13134\ : Span4Mux_s2_v
    port map (
            O => \N__53702\,
            I => \N__53500\
        );

    \I__13133\ : LocalMux
    port map (
            O => \N__53695\,
            I => \N__53500\
        );

    \I__13132\ : Span4Mux_v
    port map (
            O => \N__53690\,
            I => \N__53495\
        );

    \I__13131\ : LocalMux
    port map (
            O => \N__53687\,
            I => \N__53495\
        );

    \I__13130\ : InMux
    port map (
            O => \N__53686\,
            I => \N__53486\
        );

    \I__13129\ : InMux
    port map (
            O => \N__53685\,
            I => \N__53486\
        );

    \I__13128\ : InMux
    port map (
            O => \N__53682\,
            I => \N__53486\
        );

    \I__13127\ : InMux
    port map (
            O => \N__53681\,
            I => \N__53486\
        );

    \I__13126\ : InMux
    port map (
            O => \N__53680\,
            I => \N__53483\
        );

    \I__13125\ : LocalMux
    port map (
            O => \N__53677\,
            I => \N__53480\
        );

    \I__13124\ : InMux
    port map (
            O => \N__53676\,
            I => \N__53475\
        );

    \I__13123\ : InMux
    port map (
            O => \N__53675\,
            I => \N__53475\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__53672\,
            I => \N__53466\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__53669\,
            I => \N__53466\
        );

    \I__13120\ : LocalMux
    port map (
            O => \N__53662\,
            I => \N__53466\
        );

    \I__13119\ : Span4Mux_v
    port map (
            O => \N__53657\,
            I => \N__53466\
        );

    \I__13118\ : LocalMux
    port map (
            O => \N__53652\,
            I => \N__53461\
        );

    \I__13117\ : Span4Mux_v
    port map (
            O => \N__53647\,
            I => \N__53461\
        );

    \I__13116\ : InMux
    port map (
            O => \N__53646\,
            I => \N__53454\
        );

    \I__13115\ : InMux
    port map (
            O => \N__53645\,
            I => \N__53454\
        );

    \I__13114\ : InMux
    port map (
            O => \N__53644\,
            I => \N__53454\
        );

    \I__13113\ : LocalMux
    port map (
            O => \N__53641\,
            I => \N__53447\
        );

    \I__13112\ : LocalMux
    port map (
            O => \N__53636\,
            I => \N__53447\
        );

    \I__13111\ : LocalMux
    port map (
            O => \N__53633\,
            I => \N__53447\
        );

    \I__13110\ : Span4Mux_h
    port map (
            O => \N__53630\,
            I => \N__53442\
        );

    \I__13109\ : Span4Mux_v
    port map (
            O => \N__53625\,
            I => \N__53442\
        );

    \I__13108\ : LocalMux
    port map (
            O => \N__53620\,
            I => \N__53435\
        );

    \I__13107\ : Span4Mux_h
    port map (
            O => \N__53613\,
            I => \N__53435\
        );

    \I__13106\ : Span4Mux_h
    port map (
            O => \N__53610\,
            I => \N__53435\
        );

    \I__13105\ : Span4Mux_v
    port map (
            O => \N__53607\,
            I => \N__53430\
        );

    \I__13104\ : Span4Mux_v
    port map (
            O => \N__53594\,
            I => \N__53430\
        );

    \I__13103\ : InMux
    port map (
            O => \N__53591\,
            I => \N__53425\
        );

    \I__13102\ : InMux
    port map (
            O => \N__53590\,
            I => \N__53425\
        );

    \I__13101\ : LocalMux
    port map (
            O => \N__53587\,
            I => \N__53422\
        );

    \I__13100\ : Span4Mux_v
    port map (
            O => \N__53584\,
            I => \N__53418\
        );

    \I__13099\ : LocalMux
    port map (
            O => \N__53579\,
            I => \N__53415\
        );

    \I__13098\ : LocalMux
    port map (
            O => \N__53576\,
            I => \N__53412\
        );

    \I__13097\ : LocalMux
    port map (
            O => \N__53573\,
            I => \N__53401\
        );

    \I__13096\ : Span4Mux_h
    port map (
            O => \N__53570\,
            I => \N__53401\
        );

    \I__13095\ : Span4Mux_s2_v
    port map (
            O => \N__53565\,
            I => \N__53401\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__53562\,
            I => \N__53401\
        );

    \I__13093\ : LocalMux
    port map (
            O => \N__53559\,
            I => \N__53401\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__53552\,
            I => \N__53396\
        );

    \I__13091\ : Span4Mux_v
    port map (
            O => \N__53543\,
            I => \N__53396\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__53540\,
            I => \N__53387\
        );

    \I__13089\ : LocalMux
    port map (
            O => \N__53535\,
            I => \N__53387\
        );

    \I__13088\ : Span4Mux_h
    port map (
            O => \N__53532\,
            I => \N__53387\
        );

    \I__13087\ : LocalMux
    port map (
            O => \N__53529\,
            I => \N__53387\
        );

    \I__13086\ : Span4Mux_s2_v
    port map (
            O => \N__53526\,
            I => \N__53380\
        );

    \I__13085\ : Span4Mux_s2_v
    port map (
            O => \N__53523\,
            I => \N__53380\
        );

    \I__13084\ : LocalMux
    port map (
            O => \N__53520\,
            I => \N__53380\
        );

    \I__13083\ : Span4Mux_s2_v
    port map (
            O => \N__53517\,
            I => \N__53377\
        );

    \I__13082\ : InMux
    port map (
            O => \N__53516\,
            I => \N__53374\
        );

    \I__13081\ : Span4Mux_v
    port map (
            O => \N__53513\,
            I => \N__53365\
        );

    \I__13080\ : Span4Mux_h
    port map (
            O => \N__53510\,
            I => \N__53365\
        );

    \I__13079\ : Span4Mux_v
    port map (
            O => \N__53505\,
            I => \N__53365\
        );

    \I__13078\ : Span4Mux_v
    port map (
            O => \N__53500\,
            I => \N__53365\
        );

    \I__13077\ : Span4Mux_h
    port map (
            O => \N__53495\,
            I => \N__53358\
        );

    \I__13076\ : LocalMux
    port map (
            O => \N__53486\,
            I => \N__53358\
        );

    \I__13075\ : LocalMux
    port map (
            O => \N__53483\,
            I => \N__53358\
        );

    \I__13074\ : Span4Mux_h
    port map (
            O => \N__53480\,
            I => \N__53351\
        );

    \I__13073\ : LocalMux
    port map (
            O => \N__53475\,
            I => \N__53351\
        );

    \I__13072\ : Span4Mux_v
    port map (
            O => \N__53466\,
            I => \N__53342\
        );

    \I__13071\ : Span4Mux_h
    port map (
            O => \N__53461\,
            I => \N__53342\
        );

    \I__13070\ : LocalMux
    port map (
            O => \N__53454\,
            I => \N__53342\
        );

    \I__13069\ : Span4Mux_v
    port map (
            O => \N__53447\,
            I => \N__53342\
        );

    \I__13068\ : Span4Mux_h
    port map (
            O => \N__53442\,
            I => \N__53335\
        );

    \I__13067\ : Span4Mux_h
    port map (
            O => \N__53435\,
            I => \N__53335\
        );

    \I__13066\ : Span4Mux_h
    port map (
            O => \N__53430\,
            I => \N__53335\
        );

    \I__13065\ : LocalMux
    port map (
            O => \N__53425\,
            I => \N__53330\
        );

    \I__13064\ : Span4Mux_v
    port map (
            O => \N__53422\,
            I => \N__53330\
        );

    \I__13063\ : InMux
    port map (
            O => \N__53421\,
            I => \N__53327\
        );

    \I__13062\ : Span4Mux_h
    port map (
            O => \N__53418\,
            I => \N__53320\
        );

    \I__13061\ : Span4Mux_v
    port map (
            O => \N__53415\,
            I => \N__53320\
        );

    \I__13060\ : Span4Mux_v
    port map (
            O => \N__53412\,
            I => \N__53320\
        );

    \I__13059\ : Span4Mux_h
    port map (
            O => \N__53401\,
            I => \N__53317\
        );

    \I__13058\ : Span4Mux_h
    port map (
            O => \N__53396\,
            I => \N__53310\
        );

    \I__13057\ : Span4Mux_v
    port map (
            O => \N__53387\,
            I => \N__53310\
        );

    \I__13056\ : Span4Mux_v
    port map (
            O => \N__53380\,
            I => \N__53310\
        );

    \I__13055\ : Span4Mux_h
    port map (
            O => \N__53377\,
            I => \N__53305\
        );

    \I__13054\ : LocalMux
    port map (
            O => \N__53374\,
            I => \N__53305\
        );

    \I__13053\ : Span4Mux_h
    port map (
            O => \N__53365\,
            I => \N__53302\
        );

    \I__13052\ : Span4Mux_v
    port map (
            O => \N__53358\,
            I => \N__53299\
        );

    \I__13051\ : InMux
    port map (
            O => \N__53357\,
            I => \N__53294\
        );

    \I__13050\ : InMux
    port map (
            O => \N__53356\,
            I => \N__53294\
        );

    \I__13049\ : Span4Mux_v
    port map (
            O => \N__53351\,
            I => \N__53289\
        );

    \I__13048\ : Span4Mux_h
    port map (
            O => \N__53342\,
            I => \N__53289\
        );

    \I__13047\ : Span4Mux_v
    port map (
            O => \N__53335\,
            I => \N__53282\
        );

    \I__13046\ : Span4Mux_s3_v
    port map (
            O => \N__53330\,
            I => \N__53282\
        );

    \I__13045\ : LocalMux
    port map (
            O => \N__53327\,
            I => \N__53282\
        );

    \I__13044\ : Span4Mux_h
    port map (
            O => \N__53320\,
            I => \N__53275\
        );

    \I__13043\ : Span4Mux_v
    port map (
            O => \N__53317\,
            I => \N__53275\
        );

    \I__13042\ : Span4Mux_v
    port map (
            O => \N__53310\,
            I => \N__53275\
        );

    \I__13041\ : Span4Mux_v
    port map (
            O => \N__53305\,
            I => \N__53268\
        );

    \I__13040\ : Span4Mux_h
    port map (
            O => \N__53302\,
            I => \N__53268\
        );

    \I__13039\ : Span4Mux_v
    port map (
            O => \N__53299\,
            I => \N__53268\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__53294\,
            I => \paramsZ0Z_0\
        );

    \I__13037\ : Odrv4
    port map (
            O => \N__53289\,
            I => \paramsZ0Z_0\
        );

    \I__13036\ : Odrv4
    port map (
            O => \N__53282\,
            I => \paramsZ0Z_0\
        );

    \I__13035\ : Odrv4
    port map (
            O => \N__53275\,
            I => \paramsZ0Z_0\
        );

    \I__13034\ : Odrv4
    port map (
            O => \N__53268\,
            I => \paramsZ0Z_0\
        );

    \I__13033\ : CascadeMux
    port map (
            O => \N__53257\,
            I => \N__53251\
        );

    \I__13032\ : InMux
    port map (
            O => \N__53256\,
            I => \N__53247\
        );

    \I__13031\ : InMux
    port map (
            O => \N__53255\,
            I => \N__53244\
        );

    \I__13030\ : InMux
    port map (
            O => \N__53254\,
            I => \N__53233\
        );

    \I__13029\ : InMux
    port map (
            O => \N__53251\,
            I => \N__53225\
        );

    \I__13028\ : CascadeMux
    port map (
            O => \N__53250\,
            I => \N__53209\
        );

    \I__13027\ : LocalMux
    port map (
            O => \N__53247\,
            I => \N__53200\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__53244\,
            I => \N__53200\
        );

    \I__13025\ : CascadeMux
    port map (
            O => \N__53243\,
            I => \N__53197\
        );

    \I__13024\ : CascadeMux
    port map (
            O => \N__53242\,
            I => \N__53190\
        );

    \I__13023\ : CascadeMux
    port map (
            O => \N__53241\,
            I => \N__53187\
        );

    \I__13022\ : CascadeMux
    port map (
            O => \N__53240\,
            I => \N__53184\
        );

    \I__13021\ : CascadeMux
    port map (
            O => \N__53239\,
            I => \N__53177\
        );

    \I__13020\ : InMux
    port map (
            O => \N__53238\,
            I => \N__53170\
        );

    \I__13019\ : InMux
    port map (
            O => \N__53237\,
            I => \N__53170\
        );

    \I__13018\ : CascadeMux
    port map (
            O => \N__53236\,
            I => \N__53155\
        );

    \I__13017\ : LocalMux
    port map (
            O => \N__53233\,
            I => \N__53149\
        );

    \I__13016\ : CascadeMux
    port map (
            O => \N__53232\,
            I => \N__53146\
        );

    \I__13015\ : CascadeMux
    port map (
            O => \N__53231\,
            I => \N__53140\
        );

    \I__13014\ : CascadeMux
    port map (
            O => \N__53230\,
            I => \N__53136\
        );

    \I__13013\ : CascadeMux
    port map (
            O => \N__53229\,
            I => \N__53131\
        );

    \I__13012\ : CascadeMux
    port map (
            O => \N__53228\,
            I => \N__53126\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__53225\,
            I => \N__53123\
        );

    \I__13010\ : CascadeMux
    port map (
            O => \N__53224\,
            I => \N__53115\
        );

    \I__13009\ : CascadeMux
    port map (
            O => \N__53223\,
            I => \N__53111\
        );

    \I__13008\ : CascadeMux
    port map (
            O => \N__53222\,
            I => \N__53108\
        );

    \I__13007\ : CascadeMux
    port map (
            O => \N__53221\,
            I => \N__53105\
        );

    \I__13006\ : CascadeMux
    port map (
            O => \N__53220\,
            I => \N__53099\
        );

    \I__13005\ : CascadeMux
    port map (
            O => \N__53219\,
            I => \N__53095\
        );

    \I__13004\ : CascadeMux
    port map (
            O => \N__53218\,
            I => \N__53092\
        );

    \I__13003\ : CascadeMux
    port map (
            O => \N__53217\,
            I => \N__53087\
        );

    \I__13002\ : CascadeMux
    port map (
            O => \N__53216\,
            I => \N__53084\
        );

    \I__13001\ : CascadeMux
    port map (
            O => \N__53215\,
            I => \N__53081\
        );

    \I__13000\ : CascadeMux
    port map (
            O => \N__53214\,
            I => \N__53077\
        );

    \I__12999\ : CascadeMux
    port map (
            O => \N__53213\,
            I => \N__53074\
        );

    \I__12998\ : InMux
    port map (
            O => \N__53212\,
            I => \N__53069\
        );

    \I__12997\ : InMux
    port map (
            O => \N__53209\,
            I => \N__53069\
        );

    \I__12996\ : CascadeMux
    port map (
            O => \N__53208\,
            I => \N__53065\
        );

    \I__12995\ : CascadeMux
    port map (
            O => \N__53207\,
            I => \N__53061\
        );

    \I__12994\ : CascadeMux
    port map (
            O => \N__53206\,
            I => \N__53058\
        );

    \I__12993\ : CascadeMux
    port map (
            O => \N__53205\,
            I => \N__53055\
        );

    \I__12992\ : Span4Mux_h
    port map (
            O => \N__53200\,
            I => \N__53052\
        );

    \I__12991\ : InMux
    port map (
            O => \N__53197\,
            I => \N__53045\
        );

    \I__12990\ : InMux
    port map (
            O => \N__53196\,
            I => \N__53045\
        );

    \I__12989\ : InMux
    port map (
            O => \N__53195\,
            I => \N__53045\
        );

    \I__12988\ : InMux
    port map (
            O => \N__53194\,
            I => \N__53034\
        );

    \I__12987\ : InMux
    port map (
            O => \N__53193\,
            I => \N__53034\
        );

    \I__12986\ : InMux
    port map (
            O => \N__53190\,
            I => \N__53034\
        );

    \I__12985\ : InMux
    port map (
            O => \N__53187\,
            I => \N__53034\
        );

    \I__12984\ : InMux
    port map (
            O => \N__53184\,
            I => \N__53034\
        );

    \I__12983\ : CascadeMux
    port map (
            O => \N__53183\,
            I => \N__53031\
        );

    \I__12982\ : CascadeMux
    port map (
            O => \N__53182\,
            I => \N__53028\
        );

    \I__12981\ : CascadeMux
    port map (
            O => \N__53181\,
            I => \N__53025\
        );

    \I__12980\ : InMux
    port map (
            O => \N__53180\,
            I => \N__53018\
        );

    \I__12979\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53018\
        );

    \I__12978\ : InMux
    port map (
            O => \N__53176\,
            I => \N__53018\
        );

    \I__12977\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53015\
        );

    \I__12976\ : LocalMux
    port map (
            O => \N__53170\,
            I => \N__53011\
        );

    \I__12975\ : CascadeMux
    port map (
            O => \N__53169\,
            I => \N__53008\
        );

    \I__12974\ : CascadeMux
    port map (
            O => \N__53168\,
            I => \N__53005\
        );

    \I__12973\ : CascadeMux
    port map (
            O => \N__53167\,
            I => \N__53000\
        );

    \I__12972\ : CascadeMux
    port map (
            O => \N__53166\,
            I => \N__52997\
        );

    \I__12971\ : CascadeMux
    port map (
            O => \N__53165\,
            I => \N__52993\
        );

    \I__12970\ : CascadeMux
    port map (
            O => \N__53164\,
            I => \N__52989\
        );

    \I__12969\ : CascadeMux
    port map (
            O => \N__53163\,
            I => \N__52986\
        );

    \I__12968\ : CascadeMux
    port map (
            O => \N__53162\,
            I => \N__52979\
        );

    \I__12967\ : CascadeMux
    port map (
            O => \N__53161\,
            I => \N__52976\
        );

    \I__12966\ : CascadeMux
    port map (
            O => \N__53160\,
            I => \N__52973\
        );

    \I__12965\ : InMux
    port map (
            O => \N__53159\,
            I => \N__52967\
        );

    \I__12964\ : CascadeMux
    port map (
            O => \N__53158\,
            I => \N__52964\
        );

    \I__12963\ : InMux
    port map (
            O => \N__53155\,
            I => \N__52960\
        );

    \I__12962\ : CascadeMux
    port map (
            O => \N__53154\,
            I => \N__52957\
        );

    \I__12961\ : CascadeMux
    port map (
            O => \N__53153\,
            I => \N__52954\
        );

    \I__12960\ : CascadeMux
    port map (
            O => \N__53152\,
            I => \N__52951\
        );

    \I__12959\ : Span4Mux_s3_h
    port map (
            O => \N__53149\,
            I => \N__52948\
        );

    \I__12958\ : InMux
    port map (
            O => \N__53146\,
            I => \N__52945\
        );

    \I__12957\ : InMux
    port map (
            O => \N__53145\,
            I => \N__52942\
        );

    \I__12956\ : CascadeMux
    port map (
            O => \N__53144\,
            I => \N__52934\
        );

    \I__12955\ : CascadeMux
    port map (
            O => \N__53143\,
            I => \N__52931\
        );

    \I__12954\ : InMux
    port map (
            O => \N__53140\,
            I => \N__52928\
        );

    \I__12953\ : InMux
    port map (
            O => \N__53139\,
            I => \N__52925\
        );

    \I__12952\ : InMux
    port map (
            O => \N__53136\,
            I => \N__52922\
        );

    \I__12951\ : InMux
    port map (
            O => \N__53135\,
            I => \N__52915\
        );

    \I__12950\ : InMux
    port map (
            O => \N__53134\,
            I => \N__52915\
        );

    \I__12949\ : InMux
    port map (
            O => \N__53131\,
            I => \N__52915\
        );

    \I__12948\ : CascadeMux
    port map (
            O => \N__53130\,
            I => \N__52912\
        );

    \I__12947\ : CascadeMux
    port map (
            O => \N__53129\,
            I => \N__52909\
        );

    \I__12946\ : InMux
    port map (
            O => \N__53126\,
            I => \N__52906\
        );

    \I__12945\ : Span4Mux_s2_v
    port map (
            O => \N__53123\,
            I => \N__52903\
        );

    \I__12944\ : CascadeMux
    port map (
            O => \N__53122\,
            I => \N__52900\
        );

    \I__12943\ : CascadeMux
    port map (
            O => \N__53121\,
            I => \N__52897\
        );

    \I__12942\ : CascadeMux
    port map (
            O => \N__53120\,
            I => \N__52894\
        );

    \I__12941\ : InMux
    port map (
            O => \N__53119\,
            I => \N__52890\
        );

    \I__12940\ : InMux
    port map (
            O => \N__53118\,
            I => \N__52887\
        );

    \I__12939\ : InMux
    port map (
            O => \N__53115\,
            I => \N__52884\
        );

    \I__12938\ : CascadeMux
    port map (
            O => \N__53114\,
            I => \N__52881\
        );

    \I__12937\ : InMux
    port map (
            O => \N__53111\,
            I => \N__52876\
        );

    \I__12936\ : InMux
    port map (
            O => \N__53108\,
            I => \N__52873\
        );

    \I__12935\ : InMux
    port map (
            O => \N__53105\,
            I => \N__52870\
        );

    \I__12934\ : CascadeMux
    port map (
            O => \N__53104\,
            I => \N__52867\
        );

    \I__12933\ : CascadeMux
    port map (
            O => \N__53103\,
            I => \N__52864\
        );

    \I__12932\ : CascadeMux
    port map (
            O => \N__53102\,
            I => \N__52861\
        );

    \I__12931\ : InMux
    port map (
            O => \N__53099\,
            I => \N__52858\
        );

    \I__12930\ : InMux
    port map (
            O => \N__53098\,
            I => \N__52855\
        );

    \I__12929\ : InMux
    port map (
            O => \N__53095\,
            I => \N__52848\
        );

    \I__12928\ : InMux
    port map (
            O => \N__53092\,
            I => \N__52848\
        );

    \I__12927\ : InMux
    port map (
            O => \N__53091\,
            I => \N__52848\
        );

    \I__12926\ : InMux
    port map (
            O => \N__53090\,
            I => \N__52841\
        );

    \I__12925\ : InMux
    port map (
            O => \N__53087\,
            I => \N__52841\
        );

    \I__12924\ : InMux
    port map (
            O => \N__53084\,
            I => \N__52841\
        );

    \I__12923\ : InMux
    port map (
            O => \N__53081\,
            I => \N__52838\
        );

    \I__12922\ : InMux
    port map (
            O => \N__53080\,
            I => \N__52833\
        );

    \I__12921\ : InMux
    port map (
            O => \N__53077\,
            I => \N__52833\
        );

    \I__12920\ : InMux
    port map (
            O => \N__53074\,
            I => \N__52830\
        );

    \I__12919\ : LocalMux
    port map (
            O => \N__53069\,
            I => \N__52827\
        );

    \I__12918\ : CascadeMux
    port map (
            O => \N__53068\,
            I => \N__52824\
        );

    \I__12917\ : InMux
    port map (
            O => \N__53065\,
            I => \N__52821\
        );

    \I__12916\ : InMux
    port map (
            O => \N__53064\,
            I => \N__52816\
        );

    \I__12915\ : InMux
    port map (
            O => \N__53061\,
            I => \N__52811\
        );

    \I__12914\ : InMux
    port map (
            O => \N__53058\,
            I => \N__52811\
        );

    \I__12913\ : InMux
    port map (
            O => \N__53055\,
            I => \N__52808\
        );

    \I__12912\ : Span4Mux_h
    port map (
            O => \N__53052\,
            I => \N__52803\
        );

    \I__12911\ : LocalMux
    port map (
            O => \N__53045\,
            I => \N__52803\
        );

    \I__12910\ : LocalMux
    port map (
            O => \N__53034\,
            I => \N__52800\
        );

    \I__12909\ : InMux
    port map (
            O => \N__53031\,
            I => \N__52793\
        );

    \I__12908\ : InMux
    port map (
            O => \N__53028\,
            I => \N__52793\
        );

    \I__12907\ : InMux
    port map (
            O => \N__53025\,
            I => \N__52793\
        );

    \I__12906\ : LocalMux
    port map (
            O => \N__53018\,
            I => \N__52788\
        );

    \I__12905\ : LocalMux
    port map (
            O => \N__53015\,
            I => \N__52788\
        );

    \I__12904\ : InMux
    port map (
            O => \N__53014\,
            I => \N__52785\
        );

    \I__12903\ : Span4Mux_s2_h
    port map (
            O => \N__53011\,
            I => \N__52782\
        );

    \I__12902\ : InMux
    port map (
            O => \N__53008\,
            I => \N__52775\
        );

    \I__12901\ : InMux
    port map (
            O => \N__53005\,
            I => \N__52775\
        );

    \I__12900\ : InMux
    port map (
            O => \N__53004\,
            I => \N__52775\
        );

    \I__12899\ : InMux
    port map (
            O => \N__53003\,
            I => \N__52766\
        );

    \I__12898\ : InMux
    port map (
            O => \N__53000\,
            I => \N__52766\
        );

    \I__12897\ : InMux
    port map (
            O => \N__52997\,
            I => \N__52766\
        );

    \I__12896\ : InMux
    port map (
            O => \N__52996\,
            I => \N__52766\
        );

    \I__12895\ : InMux
    port map (
            O => \N__52993\,
            I => \N__52759\
        );

    \I__12894\ : InMux
    port map (
            O => \N__52992\,
            I => \N__52759\
        );

    \I__12893\ : InMux
    port map (
            O => \N__52989\,
            I => \N__52759\
        );

    \I__12892\ : InMux
    port map (
            O => \N__52986\,
            I => \N__52742\
        );

    \I__12891\ : InMux
    port map (
            O => \N__52985\,
            I => \N__52742\
        );

    \I__12890\ : InMux
    port map (
            O => \N__52984\,
            I => \N__52742\
        );

    \I__12889\ : InMux
    port map (
            O => \N__52983\,
            I => \N__52742\
        );

    \I__12888\ : InMux
    port map (
            O => \N__52982\,
            I => \N__52742\
        );

    \I__12887\ : InMux
    port map (
            O => \N__52979\,
            I => \N__52742\
        );

    \I__12886\ : InMux
    port map (
            O => \N__52976\,
            I => \N__52742\
        );

    \I__12885\ : InMux
    port map (
            O => \N__52973\,
            I => \N__52742\
        );

    \I__12884\ : CascadeMux
    port map (
            O => \N__52972\,
            I => \N__52738\
        );

    \I__12883\ : CascadeMux
    port map (
            O => \N__52971\,
            I => \N__52735\
        );

    \I__12882\ : CascadeMux
    port map (
            O => \N__52970\,
            I => \N__52732\
        );

    \I__12881\ : LocalMux
    port map (
            O => \N__52967\,
            I => \N__52729\
        );

    \I__12880\ : InMux
    port map (
            O => \N__52964\,
            I => \N__52726\
        );

    \I__12879\ : CascadeMux
    port map (
            O => \N__52963\,
            I => \N__52723\
        );

    \I__12878\ : LocalMux
    port map (
            O => \N__52960\,
            I => \N__52720\
        );

    \I__12877\ : InMux
    port map (
            O => \N__52957\,
            I => \N__52713\
        );

    \I__12876\ : InMux
    port map (
            O => \N__52954\,
            I => \N__52713\
        );

    \I__12875\ : InMux
    port map (
            O => \N__52951\,
            I => \N__52710\
        );

    \I__12874\ : Span4Mux_v
    port map (
            O => \N__52948\,
            I => \N__52703\
        );

    \I__12873\ : LocalMux
    port map (
            O => \N__52945\,
            I => \N__52703\
        );

    \I__12872\ : LocalMux
    port map (
            O => \N__52942\,
            I => \N__52703\
        );

    \I__12871\ : CascadeMux
    port map (
            O => \N__52941\,
            I => \N__52700\
        );

    \I__12870\ : CascadeMux
    port map (
            O => \N__52940\,
            I => \N__52697\
        );

    \I__12869\ : CascadeMux
    port map (
            O => \N__52939\,
            I => \N__52694\
        );

    \I__12868\ : CascadeMux
    port map (
            O => \N__52938\,
            I => \N__52691\
        );

    \I__12867\ : InMux
    port map (
            O => \N__52937\,
            I => \N__52688\
        );

    \I__12866\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52683\
        );

    \I__12865\ : InMux
    port map (
            O => \N__52931\,
            I => \N__52683\
        );

    \I__12864\ : LocalMux
    port map (
            O => \N__52928\,
            I => \N__52674\
        );

    \I__12863\ : LocalMux
    port map (
            O => \N__52925\,
            I => \N__52674\
        );

    \I__12862\ : LocalMux
    port map (
            O => \N__52922\,
            I => \N__52674\
        );

    \I__12861\ : LocalMux
    port map (
            O => \N__52915\,
            I => \N__52674\
        );

    \I__12860\ : InMux
    port map (
            O => \N__52912\,
            I => \N__52669\
        );

    \I__12859\ : InMux
    port map (
            O => \N__52909\,
            I => \N__52669\
        );

    \I__12858\ : LocalMux
    port map (
            O => \N__52906\,
            I => \N__52664\
        );

    \I__12857\ : Span4Mux_h
    port map (
            O => \N__52903\,
            I => \N__52664\
        );

    \I__12856\ : InMux
    port map (
            O => \N__52900\,
            I => \N__52657\
        );

    \I__12855\ : InMux
    port map (
            O => \N__52897\,
            I => \N__52657\
        );

    \I__12854\ : InMux
    port map (
            O => \N__52894\,
            I => \N__52657\
        );

    \I__12853\ : InMux
    port map (
            O => \N__52893\,
            I => \N__52654\
        );

    \I__12852\ : LocalMux
    port map (
            O => \N__52890\,
            I => \N__52647\
        );

    \I__12851\ : LocalMux
    port map (
            O => \N__52887\,
            I => \N__52647\
        );

    \I__12850\ : LocalMux
    port map (
            O => \N__52884\,
            I => \N__52647\
        );

    \I__12849\ : InMux
    port map (
            O => \N__52881\,
            I => \N__52640\
        );

    \I__12848\ : InMux
    port map (
            O => \N__52880\,
            I => \N__52640\
        );

    \I__12847\ : InMux
    port map (
            O => \N__52879\,
            I => \N__52640\
        );

    \I__12846\ : LocalMux
    port map (
            O => \N__52876\,
            I => \N__52633\
        );

    \I__12845\ : LocalMux
    port map (
            O => \N__52873\,
            I => \N__52633\
        );

    \I__12844\ : LocalMux
    port map (
            O => \N__52870\,
            I => \N__52633\
        );

    \I__12843\ : InMux
    port map (
            O => \N__52867\,
            I => \N__52630\
        );

    \I__12842\ : InMux
    port map (
            O => \N__52864\,
            I => \N__52625\
        );

    \I__12841\ : InMux
    port map (
            O => \N__52861\,
            I => \N__52625\
        );

    \I__12840\ : LocalMux
    port map (
            O => \N__52858\,
            I => \N__52620\
        );

    \I__12839\ : LocalMux
    port map (
            O => \N__52855\,
            I => \N__52620\
        );

    \I__12838\ : LocalMux
    port map (
            O => \N__52848\,
            I => \N__52617\
        );

    \I__12837\ : LocalMux
    port map (
            O => \N__52841\,
            I => \N__52610\
        );

    \I__12836\ : LocalMux
    port map (
            O => \N__52838\,
            I => \N__52610\
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__52833\,
            I => \N__52610\
        );

    \I__12834\ : LocalMux
    port map (
            O => \N__52830\,
            I => \N__52605\
        );

    \I__12833\ : Span4Mux_s2_v
    port map (
            O => \N__52827\,
            I => \N__52605\
        );

    \I__12832\ : InMux
    port map (
            O => \N__52824\,
            I => \N__52602\
        );

    \I__12831\ : LocalMux
    port map (
            O => \N__52821\,
            I => \N__52599\
        );

    \I__12830\ : InMux
    port map (
            O => \N__52820\,
            I => \N__52593\
        );

    \I__12829\ : InMux
    port map (
            O => \N__52819\,
            I => \N__52593\
        );

    \I__12828\ : LocalMux
    port map (
            O => \N__52816\,
            I => \N__52586\
        );

    \I__12827\ : LocalMux
    port map (
            O => \N__52811\,
            I => \N__52586\
        );

    \I__12826\ : LocalMux
    port map (
            O => \N__52808\,
            I => \N__52586\
        );

    \I__12825\ : Span4Mux_v
    port map (
            O => \N__52803\,
            I => \N__52581\
        );

    \I__12824\ : Span4Mux_v
    port map (
            O => \N__52800\,
            I => \N__52581\
        );

    \I__12823\ : LocalMux
    port map (
            O => \N__52793\,
            I => \N__52574\
        );

    \I__12822\ : Span4Mux_v
    port map (
            O => \N__52788\,
            I => \N__52574\
        );

    \I__12821\ : LocalMux
    port map (
            O => \N__52785\,
            I => \N__52574\
        );

    \I__12820\ : Span4Mux_v
    port map (
            O => \N__52782\,
            I => \N__52567\
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__52775\,
            I => \N__52567\
        );

    \I__12818\ : LocalMux
    port map (
            O => \N__52766\,
            I => \N__52567\
        );

    \I__12817\ : LocalMux
    port map (
            O => \N__52759\,
            I => \N__52564\
        );

    \I__12816\ : LocalMux
    port map (
            O => \N__52742\,
            I => \N__52561\
        );

    \I__12815\ : InMux
    port map (
            O => \N__52741\,
            I => \N__52558\
        );

    \I__12814\ : InMux
    port map (
            O => \N__52738\,
            I => \N__52555\
        );

    \I__12813\ : InMux
    port map (
            O => \N__52735\,
            I => \N__52550\
        );

    \I__12812\ : InMux
    port map (
            O => \N__52732\,
            I => \N__52550\
        );

    \I__12811\ : Span4Mux_s3_v
    port map (
            O => \N__52729\,
            I => \N__52545\
        );

    \I__12810\ : LocalMux
    port map (
            O => \N__52726\,
            I => \N__52545\
        );

    \I__12809\ : InMux
    port map (
            O => \N__52723\,
            I => \N__52541\
        );

    \I__12808\ : Span4Mux_h
    port map (
            O => \N__52720\,
            I => \N__52538\
        );

    \I__12807\ : InMux
    port map (
            O => \N__52719\,
            I => \N__52534\
        );

    \I__12806\ : InMux
    port map (
            O => \N__52718\,
            I => \N__52531\
        );

    \I__12805\ : LocalMux
    port map (
            O => \N__52713\,
            I => \N__52526\
        );

    \I__12804\ : LocalMux
    port map (
            O => \N__52710\,
            I => \N__52526\
        );

    \I__12803\ : Span4Mux_v
    port map (
            O => \N__52703\,
            I => \N__52523\
        );

    \I__12802\ : InMux
    port map (
            O => \N__52700\,
            I => \N__52520\
        );

    \I__12801\ : InMux
    port map (
            O => \N__52697\,
            I => \N__52517\
        );

    \I__12800\ : InMux
    port map (
            O => \N__52694\,
            I => \N__52512\
        );

    \I__12799\ : InMux
    port map (
            O => \N__52691\,
            I => \N__52512\
        );

    \I__12798\ : LocalMux
    port map (
            O => \N__52688\,
            I => \N__52509\
        );

    \I__12797\ : LocalMux
    port map (
            O => \N__52683\,
            I => \N__52498\
        );

    \I__12796\ : Span4Mux_s2_v
    port map (
            O => \N__52674\,
            I => \N__52498\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__52669\,
            I => \N__52498\
        );

    \I__12794\ : Span4Mux_h
    port map (
            O => \N__52664\,
            I => \N__52498\
        );

    \I__12793\ : LocalMux
    port map (
            O => \N__52657\,
            I => \N__52498\
        );

    \I__12792\ : LocalMux
    port map (
            O => \N__52654\,
            I => \N__52491\
        );

    \I__12791\ : Span4Mux_v
    port map (
            O => \N__52647\,
            I => \N__52491\
        );

    \I__12790\ : LocalMux
    port map (
            O => \N__52640\,
            I => \N__52491\
        );

    \I__12789\ : Span4Mux_v
    port map (
            O => \N__52633\,
            I => \N__52486\
        );

    \I__12788\ : LocalMux
    port map (
            O => \N__52630\,
            I => \N__52486\
        );

    \I__12787\ : LocalMux
    port map (
            O => \N__52625\,
            I => \N__52483\
        );

    \I__12786\ : Span4Mux_v
    port map (
            O => \N__52620\,
            I => \N__52474\
        );

    \I__12785\ : Span4Mux_s2_v
    port map (
            O => \N__52617\,
            I => \N__52474\
        );

    \I__12784\ : Span4Mux_s2_v
    port map (
            O => \N__52610\,
            I => \N__52474\
        );

    \I__12783\ : Span4Mux_h
    port map (
            O => \N__52605\,
            I => \N__52474\
        );

    \I__12782\ : LocalMux
    port map (
            O => \N__52602\,
            I => \N__52469\
        );

    \I__12781\ : Sp12to4
    port map (
            O => \N__52599\,
            I => \N__52469\
        );

    \I__12780\ : CascadeMux
    port map (
            O => \N__52598\,
            I => \N__52466\
        );

    \I__12779\ : LocalMux
    port map (
            O => \N__52593\,
            I => \N__52463\
        );

    \I__12778\ : Span4Mux_v
    port map (
            O => \N__52586\,
            I => \N__52456\
        );

    \I__12777\ : Span4Mux_h
    port map (
            O => \N__52581\,
            I => \N__52456\
        );

    \I__12776\ : Span4Mux_v
    port map (
            O => \N__52574\,
            I => \N__52456\
        );

    \I__12775\ : Span4Mux_h
    port map (
            O => \N__52567\,
            I => \N__52449\
        );

    \I__12774\ : Span4Mux_v
    port map (
            O => \N__52564\,
            I => \N__52449\
        );

    \I__12773\ : Span4Mux_v
    port map (
            O => \N__52561\,
            I => \N__52449\
        );

    \I__12772\ : LocalMux
    port map (
            O => \N__52558\,
            I => \N__52444\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__52555\,
            I => \N__52437\
        );

    \I__12770\ : LocalMux
    port map (
            O => \N__52550\,
            I => \N__52437\
        );

    \I__12769\ : Span4Mux_h
    port map (
            O => \N__52545\,
            I => \N__52437\
        );

    \I__12768\ : InMux
    port map (
            O => \N__52544\,
            I => \N__52434\
        );

    \I__12767\ : LocalMux
    port map (
            O => \N__52541\,
            I => \N__52429\
        );

    \I__12766\ : Sp12to4
    port map (
            O => \N__52538\,
            I => \N__52429\
        );

    \I__12765\ : InMux
    port map (
            O => \N__52537\,
            I => \N__52426\
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__52534\,
            I => \N__52419\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__52531\,
            I => \N__52419\
        );

    \I__12762\ : Sp12to4
    port map (
            O => \N__52526\,
            I => \N__52419\
        );

    \I__12761\ : Sp12to4
    port map (
            O => \N__52523\,
            I => \N__52416\
        );

    \I__12760\ : LocalMux
    port map (
            O => \N__52520\,
            I => \N__52401\
        );

    \I__12759\ : LocalMux
    port map (
            O => \N__52517\,
            I => \N__52401\
        );

    \I__12758\ : LocalMux
    port map (
            O => \N__52512\,
            I => \N__52401\
        );

    \I__12757\ : Span4Mux_v
    port map (
            O => \N__52509\,
            I => \N__52401\
        );

    \I__12756\ : Span4Mux_v
    port map (
            O => \N__52498\,
            I => \N__52401\
        );

    \I__12755\ : Span4Mux_v
    port map (
            O => \N__52491\,
            I => \N__52401\
        );

    \I__12754\ : Span4Mux_h
    port map (
            O => \N__52486\,
            I => \N__52401\
        );

    \I__12753\ : Span4Mux_v
    port map (
            O => \N__52483\,
            I => \N__52396\
        );

    \I__12752\ : Span4Mux_h
    port map (
            O => \N__52474\,
            I => \N__52396\
        );

    \I__12751\ : Span12Mux_s7_v
    port map (
            O => \N__52469\,
            I => \N__52393\
        );

    \I__12750\ : InMux
    port map (
            O => \N__52466\,
            I => \N__52390\
        );

    \I__12749\ : Span4Mux_h
    port map (
            O => \N__52463\,
            I => \N__52385\
        );

    \I__12748\ : Span4Mux_h
    port map (
            O => \N__52456\,
            I => \N__52385\
        );

    \I__12747\ : Sp12to4
    port map (
            O => \N__52449\,
            I => \N__52382\
        );

    \I__12746\ : InMux
    port map (
            O => \N__52448\,
            I => \N__52379\
        );

    \I__12745\ : InMux
    port map (
            O => \N__52447\,
            I => \N__52376\
        );

    \I__12744\ : Span4Mux_v
    port map (
            O => \N__52444\,
            I => \N__52371\
        );

    \I__12743\ : Span4Mux_h
    port map (
            O => \N__52437\,
            I => \N__52371\
        );

    \I__12742\ : LocalMux
    port map (
            O => \N__52434\,
            I => \N__52360\
        );

    \I__12741\ : Span12Mux_v
    port map (
            O => \N__52429\,
            I => \N__52360\
        );

    \I__12740\ : LocalMux
    port map (
            O => \N__52426\,
            I => \N__52360\
        );

    \I__12739\ : Span12Mux_s6_v
    port map (
            O => \N__52419\,
            I => \N__52360\
        );

    \I__12738\ : Span12Mux_s11_h
    port map (
            O => \N__52416\,
            I => \N__52360\
        );

    \I__12737\ : Span4Mux_v
    port map (
            O => \N__52401\,
            I => \N__52357\
        );

    \I__12736\ : Span4Mux_h
    port map (
            O => \N__52396\,
            I => \N__52354\
        );

    \I__12735\ : Span12Mux_h
    port map (
            O => \N__52393\,
            I => \N__52351\
        );

    \I__12734\ : LocalMux
    port map (
            O => \N__52390\,
            I => \N__52344\
        );

    \I__12733\ : Sp12to4
    port map (
            O => \N__52385\,
            I => \N__52344\
        );

    \I__12732\ : Span12Mux_h
    port map (
            O => \N__52382\,
            I => \N__52344\
        );

    \I__12731\ : LocalMux
    port map (
            O => \N__52379\,
            I => \opZ0Z_2\
        );

    \I__12730\ : LocalMux
    port map (
            O => \N__52376\,
            I => \opZ0Z_2\
        );

    \I__12729\ : Odrv4
    port map (
            O => \N__52371\,
            I => \opZ0Z_2\
        );

    \I__12728\ : Odrv12
    port map (
            O => \N__52360\,
            I => \opZ0Z_2\
        );

    \I__12727\ : Odrv4
    port map (
            O => \N__52357\,
            I => \opZ0Z_2\
        );

    \I__12726\ : Odrv4
    port map (
            O => \N__52354\,
            I => \opZ0Z_2\
        );

    \I__12725\ : Odrv12
    port map (
            O => \N__52351\,
            I => \opZ0Z_2\
        );

    \I__12724\ : Odrv12
    port map (
            O => \N__52344\,
            I => \opZ0Z_2\
        );

    \I__12723\ : InMux
    port map (
            O => \N__52327\,
            I => \N__52317\
        );

    \I__12722\ : InMux
    port map (
            O => \N__52326\,
            I => \N__52314\
        );

    \I__12721\ : InMux
    port map (
            O => \N__52325\,
            I => \N__52311\
        );

    \I__12720\ : InMux
    port map (
            O => \N__52324\,
            I => \N__52303\
        );

    \I__12719\ : InMux
    port map (
            O => \N__52323\,
            I => \N__52303\
        );

    \I__12718\ : InMux
    port map (
            O => \N__52322\,
            I => \N__52294\
        );

    \I__12717\ : InMux
    port map (
            O => \N__52321\,
            I => \N__52294\
        );

    \I__12716\ : InMux
    port map (
            O => \N__52320\,
            I => \N__52290\
        );

    \I__12715\ : LocalMux
    port map (
            O => \N__52317\,
            I => \N__52287\
        );

    \I__12714\ : LocalMux
    port map (
            O => \N__52314\,
            I => \N__52284\
        );

    \I__12713\ : LocalMux
    port map (
            O => \N__52311\,
            I => \N__52281\
        );

    \I__12712\ : InMux
    port map (
            O => \N__52310\,
            I => \N__52278\
        );

    \I__12711\ : InMux
    port map (
            O => \N__52309\,
            I => \N__52272\
        );

    \I__12710\ : CascadeMux
    port map (
            O => \N__52308\,
            I => \N__52269\
        );

    \I__12709\ : LocalMux
    port map (
            O => \N__52303\,
            I => \N__52266\
        );

    \I__12708\ : InMux
    port map (
            O => \N__52302\,
            I => \N__52263\
        );

    \I__12707\ : InMux
    port map (
            O => \N__52301\,
            I => \N__52260\
        );

    \I__12706\ : InMux
    port map (
            O => \N__52300\,
            I => \N__52257\
        );

    \I__12705\ : InMux
    port map (
            O => \N__52299\,
            I => \N__52250\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__52294\,
            I => \N__52247\
        );

    \I__12703\ : InMux
    port map (
            O => \N__52293\,
            I => \N__52244\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__52290\,
            I => \N__52241\
        );

    \I__12701\ : Span4Mux_v
    port map (
            O => \N__52287\,
            I => \N__52232\
        );

    \I__12700\ : Span4Mux_v
    port map (
            O => \N__52284\,
            I => \N__52232\
        );

    \I__12699\ : Span4Mux_h
    port map (
            O => \N__52281\,
            I => \N__52232\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__52278\,
            I => \N__52232\
        );

    \I__12697\ : InMux
    port map (
            O => \N__52277\,
            I => \N__52229\
        );

    \I__12696\ : InMux
    port map (
            O => \N__52276\,
            I => \N__52223\
        );

    \I__12695\ : InMux
    port map (
            O => \N__52275\,
            I => \N__52223\
        );

    \I__12694\ : LocalMux
    port map (
            O => \N__52272\,
            I => \N__52218\
        );

    \I__12693\ : InMux
    port map (
            O => \N__52269\,
            I => \N__52215\
        );

    \I__12692\ : Span4Mux_v
    port map (
            O => \N__52266\,
            I => \N__52212\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__52263\,
            I => \N__52205\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__52260\,
            I => \N__52205\
        );

    \I__12689\ : LocalMux
    port map (
            O => \N__52257\,
            I => \N__52205\
        );

    \I__12688\ : InMux
    port map (
            O => \N__52256\,
            I => \N__52200\
        );

    \I__12687\ : InMux
    port map (
            O => \N__52255\,
            I => \N__52200\
        );

    \I__12686\ : CascadeMux
    port map (
            O => \N__52254\,
            I => \N__52195\
        );

    \I__12685\ : InMux
    port map (
            O => \N__52253\,
            I => \N__52192\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__52250\,
            I => \N__52189\
        );

    \I__12683\ : Span4Mux_v
    port map (
            O => \N__52247\,
            I => \N__52184\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__52244\,
            I => \N__52184\
        );

    \I__12681\ : Span4Mux_v
    port map (
            O => \N__52241\,
            I => \N__52177\
        );

    \I__12680\ : Span4Mux_v
    port map (
            O => \N__52232\,
            I => \N__52177\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__52229\,
            I => \N__52177\
        );

    \I__12678\ : CascadeMux
    port map (
            O => \N__52228\,
            I => \N__52174\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__52223\,
            I => \N__52171\
        );

    \I__12676\ : InMux
    port map (
            O => \N__52222\,
            I => \N__52168\
        );

    \I__12675\ : InMux
    port map (
            O => \N__52221\,
            I => \N__52165\
        );

    \I__12674\ : Span4Mux_v
    port map (
            O => \N__52218\,
            I => \N__52162\
        );

    \I__12673\ : LocalMux
    port map (
            O => \N__52215\,
            I => \N__52159\
        );

    \I__12672\ : Span4Mux_h
    port map (
            O => \N__52212\,
            I => \N__52152\
        );

    \I__12671\ : Span4Mux_v
    port map (
            O => \N__52205\,
            I => \N__52152\
        );

    \I__12670\ : LocalMux
    port map (
            O => \N__52200\,
            I => \N__52152\
        );

    \I__12669\ : InMux
    port map (
            O => \N__52199\,
            I => \N__52144\
        );

    \I__12668\ : InMux
    port map (
            O => \N__52198\,
            I => \N__52144\
        );

    \I__12667\ : InMux
    port map (
            O => \N__52195\,
            I => \N__52144\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__52192\,
            I => \N__52140\
        );

    \I__12665\ : Span4Mux_s3_h
    port map (
            O => \N__52189\,
            I => \N__52136\
        );

    \I__12664\ : Span4Mux_v
    port map (
            O => \N__52184\,
            I => \N__52131\
        );

    \I__12663\ : Span4Mux_h
    port map (
            O => \N__52177\,
            I => \N__52131\
        );

    \I__12662\ : InMux
    port map (
            O => \N__52174\,
            I => \N__52128\
        );

    \I__12661\ : Span4Mux_s3_h
    port map (
            O => \N__52171\,
            I => \N__52123\
        );

    \I__12660\ : LocalMux
    port map (
            O => \N__52168\,
            I => \N__52123\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__52165\,
            I => \N__52118\
        );

    \I__12658\ : Span4Mux_v
    port map (
            O => \N__52162\,
            I => \N__52111\
        );

    \I__12657\ : Span4Mux_v
    port map (
            O => \N__52159\,
            I => \N__52111\
        );

    \I__12656\ : Span4Mux_v
    port map (
            O => \N__52152\,
            I => \N__52111\
        );

    \I__12655\ : InMux
    port map (
            O => \N__52151\,
            I => \N__52108\
        );

    \I__12654\ : LocalMux
    port map (
            O => \N__52144\,
            I => \N__52105\
        );

    \I__12653\ : InMux
    port map (
            O => \N__52143\,
            I => \N__52099\
        );

    \I__12652\ : Span4Mux_h
    port map (
            O => \N__52140\,
            I => \N__52096\
        );

    \I__12651\ : InMux
    port map (
            O => \N__52139\,
            I => \N__52093\
        );

    \I__12650\ : Span4Mux_v
    port map (
            O => \N__52136\,
            I => \N__52084\
        );

    \I__12649\ : Span4Mux_h
    port map (
            O => \N__52131\,
            I => \N__52084\
        );

    \I__12648\ : LocalMux
    port map (
            O => \N__52128\,
            I => \N__52084\
        );

    \I__12647\ : Span4Mux_v
    port map (
            O => \N__52123\,
            I => \N__52084\
        );

    \I__12646\ : InMux
    port map (
            O => \N__52122\,
            I => \N__52079\
        );

    \I__12645\ : InMux
    port map (
            O => \N__52121\,
            I => \N__52079\
        );

    \I__12644\ : Span12Mux_v
    port map (
            O => \N__52118\,
            I => \N__52070\
        );

    \I__12643\ : Sp12to4
    port map (
            O => \N__52111\,
            I => \N__52070\
        );

    \I__12642\ : LocalMux
    port map (
            O => \N__52108\,
            I => \N__52070\
        );

    \I__12641\ : Span12Mux_s4_v
    port map (
            O => \N__52105\,
            I => \N__52070\
        );

    \I__12640\ : InMux
    port map (
            O => \N__52104\,
            I => \N__52063\
        );

    \I__12639\ : InMux
    port map (
            O => \N__52103\,
            I => \N__52063\
        );

    \I__12638\ : InMux
    port map (
            O => \N__52102\,
            I => \N__52063\
        );

    \I__12637\ : LocalMux
    port map (
            O => \N__52099\,
            I => \ALU.a_9\
        );

    \I__12636\ : Odrv4
    port map (
            O => \N__52096\,
            I => \ALU.a_9\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__52093\,
            I => \ALU.a_9\
        );

    \I__12634\ : Odrv4
    port map (
            O => \N__52084\,
            I => \ALU.a_9\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__52079\,
            I => \ALU.a_9\
        );

    \I__12632\ : Odrv12
    port map (
            O => \N__52070\,
            I => \ALU.a_9\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__52063\,
            I => \ALU.a_9\
        );

    \I__12630\ : InMux
    port map (
            O => \N__52048\,
            I => \N__52045\
        );

    \I__12629\ : LocalMux
    port map (
            O => \N__52045\,
            I => \N__52042\
        );

    \I__12628\ : Span4Mux_v
    port map (
            O => \N__52042\,
            I => \N__52039\
        );

    \I__12627\ : Odrv4
    port map (
            O => \N__52039\,
            I => \ALU.r0_12_prm_4_9_s1_c_RNOZ0\
        );

    \I__12626\ : InMux
    port map (
            O => \N__52036\,
            I => \N__52030\
        );

    \I__12625\ : CascadeMux
    port map (
            O => \N__52035\,
            I => \N__52025\
        );

    \I__12624\ : InMux
    port map (
            O => \N__52034\,
            I => \N__52021\
        );

    \I__12623\ : InMux
    port map (
            O => \N__52033\,
            I => \N__52018\
        );

    \I__12622\ : LocalMux
    port map (
            O => \N__52030\,
            I => \N__52015\
        );

    \I__12621\ : CascadeMux
    port map (
            O => \N__52029\,
            I => \N__52012\
        );

    \I__12620\ : InMux
    port map (
            O => \N__52028\,
            I => \N__52009\
        );

    \I__12619\ : InMux
    port map (
            O => \N__52025\,
            I => \N__52004\
        );

    \I__12618\ : InMux
    port map (
            O => \N__52024\,
            I => \N__52004\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__52021\,
            I => \N__51997\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__52018\,
            I => \N__51992\
        );

    \I__12615\ : Span4Mux_v
    port map (
            O => \N__52015\,
            I => \N__51992\
        );

    \I__12614\ : InMux
    port map (
            O => \N__52012\,
            I => \N__51989\
        );

    \I__12613\ : LocalMux
    port map (
            O => \N__52009\,
            I => \N__51984\
        );

    \I__12612\ : LocalMux
    port map (
            O => \N__52004\,
            I => \N__51980\
        );

    \I__12611\ : InMux
    port map (
            O => \N__52003\,
            I => \N__51976\
        );

    \I__12610\ : InMux
    port map (
            O => \N__52002\,
            I => \N__51972\
        );

    \I__12609\ : InMux
    port map (
            O => \N__52001\,
            I => \N__51969\
        );

    \I__12608\ : InMux
    port map (
            O => \N__52000\,
            I => \N__51966\
        );

    \I__12607\ : Span4Mux_v
    port map (
            O => \N__51997\,
            I => \N__51959\
        );

    \I__12606\ : Span4Mux_h
    port map (
            O => \N__51992\,
            I => \N__51959\
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__51989\,
            I => \N__51959\
        );

    \I__12604\ : InMux
    port map (
            O => \N__51988\,
            I => \N__51953\
        );

    \I__12603\ : InMux
    port map (
            O => \N__51987\,
            I => \N__51953\
        );

    \I__12602\ : Span4Mux_h
    port map (
            O => \N__51984\,
            I => \N__51950\
        );

    \I__12601\ : InMux
    port map (
            O => \N__51983\,
            I => \N__51947\
        );

    \I__12600\ : Span4Mux_h
    port map (
            O => \N__51980\,
            I => \N__51944\
        );

    \I__12599\ : CascadeMux
    port map (
            O => \N__51979\,
            I => \N__51941\
        );

    \I__12598\ : LocalMux
    port map (
            O => \N__51976\,
            I => \N__51936\
        );

    \I__12597\ : InMux
    port map (
            O => \N__51975\,
            I => \N__51933\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__51972\,
            I => \N__51928\
        );

    \I__12595\ : LocalMux
    port map (
            O => \N__51969\,
            I => \N__51928\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__51966\,
            I => \N__51923\
        );

    \I__12593\ : Span4Mux_h
    port map (
            O => \N__51959\,
            I => \N__51923\
        );

    \I__12592\ : CascadeMux
    port map (
            O => \N__51958\,
            I => \N__51920\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__51953\,
            I => \N__51914\
        );

    \I__12590\ : Span4Mux_h
    port map (
            O => \N__51950\,
            I => \N__51909\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__51947\,
            I => \N__51909\
        );

    \I__12588\ : Span4Mux_h
    port map (
            O => \N__51944\,
            I => \N__51905\
        );

    \I__12587\ : InMux
    port map (
            O => \N__51941\,
            I => \N__51902\
        );

    \I__12586\ : InMux
    port map (
            O => \N__51940\,
            I => \N__51899\
        );

    \I__12585\ : InMux
    port map (
            O => \N__51939\,
            I => \N__51896\
        );

    \I__12584\ : Span4Mux_h
    port map (
            O => \N__51936\,
            I => \N__51891\
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__51933\,
            I => \N__51891\
        );

    \I__12582\ : Span12Mux_h
    port map (
            O => \N__51928\,
            I => \N__51888\
        );

    \I__12581\ : Span4Mux_h
    port map (
            O => \N__51923\,
            I => \N__51885\
        );

    \I__12580\ : InMux
    port map (
            O => \N__51920\,
            I => \N__51878\
        );

    \I__12579\ : InMux
    port map (
            O => \N__51919\,
            I => \N__51878\
        );

    \I__12578\ : InMux
    port map (
            O => \N__51918\,
            I => \N__51878\
        );

    \I__12577\ : InMux
    port map (
            O => \N__51917\,
            I => \N__51875\
        );

    \I__12576\ : Span4Mux_v
    port map (
            O => \N__51914\,
            I => \N__51870\
        );

    \I__12575\ : Span4Mux_v
    port map (
            O => \N__51909\,
            I => \N__51870\
        );

    \I__12574\ : InMux
    port map (
            O => \N__51908\,
            I => \N__51867\
        );

    \I__12573\ : Span4Mux_v
    port map (
            O => \N__51905\,
            I => \N__51856\
        );

    \I__12572\ : LocalMux
    port map (
            O => \N__51902\,
            I => \N__51856\
        );

    \I__12571\ : LocalMux
    port map (
            O => \N__51899\,
            I => \N__51856\
        );

    \I__12570\ : LocalMux
    port map (
            O => \N__51896\,
            I => \N__51856\
        );

    \I__12569\ : Span4Mux_h
    port map (
            O => \N__51891\,
            I => \N__51856\
        );

    \I__12568\ : Odrv12
    port map (
            O => \N__51888\,
            I => \ALU.b_10\
        );

    \I__12567\ : Odrv4
    port map (
            O => \N__51885\,
            I => \ALU.b_10\
        );

    \I__12566\ : LocalMux
    port map (
            O => \N__51878\,
            I => \ALU.b_10\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__51875\,
            I => \ALU.b_10\
        );

    \I__12564\ : Odrv4
    port map (
            O => \N__51870\,
            I => \ALU.b_10\
        );

    \I__12563\ : LocalMux
    port map (
            O => \N__51867\,
            I => \ALU.b_10\
        );

    \I__12562\ : Odrv4
    port map (
            O => \N__51856\,
            I => \ALU.b_10\
        );

    \I__12561\ : InMux
    port map (
            O => \N__51841\,
            I => \N__51833\
        );

    \I__12560\ : InMux
    port map (
            O => \N__51840\,
            I => \N__51822\
        );

    \I__12559\ : CascadeMux
    port map (
            O => \N__51839\,
            I => \N__51819\
        );

    \I__12558\ : CascadeMux
    port map (
            O => \N__51838\,
            I => \N__51816\
        );

    \I__12557\ : InMux
    port map (
            O => \N__51837\,
            I => \N__51812\
        );

    \I__12556\ : InMux
    port map (
            O => \N__51836\,
            I => \N__51801\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__51833\,
            I => \N__51798\
        );

    \I__12554\ : InMux
    port map (
            O => \N__51832\,
            I => \N__51791\
        );

    \I__12553\ : InMux
    port map (
            O => \N__51831\,
            I => \N__51788\
        );

    \I__12552\ : InMux
    port map (
            O => \N__51830\,
            I => \N__51781\
        );

    \I__12551\ : InMux
    port map (
            O => \N__51829\,
            I => \N__51781\
        );

    \I__12550\ : InMux
    port map (
            O => \N__51828\,
            I => \N__51781\
        );

    \I__12549\ : InMux
    port map (
            O => \N__51827\,
            I => \N__51776\
        );

    \I__12548\ : InMux
    port map (
            O => \N__51826\,
            I => \N__51776\
        );

    \I__12547\ : InMux
    port map (
            O => \N__51825\,
            I => \N__51773\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__51822\,
            I => \N__51770\
        );

    \I__12545\ : InMux
    port map (
            O => \N__51819\,
            I => \N__51767\
        );

    \I__12544\ : InMux
    port map (
            O => \N__51816\,
            I => \N__51762\
        );

    \I__12543\ : InMux
    port map (
            O => \N__51815\,
            I => \N__51762\
        );

    \I__12542\ : LocalMux
    port map (
            O => \N__51812\,
            I => \N__51759\
        );

    \I__12541\ : InMux
    port map (
            O => \N__51811\,
            I => \N__51756\
        );

    \I__12540\ : InMux
    port map (
            O => \N__51810\,
            I => \N__51751\
        );

    \I__12539\ : InMux
    port map (
            O => \N__51809\,
            I => \N__51751\
        );

    \I__12538\ : InMux
    port map (
            O => \N__51808\,
            I => \N__51748\
        );

    \I__12537\ : CascadeMux
    port map (
            O => \N__51807\,
            I => \N__51744\
        );

    \I__12536\ : CascadeMux
    port map (
            O => \N__51806\,
            I => \N__51739\
        );

    \I__12535\ : InMux
    port map (
            O => \N__51805\,
            I => \N__51736\
        );

    \I__12534\ : InMux
    port map (
            O => \N__51804\,
            I => \N__51733\
        );

    \I__12533\ : LocalMux
    port map (
            O => \N__51801\,
            I => \N__51729\
        );

    \I__12532\ : Span4Mux_v
    port map (
            O => \N__51798\,
            I => \N__51726\
        );

    \I__12531\ : InMux
    port map (
            O => \N__51797\,
            I => \N__51723\
        );

    \I__12530\ : InMux
    port map (
            O => \N__51796\,
            I => \N__51720\
        );

    \I__12529\ : InMux
    port map (
            O => \N__51795\,
            I => \N__51717\
        );

    \I__12528\ : InMux
    port map (
            O => \N__51794\,
            I => \N__51713\
        );

    \I__12527\ : LocalMux
    port map (
            O => \N__51791\,
            I => \N__51702\
        );

    \I__12526\ : LocalMux
    port map (
            O => \N__51788\,
            I => \N__51702\
        );

    \I__12525\ : LocalMux
    port map (
            O => \N__51781\,
            I => \N__51702\
        );

    \I__12524\ : LocalMux
    port map (
            O => \N__51776\,
            I => \N__51702\
        );

    \I__12523\ : LocalMux
    port map (
            O => \N__51773\,
            I => \N__51702\
        );

    \I__12522\ : Span4Mux_v
    port map (
            O => \N__51770\,
            I => \N__51699\
        );

    \I__12521\ : LocalMux
    port map (
            O => \N__51767\,
            I => \N__51696\
        );

    \I__12520\ : LocalMux
    port map (
            O => \N__51762\,
            I => \N__51691\
        );

    \I__12519\ : Span4Mux_v
    port map (
            O => \N__51759\,
            I => \N__51691\
        );

    \I__12518\ : LocalMux
    port map (
            O => \N__51756\,
            I => \N__51688\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__51751\,
            I => \N__51683\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__51748\,
            I => \N__51683\
        );

    \I__12515\ : InMux
    port map (
            O => \N__51747\,
            I => \N__51680\
        );

    \I__12514\ : InMux
    port map (
            O => \N__51744\,
            I => \N__51677\
        );

    \I__12513\ : InMux
    port map (
            O => \N__51743\,
            I => \N__51672\
        );

    \I__12512\ : InMux
    port map (
            O => \N__51742\,
            I => \N__51672\
        );

    \I__12511\ : InMux
    port map (
            O => \N__51739\,
            I => \N__51669\
        );

    \I__12510\ : LocalMux
    port map (
            O => \N__51736\,
            I => \N__51666\
        );

    \I__12509\ : LocalMux
    port map (
            O => \N__51733\,
            I => \N__51663\
        );

    \I__12508\ : InMux
    port map (
            O => \N__51732\,
            I => \N__51660\
        );

    \I__12507\ : Span12Mux_s4_h
    port map (
            O => \N__51729\,
            I => \N__51653\
        );

    \I__12506\ : Sp12to4
    port map (
            O => \N__51726\,
            I => \N__51653\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__51723\,
            I => \N__51653\
        );

    \I__12504\ : LocalMux
    port map (
            O => \N__51720\,
            I => \N__51649\
        );

    \I__12503\ : LocalMux
    port map (
            O => \N__51717\,
            I => \N__51646\
        );

    \I__12502\ : InMux
    port map (
            O => \N__51716\,
            I => \N__51643\
        );

    \I__12501\ : LocalMux
    port map (
            O => \N__51713\,
            I => \N__51638\
        );

    \I__12500\ : Span4Mux_v
    port map (
            O => \N__51702\,
            I => \N__51638\
        );

    \I__12499\ : Span4Mux_h
    port map (
            O => \N__51699\,
            I => \N__51631\
        );

    \I__12498\ : Span4Mux_v
    port map (
            O => \N__51696\,
            I => \N__51631\
        );

    \I__12497\ : Span4Mux_h
    port map (
            O => \N__51691\,
            I => \N__51631\
        );

    \I__12496\ : Span4Mux_v
    port map (
            O => \N__51688\,
            I => \N__51626\
        );

    \I__12495\ : Span4Mux_v
    port map (
            O => \N__51683\,
            I => \N__51626\
        );

    \I__12494\ : LocalMux
    port map (
            O => \N__51680\,
            I => \N__51623\
        );

    \I__12493\ : LocalMux
    port map (
            O => \N__51677\,
            I => \N__51620\
        );

    \I__12492\ : LocalMux
    port map (
            O => \N__51672\,
            I => \N__51617\
        );

    \I__12491\ : LocalMux
    port map (
            O => \N__51669\,
            I => \N__51614\
        );

    \I__12490\ : Span4Mux_v
    port map (
            O => \N__51666\,
            I => \N__51607\
        );

    \I__12489\ : Span4Mux_h
    port map (
            O => \N__51663\,
            I => \N__51607\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__51660\,
            I => \N__51607\
        );

    \I__12487\ : Span12Mux_h
    port map (
            O => \N__51653\,
            I => \N__51604\
        );

    \I__12486\ : InMux
    port map (
            O => \N__51652\,
            I => \N__51601\
        );

    \I__12485\ : Sp12to4
    port map (
            O => \N__51649\,
            I => \N__51594\
        );

    \I__12484\ : Span12Mux_s9_v
    port map (
            O => \N__51646\,
            I => \N__51594\
        );

    \I__12483\ : LocalMux
    port map (
            O => \N__51643\,
            I => \N__51594\
        );

    \I__12482\ : Span4Mux_h
    port map (
            O => \N__51638\,
            I => \N__51587\
        );

    \I__12481\ : Span4Mux_h
    port map (
            O => \N__51631\,
            I => \N__51587\
        );

    \I__12480\ : Span4Mux_h
    port map (
            O => \N__51626\,
            I => \N__51587\
        );

    \I__12479\ : Span4Mux_h
    port map (
            O => \N__51623\,
            I => \N__51582\
        );

    \I__12478\ : Span4Mux_v
    port map (
            O => \N__51620\,
            I => \N__51582\
        );

    \I__12477\ : Span4Mux_h
    port map (
            O => \N__51617\,
            I => \N__51575\
        );

    \I__12476\ : Span4Mux_v
    port map (
            O => \N__51614\,
            I => \N__51575\
        );

    \I__12475\ : Span4Mux_h
    port map (
            O => \N__51607\,
            I => \N__51575\
        );

    \I__12474\ : Odrv12
    port map (
            O => \N__51604\,
            I => \ALU.a_10\
        );

    \I__12473\ : LocalMux
    port map (
            O => \N__51601\,
            I => \ALU.a_10\
        );

    \I__12472\ : Odrv12
    port map (
            O => \N__51594\,
            I => \ALU.a_10\
        );

    \I__12471\ : Odrv4
    port map (
            O => \N__51587\,
            I => \ALU.a_10\
        );

    \I__12470\ : Odrv4
    port map (
            O => \N__51582\,
            I => \ALU.a_10\
        );

    \I__12469\ : Odrv4
    port map (
            O => \N__51575\,
            I => \ALU.a_10\
        );

    \I__12468\ : CascadeMux
    port map (
            O => \N__51562\,
            I => \N__51559\
        );

    \I__12467\ : InMux
    port map (
            O => \N__51559\,
            I => \N__51556\
        );

    \I__12466\ : LocalMux
    port map (
            O => \N__51556\,
            I => \N__51553\
        );

    \I__12465\ : Span4Mux_h
    port map (
            O => \N__51553\,
            I => \N__51550\
        );

    \I__12464\ : Span4Mux_h
    port map (
            O => \N__51550\,
            I => \N__51547\
        );

    \I__12463\ : Span4Mux_h
    port map (
            O => \N__51547\,
            I => \N__51544\
        );

    \I__12462\ : Odrv4
    port map (
            O => \N__51544\,
            I => \ALU.r0_12_prm_7_10_s0_c_RNOZ0\
        );

    \I__12461\ : CascadeMux
    port map (
            O => \N__51541\,
            I => \N__51538\
        );

    \I__12460\ : InMux
    port map (
            O => \N__51538\,
            I => \N__51534\
        );

    \I__12459\ : CascadeMux
    port map (
            O => \N__51537\,
            I => \N__51524\
        );

    \I__12458\ : LocalMux
    port map (
            O => \N__51534\,
            I => \N__51515\
        );

    \I__12457\ : CascadeMux
    port map (
            O => \N__51533\,
            I => \N__51510\
        );

    \I__12456\ : CascadeMux
    port map (
            O => \N__51532\,
            I => \N__51504\
        );

    \I__12455\ : CascadeMux
    port map (
            O => \N__51531\,
            I => \N__51501\
        );

    \I__12454\ : CascadeMux
    port map (
            O => \N__51530\,
            I => \N__51495\
        );

    \I__12453\ : CascadeMux
    port map (
            O => \N__51529\,
            I => \N__51492\
        );

    \I__12452\ : CascadeMux
    port map (
            O => \N__51528\,
            I => \N__51488\
        );

    \I__12451\ : CascadeMux
    port map (
            O => \N__51527\,
            I => \N__51485\
        );

    \I__12450\ : InMux
    port map (
            O => \N__51524\,
            I => \N__51479\
        );

    \I__12449\ : InMux
    port map (
            O => \N__51523\,
            I => \N__51476\
        );

    \I__12448\ : CascadeMux
    port map (
            O => \N__51522\,
            I => \N__51469\
        );

    \I__12447\ : CascadeMux
    port map (
            O => \N__51521\,
            I => \N__51466\
        );

    \I__12446\ : CascadeMux
    port map (
            O => \N__51520\,
            I => \N__51462\
        );

    \I__12445\ : InMux
    port map (
            O => \N__51519\,
            I => \N__51457\
        );

    \I__12444\ : InMux
    port map (
            O => \N__51518\,
            I => \N__51457\
        );

    \I__12443\ : Span4Mux_v
    port map (
            O => \N__51515\,
            I => \N__51454\
        );

    \I__12442\ : InMux
    port map (
            O => \N__51514\,
            I => \N__51447\
        );

    \I__12441\ : InMux
    port map (
            O => \N__51513\,
            I => \N__51447\
        );

    \I__12440\ : InMux
    port map (
            O => \N__51510\,
            I => \N__51447\
        );

    \I__12439\ : InMux
    port map (
            O => \N__51509\,
            I => \N__51443\
        );

    \I__12438\ : InMux
    port map (
            O => \N__51508\,
            I => \N__51438\
        );

    \I__12437\ : InMux
    port map (
            O => \N__51507\,
            I => \N__51435\
        );

    \I__12436\ : InMux
    port map (
            O => \N__51504\,
            I => \N__51430\
        );

    \I__12435\ : InMux
    port map (
            O => \N__51501\,
            I => \N__51430\
        );

    \I__12434\ : CascadeMux
    port map (
            O => \N__51500\,
            I => \N__51427\
        );

    \I__12433\ : CascadeMux
    port map (
            O => \N__51499\,
            I => \N__51424\
        );

    \I__12432\ : InMux
    port map (
            O => \N__51498\,
            I => \N__51420\
        );

    \I__12431\ : InMux
    port map (
            O => \N__51495\,
            I => \N__51415\
        );

    \I__12430\ : InMux
    port map (
            O => \N__51492\,
            I => \N__51415\
        );

    \I__12429\ : CascadeMux
    port map (
            O => \N__51491\,
            I => \N__51411\
        );

    \I__12428\ : InMux
    port map (
            O => \N__51488\,
            I => \N__51406\
        );

    \I__12427\ : InMux
    port map (
            O => \N__51485\,
            I => \N__51406\
        );

    \I__12426\ : CascadeMux
    port map (
            O => \N__51484\,
            I => \N__51403\
        );

    \I__12425\ : CascadeMux
    port map (
            O => \N__51483\,
            I => \N__51400\
        );

    \I__12424\ : CascadeMux
    port map (
            O => \N__51482\,
            I => \N__51397\
        );

    \I__12423\ : LocalMux
    port map (
            O => \N__51479\,
            I => \N__51392\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__51476\,
            I => \N__51392\
        );

    \I__12421\ : InMux
    port map (
            O => \N__51475\,
            I => \N__51389\
        );

    \I__12420\ : InMux
    port map (
            O => \N__51474\,
            I => \N__51386\
        );

    \I__12419\ : InMux
    port map (
            O => \N__51473\,
            I => \N__51381\
        );

    \I__12418\ : InMux
    port map (
            O => \N__51472\,
            I => \N__51381\
        );

    \I__12417\ : InMux
    port map (
            O => \N__51469\,
            I => \N__51378\
        );

    \I__12416\ : InMux
    port map (
            O => \N__51466\,
            I => \N__51371\
        );

    \I__12415\ : InMux
    port map (
            O => \N__51465\,
            I => \N__51371\
        );

    \I__12414\ : InMux
    port map (
            O => \N__51462\,
            I => \N__51371\
        );

    \I__12413\ : LocalMux
    port map (
            O => \N__51457\,
            I => \N__51368\
        );

    \I__12412\ : Span4Mux_h
    port map (
            O => \N__51454\,
            I => \N__51363\
        );

    \I__12411\ : LocalMux
    port map (
            O => \N__51447\,
            I => \N__51363\
        );

    \I__12410\ : CascadeMux
    port map (
            O => \N__51446\,
            I => \N__51360\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__51443\,
            I => \N__51356\
        );

    \I__12408\ : InMux
    port map (
            O => \N__51442\,
            I => \N__51353\
        );

    \I__12407\ : InMux
    port map (
            O => \N__51441\,
            I => \N__51350\
        );

    \I__12406\ : LocalMux
    port map (
            O => \N__51438\,
            I => \N__51347\
        );

    \I__12405\ : LocalMux
    port map (
            O => \N__51435\,
            I => \N__51342\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__51430\,
            I => \N__51342\
        );

    \I__12403\ : InMux
    port map (
            O => \N__51427\,
            I => \N__51337\
        );

    \I__12402\ : InMux
    port map (
            O => \N__51424\,
            I => \N__51337\
        );

    \I__12401\ : InMux
    port map (
            O => \N__51423\,
            I => \N__51334\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__51420\,
            I => \N__51329\
        );

    \I__12399\ : LocalMux
    port map (
            O => \N__51415\,
            I => \N__51329\
        );

    \I__12398\ : InMux
    port map (
            O => \N__51414\,
            I => \N__51326\
        );

    \I__12397\ : InMux
    port map (
            O => \N__51411\,
            I => \N__51323\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__51406\,
            I => \N__51320\
        );

    \I__12395\ : InMux
    port map (
            O => \N__51403\,
            I => \N__51315\
        );

    \I__12394\ : InMux
    port map (
            O => \N__51400\,
            I => \N__51315\
        );

    \I__12393\ : InMux
    port map (
            O => \N__51397\,
            I => \N__51312\
        );

    \I__12392\ : Span4Mux_v
    port map (
            O => \N__51392\,
            I => \N__51305\
        );

    \I__12391\ : LocalMux
    port map (
            O => \N__51389\,
            I => \N__51305\
        );

    \I__12390\ : LocalMux
    port map (
            O => \N__51386\,
            I => \N__51305\
        );

    \I__12389\ : LocalMux
    port map (
            O => \N__51381\,
            I => \N__51297\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__51378\,
            I => \N__51291\
        );

    \I__12387\ : LocalMux
    port map (
            O => \N__51371\,
            I => \N__51291\
        );

    \I__12386\ : Span4Mux_v
    port map (
            O => \N__51368\,
            I => \N__51286\
        );

    \I__12385\ : Span4Mux_v
    port map (
            O => \N__51363\,
            I => \N__51286\
        );

    \I__12384\ : InMux
    port map (
            O => \N__51360\,
            I => \N__51281\
        );

    \I__12383\ : InMux
    port map (
            O => \N__51359\,
            I => \N__51281\
        );

    \I__12382\ : Span4Mux_s3_v
    port map (
            O => \N__51356\,
            I => \N__51276\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__51353\,
            I => \N__51276\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__51350\,
            I => \N__51269\
        );

    \I__12379\ : Span4Mux_h
    port map (
            O => \N__51347\,
            I => \N__51269\
        );

    \I__12378\ : Span4Mux_h
    port map (
            O => \N__51342\,
            I => \N__51269\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__51337\,
            I => \N__51265\
        );

    \I__12376\ : LocalMux
    port map (
            O => \N__51334\,
            I => \N__51258\
        );

    \I__12375\ : Span4Mux_h
    port map (
            O => \N__51329\,
            I => \N__51258\
        );

    \I__12374\ : LocalMux
    port map (
            O => \N__51326\,
            I => \N__51258\
        );

    \I__12373\ : LocalMux
    port map (
            O => \N__51323\,
            I => \N__51247\
        );

    \I__12372\ : Span4Mux_h
    port map (
            O => \N__51320\,
            I => \N__51247\
        );

    \I__12371\ : LocalMux
    port map (
            O => \N__51315\,
            I => \N__51247\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__51312\,
            I => \N__51247\
        );

    \I__12369\ : Span4Mux_v
    port map (
            O => \N__51305\,
            I => \N__51247\
        );

    \I__12368\ : CascadeMux
    port map (
            O => \N__51304\,
            I => \N__51241\
        );

    \I__12367\ : InMux
    port map (
            O => \N__51303\,
            I => \N__51238\
        );

    \I__12366\ : CascadeMux
    port map (
            O => \N__51302\,
            I => \N__51235\
        );

    \I__12365\ : CascadeMux
    port map (
            O => \N__51301\,
            I => \N__51232\
        );

    \I__12364\ : InMux
    port map (
            O => \N__51300\,
            I => \N__51228\
        );

    \I__12363\ : Span4Mux_h
    port map (
            O => \N__51297\,
            I => \N__51225\
        );

    \I__12362\ : CascadeMux
    port map (
            O => \N__51296\,
            I => \N__51218\
        );

    \I__12361\ : Span4Mux_v
    port map (
            O => \N__51291\,
            I => \N__51213\
        );

    \I__12360\ : Span4Mux_v
    port map (
            O => \N__51286\,
            I => \N__51213\
        );

    \I__12359\ : LocalMux
    port map (
            O => \N__51281\,
            I => \N__51205\
        );

    \I__12358\ : Span4Mux_h
    port map (
            O => \N__51276\,
            I => \N__51205\
        );

    \I__12357\ : Span4Mux_v
    port map (
            O => \N__51269\,
            I => \N__51205\
        );

    \I__12356\ : InMux
    port map (
            O => \N__51268\,
            I => \N__51202\
        );

    \I__12355\ : Span4Mux_v
    port map (
            O => \N__51265\,
            I => \N__51199\
        );

    \I__12354\ : Span4Mux_v
    port map (
            O => \N__51258\,
            I => \N__51196\
        );

    \I__12353\ : Span4Mux_v
    port map (
            O => \N__51247\,
            I => \N__51193\
        );

    \I__12352\ : InMux
    port map (
            O => \N__51246\,
            I => \N__51190\
        );

    \I__12351\ : InMux
    port map (
            O => \N__51245\,
            I => \N__51185\
        );

    \I__12350\ : InMux
    port map (
            O => \N__51244\,
            I => \N__51185\
        );

    \I__12349\ : InMux
    port map (
            O => \N__51241\,
            I => \N__51182\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__51238\,
            I => \N__51179\
        );

    \I__12347\ : InMux
    port map (
            O => \N__51235\,
            I => \N__51172\
        );

    \I__12346\ : InMux
    port map (
            O => \N__51232\,
            I => \N__51172\
        );

    \I__12345\ : InMux
    port map (
            O => \N__51231\,
            I => \N__51172\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__51228\,
            I => \N__51167\
        );

    \I__12343\ : Span4Mux_h
    port map (
            O => \N__51225\,
            I => \N__51167\
        );

    \I__12342\ : InMux
    port map (
            O => \N__51224\,
            I => \N__51164\
        );

    \I__12341\ : InMux
    port map (
            O => \N__51223\,
            I => \N__51159\
        );

    \I__12340\ : InMux
    port map (
            O => \N__51222\,
            I => \N__51159\
        );

    \I__12339\ : InMux
    port map (
            O => \N__51221\,
            I => \N__51154\
        );

    \I__12338\ : InMux
    port map (
            O => \N__51218\,
            I => \N__51154\
        );

    \I__12337\ : Span4Mux_v
    port map (
            O => \N__51213\,
            I => \N__51151\
        );

    \I__12336\ : InMux
    port map (
            O => \N__51212\,
            I => \N__51148\
        );

    \I__12335\ : Span4Mux_v
    port map (
            O => \N__51205\,
            I => \N__51143\
        );

    \I__12334\ : LocalMux
    port map (
            O => \N__51202\,
            I => \N__51143\
        );

    \I__12333\ : Span4Mux_s0_v
    port map (
            O => \N__51199\,
            I => \N__51136\
        );

    \I__12332\ : Span4Mux_s0_v
    port map (
            O => \N__51196\,
            I => \N__51136\
        );

    \I__12331\ : Span4Mux_s0_v
    port map (
            O => \N__51193\,
            I => \N__51136\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__51190\,
            I => \N__51123\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__51185\,
            I => \N__51123\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__51182\,
            I => \N__51123\
        );

    \I__12327\ : Span12Mux_v
    port map (
            O => \N__51179\,
            I => \N__51123\
        );

    \I__12326\ : LocalMux
    port map (
            O => \N__51172\,
            I => \N__51123\
        );

    \I__12325\ : Sp12to4
    port map (
            O => \N__51167\,
            I => \N__51123\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__51164\,
            I => \paramsZ0Z_3\
        );

    \I__12323\ : LocalMux
    port map (
            O => \N__51159\,
            I => \paramsZ0Z_3\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__51154\,
            I => \paramsZ0Z_3\
        );

    \I__12321\ : Odrv4
    port map (
            O => \N__51151\,
            I => \paramsZ0Z_3\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__51148\,
            I => \paramsZ0Z_3\
        );

    \I__12319\ : Odrv4
    port map (
            O => \N__51143\,
            I => \paramsZ0Z_3\
        );

    \I__12318\ : Odrv4
    port map (
            O => \N__51136\,
            I => \paramsZ0Z_3\
        );

    \I__12317\ : Odrv12
    port map (
            O => \N__51123\,
            I => \paramsZ0Z_3\
        );

    \I__12316\ : InMux
    port map (
            O => \N__51106\,
            I => \N__51093\
        );

    \I__12315\ : InMux
    port map (
            O => \N__51105\,
            I => \N__51093\
        );

    \I__12314\ : InMux
    port map (
            O => \N__51104\,
            I => \N__51090\
        );

    \I__12313\ : InMux
    port map (
            O => \N__51103\,
            I => \N__51084\
        );

    \I__12312\ : InMux
    port map (
            O => \N__51102\,
            I => \N__51081\
        );

    \I__12311\ : InMux
    port map (
            O => \N__51101\,
            I => \N__51075\
        );

    \I__12310\ : InMux
    port map (
            O => \N__51100\,
            I => \N__51075\
        );

    \I__12309\ : InMux
    port map (
            O => \N__51099\,
            I => \N__51071\
        );

    \I__12308\ : InMux
    port map (
            O => \N__51098\,
            I => \N__51068\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__51093\,
            I => \N__51065\
        );

    \I__12306\ : LocalMux
    port map (
            O => \N__51090\,
            I => \N__51062\
        );

    \I__12305\ : InMux
    port map (
            O => \N__51089\,
            I => \N__51059\
        );

    \I__12304\ : CascadeMux
    port map (
            O => \N__51088\,
            I => \N__51055\
        );

    \I__12303\ : CascadeMux
    port map (
            O => \N__51087\,
            I => \N__51051\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__51084\,
            I => \N__51048\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__51081\,
            I => \N__51044\
        );

    \I__12300\ : InMux
    port map (
            O => \N__51080\,
            I => \N__51041\
        );

    \I__12299\ : LocalMux
    port map (
            O => \N__51075\,
            I => \N__51034\
        );

    \I__12298\ : CascadeMux
    port map (
            O => \N__51074\,
            I => \N__51029\
        );

    \I__12297\ : LocalMux
    port map (
            O => \N__51071\,
            I => \N__51021\
        );

    \I__12296\ : LocalMux
    port map (
            O => \N__51068\,
            I => \N__51016\
        );

    \I__12295\ : Span4Mux_h
    port map (
            O => \N__51065\,
            I => \N__51016\
        );

    \I__12294\ : Span4Mux_v
    port map (
            O => \N__51062\,
            I => \N__51011\
        );

    \I__12293\ : LocalMux
    port map (
            O => \N__51059\,
            I => \N__51011\
        );

    \I__12292\ : InMux
    port map (
            O => \N__51058\,
            I => \N__51004\
        );

    \I__12291\ : InMux
    port map (
            O => \N__51055\,
            I => \N__51004\
        );

    \I__12290\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51004\
        );

    \I__12289\ : InMux
    port map (
            O => \N__51051\,
            I => \N__50996\
        );

    \I__12288\ : Span4Mux_v
    port map (
            O => \N__51048\,
            I => \N__50989\
        );

    \I__12287\ : InMux
    port map (
            O => \N__51047\,
            I => \N__50986\
        );

    \I__12286\ : Span4Mux_v
    port map (
            O => \N__51044\,
            I => \N__50979\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__51041\,
            I => \N__50979\
        );

    \I__12284\ : InMux
    port map (
            O => \N__51040\,
            I => \N__50974\
        );

    \I__12283\ : InMux
    port map (
            O => \N__51039\,
            I => \N__50974\
        );

    \I__12282\ : InMux
    port map (
            O => \N__51038\,
            I => \N__50971\
        );

    \I__12281\ : InMux
    port map (
            O => \N__51037\,
            I => \N__50968\
        );

    \I__12280\ : Span4Mux_h
    port map (
            O => \N__51034\,
            I => \N__50965\
        );

    \I__12279\ : InMux
    port map (
            O => \N__51033\,
            I => \N__50962\
        );

    \I__12278\ : InMux
    port map (
            O => \N__51032\,
            I => \N__50958\
        );

    \I__12277\ : InMux
    port map (
            O => \N__51029\,
            I => \N__50955\
        );

    \I__12276\ : InMux
    port map (
            O => \N__51028\,
            I => \N__50952\
        );

    \I__12275\ : InMux
    port map (
            O => \N__51027\,
            I => \N__50949\
        );

    \I__12274\ : InMux
    port map (
            O => \N__51026\,
            I => \N__50942\
        );

    \I__12273\ : InMux
    port map (
            O => \N__51025\,
            I => \N__50942\
        );

    \I__12272\ : InMux
    port map (
            O => \N__51024\,
            I => \N__50942\
        );

    \I__12271\ : Span4Mux_v
    port map (
            O => \N__51021\,
            I => \N__50933\
        );

    \I__12270\ : Span4Mux_h
    port map (
            O => \N__51016\,
            I => \N__50933\
        );

    \I__12269\ : Span4Mux_h
    port map (
            O => \N__51011\,
            I => \N__50933\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__51004\,
            I => \N__50933\
        );

    \I__12267\ : InMux
    port map (
            O => \N__51003\,
            I => \N__50926\
        );

    \I__12266\ : InMux
    port map (
            O => \N__51002\,
            I => \N__50926\
        );

    \I__12265\ : InMux
    port map (
            O => \N__51001\,
            I => \N__50921\
        );

    \I__12264\ : InMux
    port map (
            O => \N__51000\,
            I => \N__50921\
        );

    \I__12263\ : InMux
    port map (
            O => \N__50999\,
            I => \N__50918\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__50996\,
            I => \N__50915\
        );

    \I__12261\ : InMux
    port map (
            O => \N__50995\,
            I => \N__50912\
        );

    \I__12260\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50909\
        );

    \I__12259\ : InMux
    port map (
            O => \N__50993\,
            I => \N__50904\
        );

    \I__12258\ : InMux
    port map (
            O => \N__50992\,
            I => \N__50904\
        );

    \I__12257\ : Span4Mux_h
    port map (
            O => \N__50989\,
            I => \N__50899\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__50986\,
            I => \N__50899\
        );

    \I__12255\ : InMux
    port map (
            O => \N__50985\,
            I => \N__50894\
        );

    \I__12254\ : InMux
    port map (
            O => \N__50984\,
            I => \N__50894\
        );

    \I__12253\ : Span4Mux_v
    port map (
            O => \N__50979\,
            I => \N__50889\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__50974\,
            I => \N__50889\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__50971\,
            I => \N__50882\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__50968\,
            I => \N__50882\
        );

    \I__12249\ : Span4Mux_h
    port map (
            O => \N__50965\,
            I => \N__50882\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__50962\,
            I => \N__50879\
        );

    \I__12247\ : CascadeMux
    port map (
            O => \N__50961\,
            I => \N__50875\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__50958\,
            I => \N__50860\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__50955\,
            I => \N__50860\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__50952\,
            I => \N__50860\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__50949\,
            I => \N__50860\
        );

    \I__12242\ : LocalMux
    port map (
            O => \N__50942\,
            I => \N__50860\
        );

    \I__12241\ : Span4Mux_v
    port map (
            O => \N__50933\,
            I => \N__50860\
        );

    \I__12240\ : CascadeMux
    port map (
            O => \N__50932\,
            I => \N__50857\
        );

    \I__12239\ : CascadeMux
    port map (
            O => \N__50931\,
            I => \N__50853\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__50926\,
            I => \N__50850\
        );

    \I__12237\ : LocalMux
    port map (
            O => \N__50921\,
            I => \N__50845\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__50918\,
            I => \N__50845\
        );

    \I__12235\ : Span4Mux_h
    port map (
            O => \N__50915\,
            I => \N__50834\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__50912\,
            I => \N__50834\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__50909\,
            I => \N__50834\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__50904\,
            I => \N__50834\
        );

    \I__12231\ : Span4Mux_v
    port map (
            O => \N__50899\,
            I => \N__50834\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__50894\,
            I => \N__50825\
        );

    \I__12229\ : Sp12to4
    port map (
            O => \N__50889\,
            I => \N__50825\
        );

    \I__12228\ : Sp12to4
    port map (
            O => \N__50882\,
            I => \N__50825\
        );

    \I__12227\ : Span12Mux_h
    port map (
            O => \N__50879\,
            I => \N__50825\
        );

    \I__12226\ : InMux
    port map (
            O => \N__50878\,
            I => \N__50822\
        );

    \I__12225\ : InMux
    port map (
            O => \N__50875\,
            I => \N__50819\
        );

    \I__12224\ : InMux
    port map (
            O => \N__50874\,
            I => \N__50816\
        );

    \I__12223\ : InMux
    port map (
            O => \N__50873\,
            I => \N__50813\
        );

    \I__12222\ : Span4Mux_v
    port map (
            O => \N__50860\,
            I => \N__50810\
        );

    \I__12221\ : InMux
    port map (
            O => \N__50857\,
            I => \N__50803\
        );

    \I__12220\ : InMux
    port map (
            O => \N__50856\,
            I => \N__50803\
        );

    \I__12219\ : InMux
    port map (
            O => \N__50853\,
            I => \N__50803\
        );

    \I__12218\ : Span4Mux_h
    port map (
            O => \N__50850\,
            I => \N__50800\
        );

    \I__12217\ : Span4Mux_v
    port map (
            O => \N__50845\,
            I => \N__50795\
        );

    \I__12216\ : Span4Mux_v
    port map (
            O => \N__50834\,
            I => \N__50795\
        );

    \I__12215\ : Span12Mux_v
    port map (
            O => \N__50825\,
            I => \N__50792\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__50822\,
            I => \paramsZ0Z_2\
        );

    \I__12213\ : LocalMux
    port map (
            O => \N__50819\,
            I => \paramsZ0Z_2\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__50816\,
            I => \paramsZ0Z_2\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__50813\,
            I => \paramsZ0Z_2\
        );

    \I__12210\ : Odrv4
    port map (
            O => \N__50810\,
            I => \paramsZ0Z_2\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__50803\,
            I => \paramsZ0Z_2\
        );

    \I__12208\ : Odrv4
    port map (
            O => \N__50800\,
            I => \paramsZ0Z_2\
        );

    \I__12207\ : Odrv4
    port map (
            O => \N__50795\,
            I => \paramsZ0Z_2\
        );

    \I__12206\ : Odrv12
    port map (
            O => \N__50792\,
            I => \paramsZ0Z_2\
        );

    \I__12205\ : InMux
    port map (
            O => \N__50773\,
            I => \N__50769\
        );

    \I__12204\ : InMux
    port map (
            O => \N__50772\,
            I => \N__50766\
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__50769\,
            I => \N__50762\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__50766\,
            I => \N__50759\
        );

    \I__12201\ : InMux
    port map (
            O => \N__50765\,
            I => \N__50756\
        );

    \I__12200\ : Span4Mux_v
    port map (
            O => \N__50762\,
            I => \N__50753\
        );

    \I__12199\ : Span4Mux_h
    port map (
            O => \N__50759\,
            I => \N__50749\
        );

    \I__12198\ : LocalMux
    port map (
            O => \N__50756\,
            I => \N__50744\
        );

    \I__12197\ : Span4Mux_v
    port map (
            O => \N__50753\,
            I => \N__50744\
        );

    \I__12196\ : InMux
    port map (
            O => \N__50752\,
            I => \N__50741\
        );

    \I__12195\ : Span4Mux_h
    port map (
            O => \N__50749\,
            I => \N__50737\
        );

    \I__12194\ : Span4Mux_h
    port map (
            O => \N__50744\,
            I => \N__50734\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__50741\,
            I => \N__50731\
        );

    \I__12192\ : InMux
    port map (
            O => \N__50740\,
            I => \N__50728\
        );

    \I__12191\ : Odrv4
    port map (
            O => \N__50737\,
            I => \ALU.r4_RNII2A0LZ0Z_1\
        );

    \I__12190\ : Odrv4
    port map (
            O => \N__50734\,
            I => \ALU.r4_RNII2A0LZ0Z_1\
        );

    \I__12189\ : Odrv4
    port map (
            O => \N__50731\,
            I => \ALU.r4_RNII2A0LZ0Z_1\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__50728\,
            I => \ALU.r4_RNII2A0LZ0Z_1\
        );

    \I__12187\ : CascadeMux
    port map (
            O => \N__50719\,
            I => \N__50716\
        );

    \I__12186\ : InMux
    port map (
            O => \N__50716\,
            I => \N__50713\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__50713\,
            I => \N__50710\
        );

    \I__12184\ : Odrv12
    port map (
            O => \N__50710\,
            I => \ALU.lshift_3\
        );

    \I__12183\ : CascadeMux
    port map (
            O => \N__50707\,
            I => \N__50702\
        );

    \I__12182\ : InMux
    port map (
            O => \N__50706\,
            I => \N__50697\
        );

    \I__12181\ : InMux
    port map (
            O => \N__50705\,
            I => \N__50694\
        );

    \I__12180\ : InMux
    port map (
            O => \N__50702\,
            I => \N__50691\
        );

    \I__12179\ : InMux
    port map (
            O => \N__50701\,
            I => \N__50686\
        );

    \I__12178\ : InMux
    port map (
            O => \N__50700\,
            I => \N__50686\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__50697\,
            I => \N__50683\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__50694\,
            I => \N__50680\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__50691\,
            I => \N__50676\
        );

    \I__12174\ : LocalMux
    port map (
            O => \N__50686\,
            I => \N__50673\
        );

    \I__12173\ : Span4Mux_v
    port map (
            O => \N__50683\,
            I => \N__50670\
        );

    \I__12172\ : Span4Mux_h
    port map (
            O => \N__50680\,
            I => \N__50666\
        );

    \I__12171\ : CascadeMux
    port map (
            O => \N__50679\,
            I => \N__50663\
        );

    \I__12170\ : Span12Mux_h
    port map (
            O => \N__50676\,
            I => \N__50660\
        );

    \I__12169\ : Span4Mux_v
    port map (
            O => \N__50673\,
            I => \N__50657\
        );

    \I__12168\ : Span4Mux_v
    port map (
            O => \N__50670\,
            I => \N__50654\
        );

    \I__12167\ : CascadeMux
    port map (
            O => \N__50669\,
            I => \N__50651\
        );

    \I__12166\ : Span4Mux_v
    port map (
            O => \N__50666\,
            I => \N__50648\
        );

    \I__12165\ : InMux
    port map (
            O => \N__50663\,
            I => \N__50645\
        );

    \I__12164\ : Span12Mux_v
    port map (
            O => \N__50660\,
            I => \N__50642\
        );

    \I__12163\ : Span4Mux_v
    port map (
            O => \N__50657\,
            I => \N__50637\
        );

    \I__12162\ : Span4Mux_v
    port map (
            O => \N__50654\,
            I => \N__50637\
        );

    \I__12161\ : InMux
    port map (
            O => \N__50651\,
            I => \N__50634\
        );

    \I__12160\ : Odrv4
    port map (
            O => \N__50648\,
            I => \ALU.lshift63Z0Z_2\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__50645\,
            I => \ALU.lshift63Z0Z_2\
        );

    \I__12158\ : Odrv12
    port map (
            O => \N__50642\,
            I => \ALU.lshift63Z0Z_2\
        );

    \I__12157\ : Odrv4
    port map (
            O => \N__50637\,
            I => \ALU.lshift63Z0Z_2\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__50634\,
            I => \ALU.lshift63Z0Z_2\
        );

    \I__12155\ : InMux
    port map (
            O => \N__50623\,
            I => \N__50618\
        );

    \I__12154\ : InMux
    port map (
            O => \N__50622\,
            I => \N__50615\
        );

    \I__12153\ : InMux
    port map (
            O => \N__50621\,
            I => \N__50612\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__50618\,
            I => \N__50607\
        );

    \I__12151\ : LocalMux
    port map (
            O => \N__50615\,
            I => \N__50604\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__50612\,
            I => \N__50601\
        );

    \I__12149\ : InMux
    port map (
            O => \N__50611\,
            I => \N__50596\
        );

    \I__12148\ : InMux
    port map (
            O => \N__50610\,
            I => \N__50596\
        );

    \I__12147\ : Span4Mux_v
    port map (
            O => \N__50607\,
            I => \N__50593\
        );

    \I__12146\ : Span4Mux_v
    port map (
            O => \N__50604\,
            I => \N__50590\
        );

    \I__12145\ : Span4Mux_v
    port map (
            O => \N__50601\,
            I => \N__50587\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__50596\,
            I => \N__50584\
        );

    \I__12143\ : Span4Mux_h
    port map (
            O => \N__50593\,
            I => \N__50581\
        );

    \I__12142\ : Span4Mux_h
    port map (
            O => \N__50590\,
            I => \N__50578\
        );

    \I__12141\ : Sp12to4
    port map (
            O => \N__50587\,
            I => \N__50573\
        );

    \I__12140\ : Sp12to4
    port map (
            O => \N__50584\,
            I => \N__50573\
        );

    \I__12139\ : Sp12to4
    port map (
            O => \N__50581\,
            I => \N__50568\
        );

    \I__12138\ : Sp12to4
    port map (
            O => \N__50578\,
            I => \N__50568\
        );

    \I__12137\ : Span12Mux_h
    port map (
            O => \N__50573\,
            I => \N__50565\
        );

    \I__12136\ : Odrv12
    port map (
            O => \N__50568\,
            I => \ALU.r5_RNIAG9A9Z0Z_15\
        );

    \I__12135\ : Odrv12
    port map (
            O => \N__50565\,
            I => \ALU.r5_RNIAG9A9Z0Z_15\
        );

    \I__12134\ : InMux
    port map (
            O => \N__50560\,
            I => \N__50557\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__50557\,
            I => \ALU.r0_12_prm_8_14_s1_c_RNOZ0Z_1\
        );

    \I__12132\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50551\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__50551\,
            I => op_i_0
        );

    \I__12130\ : InMux
    port map (
            O => \N__50548\,
            I => \N__50544\
        );

    \I__12129\ : InMux
    port map (
            O => \N__50547\,
            I => \N__50541\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__50544\,
            I => \N__50538\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__50541\,
            I => \N__50533\
        );

    \I__12126\ : Span4Mux_h
    port map (
            O => \N__50538\,
            I => \N__50533\
        );

    \I__12125\ : Span4Mux_v
    port map (
            O => \N__50533\,
            I => \N__50530\
        );

    \I__12124\ : Span4Mux_h
    port map (
            O => \N__50530\,
            I => \N__50527\
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__50527\,
            I => \ALU.un2_addsub_cry_0_c_RNIJPSHDZ0\
        );

    \I__12122\ : CascadeMux
    port map (
            O => \N__50524\,
            I => \N__50521\
        );

    \I__12121\ : InMux
    port map (
            O => \N__50521\,
            I => \N__50518\
        );

    \I__12120\ : LocalMux
    port map (
            O => \N__50518\,
            I => \N__50515\
        );

    \I__12119\ : Span4Mux_h
    port map (
            O => \N__50515\,
            I => \N__50512\
        );

    \I__12118\ : Odrv4
    port map (
            O => \N__50512\,
            I => \ALU.r0_12_prm_2_1_c_RNOZ0\
        );

    \I__12117\ : InMux
    port map (
            O => \N__50509\,
            I => op_1_cry_1
        );

    \I__12116\ : InMux
    port map (
            O => \N__50506\,
            I => op_1_cry_2
        );

    \I__12115\ : InMux
    port map (
            O => \N__50503\,
            I => op_1_cry_3
        );

    \I__12114\ : CascadeMux
    port map (
            O => \N__50500\,
            I => \N__50494\
        );

    \I__12113\ : CascadeMux
    port map (
            O => \N__50499\,
            I => \N__50490\
        );

    \I__12112\ : CascadeMux
    port map (
            O => \N__50498\,
            I => \N__50486\
        );

    \I__12111\ : InMux
    port map (
            O => \N__50497\,
            I => \N__50467\
        );

    \I__12110\ : InMux
    port map (
            O => \N__50494\,
            I => \N__50467\
        );

    \I__12109\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50467\
        );

    \I__12108\ : InMux
    port map (
            O => \N__50490\,
            I => \N__50467\
        );

    \I__12107\ : InMux
    port map (
            O => \N__50489\,
            I => \N__50467\
        );

    \I__12106\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50467\
        );

    \I__12105\ : InMux
    port map (
            O => \N__50485\,
            I => \N__50467\
        );

    \I__12104\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50467\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__50467\,
            I => \N__50463\
        );

    \I__12102\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50458\
        );

    \I__12101\ : Span4Mux_v
    port map (
            O => \N__50463\,
            I => \N__50455\
        );

    \I__12100\ : InMux
    port map (
            O => \N__50462\,
            I => \N__50450\
        );

    \I__12099\ : InMux
    port map (
            O => \N__50461\,
            I => \N__50450\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__50458\,
            I => \yZ0Z_0\
        );

    \I__12097\ : Odrv4
    port map (
            O => \N__50455\,
            I => \yZ0Z_0\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__50450\,
            I => \yZ0Z_0\
        );

    \I__12095\ : InMux
    port map (
            O => \N__50443\,
            I => \N__50419\
        );

    \I__12094\ : InMux
    port map (
            O => \N__50442\,
            I => \N__50419\
        );

    \I__12093\ : InMux
    port map (
            O => \N__50441\,
            I => \N__50419\
        );

    \I__12092\ : InMux
    port map (
            O => \N__50440\,
            I => \N__50419\
        );

    \I__12091\ : InMux
    port map (
            O => \N__50439\,
            I => \N__50419\
        );

    \I__12090\ : InMux
    port map (
            O => \N__50438\,
            I => \N__50419\
        );

    \I__12089\ : InMux
    port map (
            O => \N__50437\,
            I => \N__50419\
        );

    \I__12088\ : InMux
    port map (
            O => \N__50436\,
            I => \N__50419\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__50419\,
            I => \N__50416\
        );

    \I__12086\ : Span4Mux_v
    port map (
            O => \N__50416\,
            I => \N__50413\
        );

    \I__12085\ : Span4Mux_v
    port map (
            O => \N__50413\,
            I => \N__50408\
        );

    \I__12084\ : InMux
    port map (
            O => \N__50412\,
            I => \N__50403\
        );

    \I__12083\ : InMux
    port map (
            O => \N__50411\,
            I => \N__50403\
        );

    \I__12082\ : Odrv4
    port map (
            O => \N__50408\,
            I => \yZ0Z_1\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__50403\,
            I => \yZ0Z_1\
        );

    \I__12080\ : InMux
    port map (
            O => \N__50398\,
            I => \N__50395\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__50395\,
            I => \N__50392\
        );

    \I__12078\ : Odrv4
    port map (
            O => \N__50392\,
            I => \TXbufferZ0Z_7\
        );

    \I__12077\ : InMux
    port map (
            O => \N__50389\,
            I => \N__50386\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__50386\,
            I => \N__50383\
        );

    \I__12075\ : Span4Mux_v
    port map (
            O => \N__50383\,
            I => \N__50380\
        );

    \I__12074\ : Span4Mux_h
    port map (
            O => \N__50380\,
            I => \N__50377\
        );

    \I__12073\ : Span4Mux_h
    port map (
            O => \N__50377\,
            I => \N__50374\
        );

    \I__12072\ : Odrv4
    port map (
            O => \N__50374\,
            I => \TXbufferZ0Z_1\
        );

    \I__12071\ : InMux
    port map (
            O => \N__50371\,
            I => \N__50368\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__50368\,
            I => \N__50365\
        );

    \I__12069\ : Span4Mux_h
    port map (
            O => \N__50365\,
            I => \N__50362\
        );

    \I__12068\ : Span4Mux_h
    port map (
            O => \N__50362\,
            I => \N__50359\
        );

    \I__12067\ : Span4Mux_h
    port map (
            O => \N__50359\,
            I => \N__50356\
        );

    \I__12066\ : Span4Mux_v
    port map (
            O => \N__50356\,
            I => \N__50353\
        );

    \I__12065\ : Odrv4
    port map (
            O => \N__50353\,
            I => \TXbufferZ0Z_2\
        );

    \I__12064\ : InMux
    port map (
            O => \N__50350\,
            I => \N__50347\
        );

    \I__12063\ : LocalMux
    port map (
            O => \N__50347\,
            I => \FTDI.TXshiftZ0Z_2\
        );

    \I__12062\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50341\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__50341\,
            I => \N__50338\
        );

    \I__12060\ : Sp12to4
    port map (
            O => \N__50338\,
            I => \N__50335\
        );

    \I__12059\ : Span12Mux_s11_v
    port map (
            O => \N__50335\,
            I => \N__50332\
        );

    \I__12058\ : Span12Mux_h
    port map (
            O => \N__50332\,
            I => \N__50329\
        );

    \I__12057\ : Odrv12
    port map (
            O => \N__50329\,
            I => \TXbufferZ0Z_4\
        );

    \I__12056\ : InMux
    port map (
            O => \N__50326\,
            I => \N__50323\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__50323\,
            I => \FTDI.TXshiftZ0Z_4\
        );

    \I__12054\ : InMux
    port map (
            O => \N__50320\,
            I => \N__50317\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__50317\,
            I => \N__50314\
        );

    \I__12052\ : Span12Mux_h
    port map (
            O => \N__50314\,
            I => \N__50311\
        );

    \I__12051\ : Span12Mux_v
    port map (
            O => \N__50311\,
            I => \N__50308\
        );

    \I__12050\ : Span12Mux_h
    port map (
            O => \N__50308\,
            I => \N__50305\
        );

    \I__12049\ : Odrv12
    port map (
            O => \N__50305\,
            I => \TXbufferZ0Z_3\
        );

    \I__12048\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50299\
        );

    \I__12047\ : LocalMux
    port map (
            O => \N__50299\,
            I => \FTDI.TXshiftZ0Z_3\
        );

    \I__12046\ : InMux
    port map (
            O => \N__50296\,
            I => \N__50293\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__50293\,
            I => \N__50290\
        );

    \I__12044\ : Odrv4
    port map (
            O => \N__50290\,
            I => \FTDI.TXshiftZ0Z_7\
        );

    \I__12043\ : InMux
    port map (
            O => \N__50287\,
            I => \N__50284\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__50284\,
            I => \N__50281\
        );

    \I__12041\ : Span12Mux_v
    port map (
            O => \N__50281\,
            I => \N__50278\
        );

    \I__12040\ : Span12Mux_h
    port map (
            O => \N__50278\,
            I => \N__50275\
        );

    \I__12039\ : Odrv12
    port map (
            O => \N__50275\,
            I => \TXbufferZ0Z_6\
        );

    \I__12038\ : InMux
    port map (
            O => \N__50272\,
            I => \N__50269\
        );

    \I__12037\ : LocalMux
    port map (
            O => \N__50269\,
            I => \FTDI.TXshiftZ0Z_6\
        );

    \I__12036\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50263\
        );

    \I__12035\ : LocalMux
    port map (
            O => \N__50263\,
            I => \N__50260\
        );

    \I__12034\ : Span4Mux_v
    port map (
            O => \N__50260\,
            I => \N__50257\
        );

    \I__12033\ : Span4Mux_h
    port map (
            O => \N__50257\,
            I => \N__50254\
        );

    \I__12032\ : Span4Mux_h
    port map (
            O => \N__50254\,
            I => \N__50251\
        );

    \I__12031\ : Odrv4
    port map (
            O => \N__50251\,
            I => \TXbufferZ0Z_5\
        );

    \I__12030\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50245\
        );

    \I__12029\ : LocalMux
    port map (
            O => \N__50245\,
            I => \FTDI.TXshiftZ0Z_5\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50242\,
            I => \N__50239\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__50239\,
            I => \ALU.r0_12_prm_1_3_c_RNOZ0\
        );

    \I__12026\ : CascadeMux
    port map (
            O => \N__50236\,
            I => \N__50233\
        );

    \I__12025\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50229\
        );

    \I__12024\ : InMux
    port map (
            O => \N__50232\,
            I => \N__50226\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__50229\,
            I => \N__50223\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__50226\,
            I => \N__50220\
        );

    \I__12021\ : Span4Mux_v
    port map (
            O => \N__50223\,
            I => \N__50217\
        );

    \I__12020\ : Span4Mux_v
    port map (
            O => \N__50220\,
            I => \N__50214\
        );

    \I__12019\ : Span4Mux_h
    port map (
            O => \N__50217\,
            I => \N__50211\
        );

    \I__12018\ : Span4Mux_h
    port map (
            O => \N__50214\,
            I => \N__50208\
        );

    \I__12017\ : Odrv4
    port map (
            O => \N__50211\,
            I => \ALU.un9_addsub_cry_2_c_RNIOR8AJZ0\
        );

    \I__12016\ : Odrv4
    port map (
            O => \N__50208\,
            I => \ALU.un9_addsub_cry_2_c_RNIOR8AJZ0\
        );

    \I__12015\ : InMux
    port map (
            O => \N__50203\,
            I => \ALU.r0_12_3\
        );

    \I__12014\ : InMux
    port map (
            O => \N__50200\,
            I => \N__50196\
        );

    \I__12013\ : InMux
    port map (
            O => \N__50199\,
            I => \N__50193\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__50196\,
            I => \N__50189\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__50193\,
            I => \N__50185\
        );

    \I__12010\ : InMux
    port map (
            O => \N__50192\,
            I => \N__50182\
        );

    \I__12009\ : Span4Mux_h
    port map (
            O => \N__50189\,
            I => \N__50179\
        );

    \I__12008\ : InMux
    port map (
            O => \N__50188\,
            I => \N__50176\
        );

    \I__12007\ : Span4Mux_v
    port map (
            O => \N__50185\,
            I => \N__50172\
        );

    \I__12006\ : LocalMux
    port map (
            O => \N__50182\,
            I => \N__50168\
        );

    \I__12005\ : Span4Mux_h
    port map (
            O => \N__50179\,
            I => \N__50163\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__50176\,
            I => \N__50163\
        );

    \I__12003\ : InMux
    port map (
            O => \N__50175\,
            I => \N__50160\
        );

    \I__12002\ : Span4Mux_h
    port map (
            O => \N__50172\,
            I => \N__50156\
        );

    \I__12001\ : InMux
    port map (
            O => \N__50171\,
            I => \N__50153\
        );

    \I__12000\ : Span4Mux_h
    port map (
            O => \N__50168\,
            I => \N__50150\
        );

    \I__11999\ : Span4Mux_v
    port map (
            O => \N__50163\,
            I => \N__50145\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__50160\,
            I => \N__50145\
        );

    \I__11997\ : InMux
    port map (
            O => \N__50159\,
            I => \N__50142\
        );

    \I__11996\ : Span4Mux_h
    port map (
            O => \N__50156\,
            I => \N__50137\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__50153\,
            I => \N__50137\
        );

    \I__11994\ : Span4Mux_h
    port map (
            O => \N__50150\,
            I => \N__50129\
        );

    \I__11993\ : Span4Mux_h
    port map (
            O => \N__50145\,
            I => \N__50129\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__50142\,
            I => \N__50129\
        );

    \I__11991\ : Span4Mux_h
    port map (
            O => \N__50137\,
            I => \N__50126\
        );

    \I__11990\ : InMux
    port map (
            O => \N__50136\,
            I => \N__50123\
        );

    \I__11989\ : Span4Mux_h
    port map (
            O => \N__50129\,
            I => \N__50120\
        );

    \I__11988\ : Sp12to4
    port map (
            O => \N__50126\,
            I => \N__50115\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__50123\,
            I => \N__50115\
        );

    \I__11986\ : Odrv4
    port map (
            O => \N__50120\,
            I => \ALU.r0_12_3_THRU_CO\
        );

    \I__11985\ : Odrv12
    port map (
            O => \N__50115\,
            I => \ALU.r0_12_3_THRU_CO\
        );

    \I__11984\ : CascadeMux
    port map (
            O => \N__50110\,
            I => \N__50107\
        );

    \I__11983\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50104\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__50104\,
            I => \N__50100\
        );

    \I__11981\ : InMux
    port map (
            O => \N__50103\,
            I => \N__50097\
        );

    \I__11980\ : Span4Mux_h
    port map (
            O => \N__50100\,
            I => \N__50094\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__50097\,
            I => \N__50091\
        );

    \I__11978\ : Span4Mux_h
    port map (
            O => \N__50094\,
            I => \N__50088\
        );

    \I__11977\ : Span4Mux_h
    port map (
            O => \N__50091\,
            I => \N__50085\
        );

    \I__11976\ : Span4Mux_h
    port map (
            O => \N__50088\,
            I => \N__50082\
        );

    \I__11975\ : Span4Mux_h
    port map (
            O => \N__50085\,
            I => \N__50079\
        );

    \I__11974\ : Odrv4
    port map (
            O => \N__50082\,
            I => \ALU.un2_addsub_cry_2_c_RNI3K9SGZ0\
        );

    \I__11973\ : Odrv4
    port map (
            O => \N__50079\,
            I => \ALU.un2_addsub_cry_2_c_RNI3K9SGZ0\
        );

    \I__11972\ : InMux
    port map (
            O => \N__50074\,
            I => \N__50071\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__50071\,
            I => \ALU.r0_12_prm_2_3_c_RNOZ0\
        );

    \I__11970\ : InMux
    port map (
            O => \N__50068\,
            I => \N__50065\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__50065\,
            I => \ALU.r0_12_prm_3_3_c_RNOZ0\
        );

    \I__11968\ : InMux
    port map (
            O => \N__50062\,
            I => \N__50056\
        );

    \I__11967\ : InMux
    port map (
            O => \N__50061\,
            I => \N__50056\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__50056\,
            I => \N__50053\
        );

    \I__11965\ : Span4Mux_h
    port map (
            O => \N__50053\,
            I => \N__50049\
        );

    \I__11964\ : InMux
    port map (
            O => \N__50052\,
            I => \N__50046\
        );

    \I__11963\ : Span4Mux_h
    port map (
            O => \N__50049\,
            I => \N__50041\
        );

    \I__11962\ : LocalMux
    port map (
            O => \N__50046\,
            I => \N__50041\
        );

    \I__11961\ : Span4Mux_h
    port map (
            O => \N__50041\,
            I => \N__50038\
        );

    \I__11960\ : Odrv4
    port map (
            O => \N__50038\,
            I => \ALU.madd_axb_2\
        );

    \I__11959\ : CascadeMux
    port map (
            O => \N__50035\,
            I => \N__50032\
        );

    \I__11958\ : InMux
    port map (
            O => \N__50032\,
            I => \N__50026\
        );

    \I__11957\ : InMux
    port map (
            O => \N__50031\,
            I => \N__50026\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__50026\,
            I => \N__50023\
        );

    \I__11955\ : Span4Mux_h
    port map (
            O => \N__50023\,
            I => \N__50020\
        );

    \I__11954\ : Span4Mux_h
    port map (
            O => \N__50020\,
            I => \N__50017\
        );

    \I__11953\ : Span4Mux_h
    port map (
            O => \N__50017\,
            I => \N__50014\
        );

    \I__11952\ : Odrv4
    port map (
            O => \N__50014\,
            I => \ALU.madd_cry_1_THRU_CO\
        );

    \I__11951\ : CascadeMux
    port map (
            O => \N__50011\,
            I => \N__50008\
        );

    \I__11950\ : InMux
    port map (
            O => \N__50008\,
            I => \N__50005\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__50005\,
            I => \ALU.mult_3\
        );

    \I__11948\ : InMux
    port map (
            O => \N__50002\,
            I => \N__49999\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__49999\,
            I => \N__49996\
        );

    \I__11946\ : Span12Mux_v
    port map (
            O => \N__49996\,
            I => \N__49993\
        );

    \I__11945\ : Span12Mux_h
    port map (
            O => \N__49993\,
            I => \N__49990\
        );

    \I__11944\ : Odrv12
    port map (
            O => \N__49990\,
            I => \TXbuffer_RNO_1Z0Z_7\
        );

    \I__11943\ : InMux
    port map (
            O => \N__49987\,
            I => \N__49984\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__49984\,
            I => \N__49981\
        );

    \I__11941\ : Odrv12
    port map (
            O => \N__49981\,
            I => \TXbuffer_RNO_0Z0Z_7\
        );

    \I__11940\ : CascadeMux
    port map (
            O => \N__49978\,
            I => \N__49975\
        );

    \I__11939\ : InMux
    port map (
            O => \N__49975\,
            I => \N__49971\
        );

    \I__11938\ : CascadeMux
    port map (
            O => \N__49974\,
            I => \N__49964\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__49971\,
            I => \N__49961\
        );

    \I__11936\ : InMux
    port map (
            O => \N__49970\,
            I => \N__49958\
        );

    \I__11935\ : InMux
    port map (
            O => \N__49969\,
            I => \N__49955\
        );

    \I__11934\ : InMux
    port map (
            O => \N__49968\,
            I => \N__49952\
        );

    \I__11933\ : CascadeMux
    port map (
            O => \N__49967\,
            I => \N__49949\
        );

    \I__11932\ : InMux
    port map (
            O => \N__49964\,
            I => \N__49946\
        );

    \I__11931\ : Span4Mux_v
    port map (
            O => \N__49961\,
            I => \N__49941\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__49958\,
            I => \N__49941\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__49955\,
            I => \N__49933\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__49952\,
            I => \N__49929\
        );

    \I__11927\ : InMux
    port map (
            O => \N__49949\,
            I => \N__49926\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__49946\,
            I => \N__49922\
        );

    \I__11925\ : Span4Mux_v
    port map (
            O => \N__49941\,
            I => \N__49919\
        );

    \I__11924\ : InMux
    port map (
            O => \N__49940\,
            I => \N__49916\
        );

    \I__11923\ : InMux
    port map (
            O => \N__49939\,
            I => \N__49911\
        );

    \I__11922\ : InMux
    port map (
            O => \N__49938\,
            I => \N__49911\
        );

    \I__11921\ : InMux
    port map (
            O => \N__49937\,
            I => \N__49906\
        );

    \I__11920\ : InMux
    port map (
            O => \N__49936\,
            I => \N__49906\
        );

    \I__11919\ : Span4Mux_v
    port map (
            O => \N__49933\,
            I => \N__49903\
        );

    \I__11918\ : InMux
    port map (
            O => \N__49932\,
            I => \N__49899\
        );

    \I__11917\ : Span4Mux_v
    port map (
            O => \N__49929\,
            I => \N__49896\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__49926\,
            I => \N__49893\
        );

    \I__11915\ : InMux
    port map (
            O => \N__49925\,
            I => \N__49890\
        );

    \I__11914\ : Span12Mux_h
    port map (
            O => \N__49922\,
            I => \N__49881\
        );

    \I__11913\ : Sp12to4
    port map (
            O => \N__49919\,
            I => \N__49881\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__49916\,
            I => \N__49881\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__49911\,
            I => \N__49874\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__49906\,
            I => \N__49874\
        );

    \I__11909\ : Span4Mux_h
    port map (
            O => \N__49903\,
            I => \N__49874\
        );

    \I__11908\ : InMux
    port map (
            O => \N__49902\,
            I => \N__49871\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__49899\,
            I => \N__49868\
        );

    \I__11906\ : Span4Mux_h
    port map (
            O => \N__49896\,
            I => \N__49865\
        );

    \I__11905\ : Span4Mux_h
    port map (
            O => \N__49893\,
            I => \N__49860\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__49890\,
            I => \N__49860\
        );

    \I__11903\ : InMux
    port map (
            O => \N__49889\,
            I => \N__49857\
        );

    \I__11902\ : InMux
    port map (
            O => \N__49888\,
            I => \N__49854\
        );

    \I__11901\ : Span12Mux_h
    port map (
            O => \N__49881\,
            I => \N__49850\
        );

    \I__11900\ : Span4Mux_v
    port map (
            O => \N__49874\,
            I => \N__49847\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__49871\,
            I => \N__49842\
        );

    \I__11898\ : Span4Mux_v
    port map (
            O => \N__49868\,
            I => \N__49842\
        );

    \I__11897\ : Span4Mux_v
    port map (
            O => \N__49865\,
            I => \N__49837\
        );

    \I__11896\ : Span4Mux_h
    port map (
            O => \N__49860\,
            I => \N__49837\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__49857\,
            I => \N__49832\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__49854\,
            I => \N__49832\
        );

    \I__11893\ : InMux
    port map (
            O => \N__49853\,
            I => \N__49829\
        );

    \I__11892\ : Odrv12
    port map (
            O => \N__49850\,
            I => \clkdivZ0Z_4\
        );

    \I__11891\ : Odrv4
    port map (
            O => \N__49847\,
            I => \clkdivZ0Z_4\
        );

    \I__11890\ : Odrv4
    port map (
            O => \N__49842\,
            I => \clkdivZ0Z_4\
        );

    \I__11889\ : Odrv4
    port map (
            O => \N__49837\,
            I => \clkdivZ0Z_4\
        );

    \I__11888\ : Odrv4
    port map (
            O => \N__49832\,
            I => \clkdivZ0Z_4\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__49829\,
            I => \clkdivZ0Z_4\
        );

    \I__11886\ : InMux
    port map (
            O => \N__49816\,
            I => \N__49813\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__49813\,
            I => \N__49810\
        );

    \I__11884\ : Odrv12
    port map (
            O => \N__49810\,
            I => \TXbuffer_18_15_ns_1_7\
        );

    \I__11883\ : CascadeMux
    port map (
            O => \N__49807\,
            I => \N__49804\
        );

    \I__11882\ : InMux
    port map (
            O => \N__49804\,
            I => \N__49797\
        );

    \I__11881\ : CascadeMux
    port map (
            O => \N__49803\,
            I => \N__49792\
        );

    \I__11880\ : CascadeMux
    port map (
            O => \N__49802\,
            I => \N__49788\
        );

    \I__11879\ : CascadeMux
    port map (
            O => \N__49801\,
            I => \N__49784\
        );

    \I__11878\ : CascadeMux
    port map (
            O => \N__49800\,
            I => \N__49781\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__49797\,
            I => \N__49778\
        );

    \I__11876\ : InMux
    port map (
            O => \N__49796\,
            I => \N__49761\
        );

    \I__11875\ : InMux
    port map (
            O => \N__49795\,
            I => \N__49761\
        );

    \I__11874\ : InMux
    port map (
            O => \N__49792\,
            I => \N__49761\
        );

    \I__11873\ : InMux
    port map (
            O => \N__49791\,
            I => \N__49761\
        );

    \I__11872\ : InMux
    port map (
            O => \N__49788\,
            I => \N__49761\
        );

    \I__11871\ : InMux
    port map (
            O => \N__49787\,
            I => \N__49761\
        );

    \I__11870\ : InMux
    port map (
            O => \N__49784\,
            I => \N__49761\
        );

    \I__11869\ : InMux
    port map (
            O => \N__49781\,
            I => \N__49761\
        );

    \I__11868\ : Odrv4
    port map (
            O => \N__49778\,
            I => \yZ0Z_2\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__49761\,
            I => \yZ0Z_2\
        );

    \I__11866\ : CEMux
    port map (
            O => \N__49756\,
            I => \N__49753\
        );

    \I__11865\ : LocalMux
    port map (
            O => \N__49753\,
            I => \N__49750\
        );

    \I__11864\ : Span4Mux_v
    port map (
            O => \N__49750\,
            I => \N__49747\
        );

    \I__11863\ : Span4Mux_h
    port map (
            O => \N__49747\,
            I => \N__49743\
        );

    \I__11862\ : CEMux
    port map (
            O => \N__49746\,
            I => \N__49740\
        );

    \I__11861\ : Span4Mux_h
    port map (
            O => \N__49743\,
            I => \N__49734\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__49740\,
            I => \N__49734\
        );

    \I__11859\ : CEMux
    port map (
            O => \N__49739\,
            I => \N__49727\
        );

    \I__11858\ : Span4Mux_v
    port map (
            O => \N__49734\,
            I => \N__49723\
        );

    \I__11857\ : CEMux
    port map (
            O => \N__49733\,
            I => \N__49720\
        );

    \I__11856\ : CEMux
    port map (
            O => \N__49732\,
            I => \N__49713\
        );

    \I__11855\ : CEMux
    port map (
            O => \N__49731\,
            I => \N__49710\
        );

    \I__11854\ : CEMux
    port map (
            O => \N__49730\,
            I => \N__49707\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__49727\,
            I => \N__49704\
        );

    \I__11852\ : CEMux
    port map (
            O => \N__49726\,
            I => \N__49701\
        );

    \I__11851\ : Span4Mux_h
    port map (
            O => \N__49723\,
            I => \N__49698\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__49720\,
            I => \N__49695\
        );

    \I__11849\ : CEMux
    port map (
            O => \N__49719\,
            I => \N__49692\
        );

    \I__11848\ : CEMux
    port map (
            O => \N__49718\,
            I => \N__49689\
        );

    \I__11847\ : CEMux
    port map (
            O => \N__49717\,
            I => \N__49686\
        );

    \I__11846\ : CEMux
    port map (
            O => \N__49716\,
            I => \N__49682\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__49713\,
            I => \N__49679\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__49710\,
            I => \N__49676\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__49707\,
            I => \N__49673\
        );

    \I__11842\ : Span4Mux_v
    port map (
            O => \N__49704\,
            I => \N__49670\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__49701\,
            I => \N__49667\
        );

    \I__11840\ : Span4Mux_s0_h
    port map (
            O => \N__49698\,
            I => \N__49664\
        );

    \I__11839\ : Span4Mux_h
    port map (
            O => \N__49695\,
            I => \N__49661\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__49692\,
            I => \N__49658\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__49689\,
            I => \N__49655\
        );

    \I__11836\ : LocalMux
    port map (
            O => \N__49686\,
            I => \N__49652\
        );

    \I__11835\ : CEMux
    port map (
            O => \N__49685\,
            I => \N__49649\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__49682\,
            I => \N__49646\
        );

    \I__11833\ : Span4Mux_v
    port map (
            O => \N__49679\,
            I => \N__49643\
        );

    \I__11832\ : Span4Mux_v
    port map (
            O => \N__49676\,
            I => \N__49640\
        );

    \I__11831\ : Span4Mux_h
    port map (
            O => \N__49673\,
            I => \N__49637\
        );

    \I__11830\ : Span4Mux_s3_h
    port map (
            O => \N__49670\,
            I => \N__49634\
        );

    \I__11829\ : Span4Mux_h
    port map (
            O => \N__49667\,
            I => \N__49631\
        );

    \I__11828\ : Span4Mux_v
    port map (
            O => \N__49664\,
            I => \N__49626\
        );

    \I__11827\ : Span4Mux_s0_h
    port map (
            O => \N__49661\,
            I => \N__49626\
        );

    \I__11826\ : Span4Mux_v
    port map (
            O => \N__49658\,
            I => \N__49619\
        );

    \I__11825\ : Span4Mux_v
    port map (
            O => \N__49655\,
            I => \N__49619\
        );

    \I__11824\ : Span4Mux_h
    port map (
            O => \N__49652\,
            I => \N__49619\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__49649\,
            I => \N__49616\
        );

    \I__11822\ : Span4Mux_v
    port map (
            O => \N__49646\,
            I => \N__49609\
        );

    \I__11821\ : Span4Mux_h
    port map (
            O => \N__49643\,
            I => \N__49609\
        );

    \I__11820\ : Span4Mux_h
    port map (
            O => \N__49640\,
            I => \N__49609\
        );

    \I__11819\ : Span4Mux_h
    port map (
            O => \N__49637\,
            I => \N__49606\
        );

    \I__11818\ : Span4Mux_h
    port map (
            O => \N__49634\,
            I => \N__49603\
        );

    \I__11817\ : Span4Mux_h
    port map (
            O => \N__49631\,
            I => \N__49600\
        );

    \I__11816\ : Span4Mux_v
    port map (
            O => \N__49626\,
            I => \N__49597\
        );

    \I__11815\ : Span4Mux_h
    port map (
            O => \N__49619\,
            I => \N__49594\
        );

    \I__11814\ : Span4Mux_h
    port map (
            O => \N__49616\,
            I => \N__49591\
        );

    \I__11813\ : Span4Mux_h
    port map (
            O => \N__49609\,
            I => \N__49588\
        );

    \I__11812\ : Span4Mux_v
    port map (
            O => \N__49606\,
            I => \N__49583\
        );

    \I__11811\ : Span4Mux_h
    port map (
            O => \N__49603\,
            I => \N__49583\
        );

    \I__11810\ : Sp12to4
    port map (
            O => \N__49600\,
            I => \N__49580\
        );

    \I__11809\ : Sp12to4
    port map (
            O => \N__49597\,
            I => \N__49577\
        );

    \I__11808\ : Span4Mux_h
    port map (
            O => \N__49594\,
            I => \N__49574\
        );

    \I__11807\ : Span4Mux_h
    port map (
            O => \N__49591\,
            I => \N__49569\
        );

    \I__11806\ : Span4Mux_h
    port map (
            O => \N__49588\,
            I => \N__49569\
        );

    \I__11805\ : Span4Mux_h
    port map (
            O => \N__49583\,
            I => \N__49566\
        );

    \I__11804\ : Span12Mux_v
    port map (
            O => \N__49580\,
            I => \N__49561\
        );

    \I__11803\ : Span12Mux_s11_h
    port map (
            O => \N__49577\,
            I => \N__49561\
        );

    \I__11802\ : Span4Mux_v
    port map (
            O => \N__49574\,
            I => \N__49558\
        );

    \I__11801\ : Odrv4
    port map (
            O => \N__49569\,
            I => \ALU.un1_yindexZ0Z_8\
        );

    \I__11800\ : Odrv4
    port map (
            O => \N__49566\,
            I => \ALU.un1_yindexZ0Z_8\
        );

    \I__11799\ : Odrv12
    port map (
            O => \N__49561\,
            I => \ALU.un1_yindexZ0Z_8\
        );

    \I__11798\ : Odrv4
    port map (
            O => \N__49558\,
            I => \ALU.un1_yindexZ0Z_8\
        );

    \I__11797\ : CascadeMux
    port map (
            O => \N__49549\,
            I => \N__49546\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49546\,
            I => \N__49542\
        );

    \I__11795\ : InMux
    port map (
            O => \N__49545\,
            I => \N__49539\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__49542\,
            I => \ALU.rshift_3\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__49539\,
            I => \ALU.rshift_3\
        );

    \I__11792\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49531\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__49531\,
            I => \N__49528\
        );

    \I__11790\ : Span4Mux_h
    port map (
            O => \N__49528\,
            I => \N__49525\
        );

    \I__11789\ : Odrv4
    port map (
            O => \N__49525\,
            I => \ALU.r0_12_prm_8_3_c_RNOZ0\
        );

    \I__11788\ : InMux
    port map (
            O => \N__49522\,
            I => \N__49519\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__49519\,
            I => \ALU.r0_12_prm_7_3_c_RNOZ0\
        );

    \I__11786\ : CascadeMux
    port map (
            O => \N__49516\,
            I => \N__49513\
        );

    \I__11785\ : InMux
    port map (
            O => \N__49513\,
            I => \N__49509\
        );

    \I__11784\ : InMux
    port map (
            O => \N__49512\,
            I => \N__49506\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__49509\,
            I => \N__49501\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49506\,
            I => \N__49501\
        );

    \I__11781\ : Span4Mux_v
    port map (
            O => \N__49501\,
            I => \N__49498\
        );

    \I__11780\ : Span4Mux_h
    port map (
            O => \N__49498\,
            I => \N__49495\
        );

    \I__11779\ : Odrv4
    port map (
            O => \N__49495\,
            I => \ALU.a3_b_3\
        );

    \I__11778\ : InMux
    port map (
            O => \N__49492\,
            I => \N__49489\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__49489\,
            I => \N__49486\
        );

    \I__11776\ : Span12Mux_h
    port map (
            O => \N__49486\,
            I => \N__49483\
        );

    \I__11775\ : Odrv12
    port map (
            O => \N__49483\,
            I => \ALU.un14_log_0_i_3\
        );

    \I__11774\ : CascadeMux
    port map (
            O => \N__49480\,
            I => \N__49477\
        );

    \I__11773\ : InMux
    port map (
            O => \N__49477\,
            I => \N__49474\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__49474\,
            I => \N__49471\
        );

    \I__11771\ : Span12Mux_h
    port map (
            O => \N__49471\,
            I => \N__49468\
        );

    \I__11770\ : Odrv12
    port map (
            O => \N__49468\,
            I => \ALU.r0_12_prm_6_3_c_RNOZ0\
        );

    \I__11769\ : InMux
    port map (
            O => \N__49465\,
            I => \N__49462\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__49462\,
            I => \ALU.r0_12_prm_5_3_c_RNOZ0\
        );

    \I__11767\ : CascadeMux
    port map (
            O => \N__49459\,
            I => \N__49456\
        );

    \I__11766\ : InMux
    port map (
            O => \N__49456\,
            I => \N__49453\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__49453\,
            I => \N__49450\
        );

    \I__11764\ : Span4Mux_h
    port map (
            O => \N__49450\,
            I => \N__49447\
        );

    \I__11763\ : Odrv4
    port map (
            O => \N__49447\,
            I => \ALU.r0_12_prm_5_3_c_RNOZ0Z_0\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49444\,
            I => \N__49441\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__49441\,
            I => \N__49438\
        );

    \I__11760\ : Span4Mux_v
    port map (
            O => \N__49438\,
            I => \N__49435\
        );

    \I__11759\ : Span4Mux_v
    port map (
            O => \N__49435\,
            I => \N__49432\
        );

    \I__11758\ : Span4Mux_h
    port map (
            O => \N__49432\,
            I => \N__49429\
        );

    \I__11757\ : Odrv4
    port map (
            O => \N__49429\,
            I => \ALU.r4_RNIUH636Z0Z_3\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49426\,
            I => \N__49420\
        );

    \I__11755\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49413\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49424\,
            I => \N__49409\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49405\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49402\
        );

    \I__11751\ : InMux
    port map (
            O => \N__49419\,
            I => \N__49399\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49418\,
            I => \N__49394\
        );

    \I__11749\ : InMux
    port map (
            O => \N__49417\,
            I => \N__49390\
        );

    \I__11748\ : InMux
    port map (
            O => \N__49416\,
            I => \N__49387\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__49413\,
            I => \N__49384\
        );

    \I__11746\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49381\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__49409\,
            I => \N__49378\
        );

    \I__11744\ : InMux
    port map (
            O => \N__49408\,
            I => \N__49375\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__49405\,
            I => \N__49372\
        );

    \I__11742\ : Span4Mux_h
    port map (
            O => \N__49402\,
            I => \N__49367\
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__49399\,
            I => \N__49367\
        );

    \I__11740\ : InMux
    port map (
            O => \N__49398\,
            I => \N__49357\
        );

    \I__11739\ : InMux
    port map (
            O => \N__49397\,
            I => \N__49354\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__49394\,
            I => \N__49345\
        );

    \I__11737\ : InMux
    port map (
            O => \N__49393\,
            I => \N__49342\
        );

    \I__11736\ : LocalMux
    port map (
            O => \N__49390\,
            I => \N__49338\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__49387\,
            I => \N__49335\
        );

    \I__11734\ : Span4Mux_v
    port map (
            O => \N__49384\,
            I => \N__49326\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__49381\,
            I => \N__49326\
        );

    \I__11732\ : Span4Mux_h
    port map (
            O => \N__49378\,
            I => \N__49326\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__49375\,
            I => \N__49326\
        );

    \I__11730\ : Span4Mux_h
    port map (
            O => \N__49372\,
            I => \N__49319\
        );

    \I__11729\ : Span4Mux_v
    port map (
            O => \N__49367\,
            I => \N__49319\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49316\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49365\,
            I => \N__49309\
        );

    \I__11726\ : InMux
    port map (
            O => \N__49364\,
            I => \N__49309\
        );

    \I__11725\ : InMux
    port map (
            O => \N__49363\,
            I => \N__49309\
        );

    \I__11724\ : InMux
    port map (
            O => \N__49362\,
            I => \N__49306\
        );

    \I__11723\ : InMux
    port map (
            O => \N__49361\,
            I => \N__49303\
        );

    \I__11722\ : InMux
    port map (
            O => \N__49360\,
            I => \N__49300\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__49357\,
            I => \N__49297\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__49354\,
            I => \N__49294\
        );

    \I__11719\ : InMux
    port map (
            O => \N__49353\,
            I => \N__49289\
        );

    \I__11718\ : InMux
    port map (
            O => \N__49352\,
            I => \N__49289\
        );

    \I__11717\ : InMux
    port map (
            O => \N__49351\,
            I => \N__49283\
        );

    \I__11716\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49283\
        );

    \I__11715\ : InMux
    port map (
            O => \N__49349\,
            I => \N__49278\
        );

    \I__11714\ : InMux
    port map (
            O => \N__49348\,
            I => \N__49278\
        );

    \I__11713\ : Span4Mux_v
    port map (
            O => \N__49345\,
            I => \N__49274\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__49342\,
            I => \N__49271\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49341\,
            I => \N__49268\
        );

    \I__11710\ : Span4Mux_v
    port map (
            O => \N__49338\,
            I => \N__49265\
        );

    \I__11709\ : Span4Mux_h
    port map (
            O => \N__49335\,
            I => \N__49260\
        );

    \I__11708\ : Span4Mux_v
    port map (
            O => \N__49326\,
            I => \N__49260\
        );

    \I__11707\ : InMux
    port map (
            O => \N__49325\,
            I => \N__49255\
        );

    \I__11706\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49255\
        );

    \I__11705\ : Span4Mux_h
    port map (
            O => \N__49319\,
            I => \N__49250\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__49316\,
            I => \N__49247\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__49309\,
            I => \N__49242\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__49306\,
            I => \N__49242\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__49303\,
            I => \N__49239\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__49300\,
            I => \N__49227\
        );

    \I__11699\ : Span4Mux_s0_v
    port map (
            O => \N__49297\,
            I => \N__49227\
        );

    \I__11698\ : Span4Mux_v
    port map (
            O => \N__49294\,
            I => \N__49227\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__49289\,
            I => \N__49227\
        );

    \I__11696\ : InMux
    port map (
            O => \N__49288\,
            I => \N__49224\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__49283\,
            I => \N__49219\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__49278\,
            I => \N__49219\
        );

    \I__11693\ : InMux
    port map (
            O => \N__49277\,
            I => \N__49216\
        );

    \I__11692\ : Span4Mux_h
    port map (
            O => \N__49274\,
            I => \N__49213\
        );

    \I__11691\ : Span12Mux_v
    port map (
            O => \N__49271\,
            I => \N__49202\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__49268\,
            I => \N__49202\
        );

    \I__11689\ : Sp12to4
    port map (
            O => \N__49265\,
            I => \N__49202\
        );

    \I__11688\ : Sp12to4
    port map (
            O => \N__49260\,
            I => \N__49202\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__49255\,
            I => \N__49202\
        );

    \I__11686\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49197\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49197\
        );

    \I__11684\ : Span4Mux_v
    port map (
            O => \N__49250\,
            I => \N__49192\
        );

    \I__11683\ : Span4Mux_h
    port map (
            O => \N__49247\,
            I => \N__49192\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__49242\,
            I => \N__49187\
        );

    \I__11681\ : Span4Mux_s3_v
    port map (
            O => \N__49239\,
            I => \N__49187\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49238\,
            I => \N__49184\
        );

    \I__11679\ : InMux
    port map (
            O => \N__49237\,
            I => \N__49179\
        );

    \I__11678\ : InMux
    port map (
            O => \N__49236\,
            I => \N__49179\
        );

    \I__11677\ : Span4Mux_h
    port map (
            O => \N__49227\,
            I => \N__49170\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__49224\,
            I => \N__49170\
        );

    \I__11675\ : Span4Mux_h
    port map (
            O => \N__49219\,
            I => \N__49170\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__49216\,
            I => \N__49170\
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__49213\,
            I => \ALU.a_3\
        );

    \I__11672\ : Odrv12
    port map (
            O => \N__49202\,
            I => \ALU.a_3\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__49197\,
            I => \ALU.a_3\
        );

    \I__11670\ : Odrv4
    port map (
            O => \N__49192\,
            I => \ALU.a_3\
        );

    \I__11669\ : Odrv4
    port map (
            O => \N__49187\,
            I => \ALU.a_3\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__49184\,
            I => \ALU.a_3\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__49179\,
            I => \ALU.a_3\
        );

    \I__11666\ : Odrv4
    port map (
            O => \N__49170\,
            I => \ALU.a_3\
        );

    \I__11665\ : CascadeMux
    port map (
            O => \N__49153\,
            I => \N__49150\
        );

    \I__11664\ : InMux
    port map (
            O => \N__49150\,
            I => \N__49147\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__49147\,
            I => \N__49144\
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__49144\,
            I => \ALU.a_i_3\
        );

    \I__11661\ : InMux
    port map (
            O => \N__49141\,
            I => \N__49137\
        );

    \I__11660\ : InMux
    port map (
            O => \N__49140\,
            I => \N__49133\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__49137\,
            I => \N__49129\
        );

    \I__11658\ : InMux
    port map (
            O => \N__49136\,
            I => \N__49126\
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__49133\,
            I => \N__49123\
        );

    \I__11656\ : InMux
    port map (
            O => \N__49132\,
            I => \N__49120\
        );

    \I__11655\ : Span4Mux_h
    port map (
            O => \N__49129\,
            I => \N__49115\
        );

    \I__11654\ : LocalMux
    port map (
            O => \N__49126\,
            I => \N__49115\
        );

    \I__11653\ : Span4Mux_h
    port map (
            O => \N__49123\,
            I => \N__49108\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__49120\,
            I => \N__49108\
        );

    \I__11651\ : Span4Mux_h
    port map (
            O => \N__49115\,
            I => \N__49108\
        );

    \I__11650\ : Odrv4
    port map (
            O => \N__49108\,
            I => \ALU.un2_addsub_cry_13_c_RNIR5I0EZ0\
        );

    \I__11649\ : CascadeMux
    port map (
            O => \N__49105\,
            I => \N__49102\
        );

    \I__11648\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49099\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__49099\,
            I => \ALU.r0_12_prm_2_14_s1_c_RNOZ0\
        );

    \I__11646\ : InMux
    port map (
            O => \N__49096\,
            I => \N__49093\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__49093\,
            I => \N__49090\
        );

    \I__11644\ : Span4Mux_v
    port map (
            O => \N__49090\,
            I => \N__49087\
        );

    \I__11643\ : Odrv4
    port map (
            O => \N__49087\,
            I => \ALU.r0_12_prm_1_14_s1_c_RNOZ0\
        );

    \I__11642\ : CascadeMux
    port map (
            O => \N__49084\,
            I => \N__49080\
        );

    \I__11641\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49077\
        );

    \I__11640\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49074\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__49077\,
            I => \N__49070\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__49074\,
            I => \N__49067\
        );

    \I__11637\ : InMux
    port map (
            O => \N__49073\,
            I => \N__49064\
        );

    \I__11636\ : Span4Mux_v
    port map (
            O => \N__49070\,
            I => \N__49061\
        );

    \I__11635\ : Span4Mux_v
    port map (
            O => \N__49067\,
            I => \N__49058\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__49064\,
            I => \N__49055\
        );

    \I__11633\ : Span4Mux_h
    port map (
            O => \N__49061\,
            I => \N__49049\
        );

    \I__11632\ : Span4Mux_h
    port map (
            O => \N__49058\,
            I => \N__49049\
        );

    \I__11631\ : Span4Mux_v
    port map (
            O => \N__49055\,
            I => \N__49046\
        );

    \I__11630\ : InMux
    port map (
            O => \N__49054\,
            I => \N__49043\
        );

    \I__11629\ : Odrv4
    port map (
            O => \N__49049\,
            I => \ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9\
        );

    \I__11628\ : Odrv4
    port map (
            O => \N__49046\,
            I => \ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__49043\,
            I => \ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9\
        );

    \I__11626\ : InMux
    port map (
            O => \N__49036\,
            I => \ALU.r0_12_s1_14\
        );

    \I__11625\ : InMux
    port map (
            O => \N__49033\,
            I => \N__49030\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__49030\,
            I => \N__49027\
        );

    \I__11623\ : Span4Mux_h
    port map (
            O => \N__49027\,
            I => \N__49024\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__49024\,
            I => \N__49021\
        );

    \I__11621\ : Odrv4
    port map (
            O => \N__49021\,
            I => \ALU.r0_12_s1_14_THRU_CO\
        );

    \I__11620\ : CascadeMux
    port map (
            O => \N__49018\,
            I => \N__49009\
        );

    \I__11619\ : InMux
    port map (
            O => \N__49017\,
            I => \N__49005\
        );

    \I__11618\ : InMux
    port map (
            O => \N__49016\,
            I => \N__48995\
        );

    \I__11617\ : InMux
    port map (
            O => \N__49015\,
            I => \N__48990\
        );

    \I__11616\ : InMux
    port map (
            O => \N__49014\,
            I => \N__48990\
        );

    \I__11615\ : InMux
    port map (
            O => \N__49013\,
            I => \N__48984\
        );

    \I__11614\ : InMux
    port map (
            O => \N__49012\,
            I => \N__48980\
        );

    \I__11613\ : InMux
    port map (
            O => \N__49009\,
            I => \N__48977\
        );

    \I__11612\ : InMux
    port map (
            O => \N__49008\,
            I => \N__48974\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48971\
        );

    \I__11610\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48968\
        );

    \I__11609\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48965\
        );

    \I__11608\ : InMux
    port map (
            O => \N__49002\,
            I => \N__48962\
        );

    \I__11607\ : InMux
    port map (
            O => \N__49001\,
            I => \N__48959\
        );

    \I__11606\ : InMux
    port map (
            O => \N__49000\,
            I => \N__48956\
        );

    \I__11605\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48950\
        );

    \I__11604\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48950\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__48995\,
            I => \N__48946\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__48990\,
            I => \N__48940\
        );

    \I__11601\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48937\
        );

    \I__11600\ : CascadeMux
    port map (
            O => \N__48988\,
            I => \N__48929\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__48987\,
            I => \N__48923\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__48984\,
            I => \N__48917\
        );

    \I__11597\ : InMux
    port map (
            O => \N__48983\,
            I => \N__48904\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__48980\,
            I => \N__48901\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__48977\,
            I => \N__48894\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__48974\,
            I => \N__48894\
        );

    \I__11593\ : Span4Mux_v
    port map (
            O => \N__48971\,
            I => \N__48894\
        );

    \I__11592\ : LocalMux
    port map (
            O => \N__48968\,
            I => \N__48891\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__48965\,
            I => \N__48888\
        );

    \I__11590\ : LocalMux
    port map (
            O => \N__48962\,
            I => \N__48885\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__48959\,
            I => \N__48880\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__48956\,
            I => \N__48880\
        );

    \I__11587\ : InMux
    port map (
            O => \N__48955\,
            I => \N__48877\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__48950\,
            I => \N__48874\
        );

    \I__11585\ : InMux
    port map (
            O => \N__48949\,
            I => \N__48871\
        );

    \I__11584\ : Span4Mux_v
    port map (
            O => \N__48946\,
            I => \N__48867\
        );

    \I__11583\ : InMux
    port map (
            O => \N__48945\,
            I => \N__48860\
        );

    \I__11582\ : InMux
    port map (
            O => \N__48944\,
            I => \N__48860\
        );

    \I__11581\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48860\
        );

    \I__11580\ : Span4Mux_s2_v
    port map (
            O => \N__48940\,
            I => \N__48855\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48855\
        );

    \I__11578\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48846\
        );

    \I__11577\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48846\
        );

    \I__11576\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48846\
        );

    \I__11575\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48846\
        );

    \I__11574\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48839\
        );

    \I__11573\ : InMux
    port map (
            O => \N__48929\,
            I => \N__48839\
        );

    \I__11572\ : InMux
    port map (
            O => \N__48928\,
            I => \N__48839\
        );

    \I__11571\ : InMux
    port map (
            O => \N__48927\,
            I => \N__48834\
        );

    \I__11570\ : InMux
    port map (
            O => \N__48926\,
            I => \N__48834\
        );

    \I__11569\ : InMux
    port map (
            O => \N__48923\,
            I => \N__48831\
        );

    \I__11568\ : InMux
    port map (
            O => \N__48922\,
            I => \N__48827\
        );

    \I__11567\ : InMux
    port map (
            O => \N__48921\,
            I => \N__48822\
        );

    \I__11566\ : InMux
    port map (
            O => \N__48920\,
            I => \N__48822\
        );

    \I__11565\ : Span4Mux_s3_h
    port map (
            O => \N__48917\,
            I => \N__48819\
        );

    \I__11564\ : InMux
    port map (
            O => \N__48916\,
            I => \N__48816\
        );

    \I__11563\ : InMux
    port map (
            O => \N__48915\,
            I => \N__48809\
        );

    \I__11562\ : InMux
    port map (
            O => \N__48914\,
            I => \N__48809\
        );

    \I__11561\ : InMux
    port map (
            O => \N__48913\,
            I => \N__48809\
        );

    \I__11560\ : InMux
    port map (
            O => \N__48912\,
            I => \N__48802\
        );

    \I__11559\ : InMux
    port map (
            O => \N__48911\,
            I => \N__48802\
        );

    \I__11558\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48802\
        );

    \I__11557\ : InMux
    port map (
            O => \N__48909\,
            I => \N__48799\
        );

    \I__11556\ : InMux
    port map (
            O => \N__48908\,
            I => \N__48794\
        );

    \I__11555\ : InMux
    port map (
            O => \N__48907\,
            I => \N__48794\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__48904\,
            I => \N__48785\
        );

    \I__11553\ : Span4Mux_h
    port map (
            O => \N__48901\,
            I => \N__48785\
        );

    \I__11552\ : Span4Mux_v
    port map (
            O => \N__48894\,
            I => \N__48785\
        );

    \I__11551\ : Span4Mux_s2_h
    port map (
            O => \N__48891\,
            I => \N__48782\
        );

    \I__11550\ : Span4Mux_s1_v
    port map (
            O => \N__48888\,
            I => \N__48779\
        );

    \I__11549\ : Span4Mux_s1_v
    port map (
            O => \N__48885\,
            I => \N__48770\
        );

    \I__11548\ : Span4Mux_h
    port map (
            O => \N__48880\,
            I => \N__48770\
        );

    \I__11547\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48770\
        );

    \I__11546\ : Span4Mux_v
    port map (
            O => \N__48874\,
            I => \N__48770\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__48871\,
            I => \N__48767\
        );

    \I__11544\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48764\
        );

    \I__11543\ : Span4Mux_h
    port map (
            O => \N__48867\,
            I => \N__48750\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__48860\,
            I => \N__48750\
        );

    \I__11541\ : Span4Mux_v
    port map (
            O => \N__48855\,
            I => \N__48750\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__48846\,
            I => \N__48750\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__48839\,
            I => \N__48747\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__48834\,
            I => \N__48742\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__48831\,
            I => \N__48742\
        );

    \I__11536\ : InMux
    port map (
            O => \N__48830\,
            I => \N__48739\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__48827\,
            I => \N__48736\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__48822\,
            I => \N__48727\
        );

    \I__11533\ : Span4Mux_v
    port map (
            O => \N__48819\,
            I => \N__48727\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__48816\,
            I => \N__48727\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__48809\,
            I => \N__48727\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__48802\,
            I => \N__48724\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__48799\,
            I => \N__48719\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__48794\,
            I => \N__48719\
        );

    \I__11527\ : InMux
    port map (
            O => \N__48793\,
            I => \N__48716\
        );

    \I__11526\ : InMux
    port map (
            O => \N__48792\,
            I => \N__48713\
        );

    \I__11525\ : Span4Mux_h
    port map (
            O => \N__48785\,
            I => \N__48708\
        );

    \I__11524\ : Span4Mux_h
    port map (
            O => \N__48782\,
            I => \N__48708\
        );

    \I__11523\ : Span4Mux_h
    port map (
            O => \N__48779\,
            I => \N__48699\
        );

    \I__11522\ : Span4Mux_h
    port map (
            O => \N__48770\,
            I => \N__48699\
        );

    \I__11521\ : Span4Mux_s1_v
    port map (
            O => \N__48767\,
            I => \N__48699\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__48764\,
            I => \N__48699\
        );

    \I__11519\ : InMux
    port map (
            O => \N__48763\,
            I => \N__48690\
        );

    \I__11518\ : InMux
    port map (
            O => \N__48762\,
            I => \N__48690\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48761\,
            I => \N__48690\
        );

    \I__11516\ : InMux
    port map (
            O => \N__48760\,
            I => \N__48690\
        );

    \I__11515\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48687\
        );

    \I__11514\ : Span4Mux_h
    port map (
            O => \N__48750\,
            I => \N__48674\
        );

    \I__11513\ : Span4Mux_s3_h
    port map (
            O => \N__48747\,
            I => \N__48674\
        );

    \I__11512\ : Span4Mux_s2_v
    port map (
            O => \N__48742\,
            I => \N__48674\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48674\
        );

    \I__11510\ : Span4Mux_s2_v
    port map (
            O => \N__48736\,
            I => \N__48674\
        );

    \I__11509\ : Span4Mux_v
    port map (
            O => \N__48727\,
            I => \N__48674\
        );

    \I__11508\ : Odrv4
    port map (
            O => \N__48724\,
            I => \ALU.aZ0Z_0\
        );

    \I__11507\ : Odrv12
    port map (
            O => \N__48719\,
            I => \ALU.aZ0Z_0\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__48716\,
            I => \ALU.aZ0Z_0\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__48713\,
            I => \ALU.aZ0Z_0\
        );

    \I__11504\ : Odrv4
    port map (
            O => \N__48708\,
            I => \ALU.aZ0Z_0\
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__48699\,
            I => \ALU.aZ0Z_0\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__48690\,
            I => \ALU.aZ0Z_0\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__48687\,
            I => \ALU.aZ0Z_0\
        );

    \I__11500\ : Odrv4
    port map (
            O => \N__48674\,
            I => \ALU.aZ0Z_0\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48649\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48654\,
            I => \N__48644\
        );

    \I__11497\ : InMux
    port map (
            O => \N__48653\,
            I => \N__48641\
        );

    \I__11496\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48635\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__48649\,
            I => \N__48632\
        );

    \I__11494\ : InMux
    port map (
            O => \N__48648\,
            I => \N__48629\
        );

    \I__11493\ : InMux
    port map (
            O => \N__48647\,
            I => \N__48626\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__48644\,
            I => \N__48621\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__48641\,
            I => \N__48621\
        );

    \I__11490\ : InMux
    port map (
            O => \N__48640\,
            I => \N__48618\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48605\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48602\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__48635\,
            I => \N__48597\
        );

    \I__11486\ : Span4Mux_v
    port map (
            O => \N__48632\,
            I => \N__48597\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__48629\,
            I => \N__48594\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__48626\,
            I => \N__48587\
        );

    \I__11483\ : Span4Mux_v
    port map (
            O => \N__48621\,
            I => \N__48587\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__48618\,
            I => \N__48587\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48617\,
            I => \N__48582\
        );

    \I__11480\ : InMux
    port map (
            O => \N__48616\,
            I => \N__48582\
        );

    \I__11479\ : InMux
    port map (
            O => \N__48615\,
            I => \N__48577\
        );

    \I__11478\ : InMux
    port map (
            O => \N__48614\,
            I => \N__48577\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48613\,
            I => \N__48572\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48612\,
            I => \N__48564\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48611\,
            I => \N__48561\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48610\,
            I => \N__48554\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48609\,
            I => \N__48554\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48608\,
            I => \N__48554\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__48605\,
            I => \N__48550\
        );

    \I__11470\ : LocalMux
    port map (
            O => \N__48602\,
            I => \N__48545\
        );

    \I__11469\ : Span4Mux_v
    port map (
            O => \N__48597\,
            I => \N__48545\
        );

    \I__11468\ : Span4Mux_h
    port map (
            O => \N__48594\,
            I => \N__48536\
        );

    \I__11467\ : Span4Mux_v
    port map (
            O => \N__48587\,
            I => \N__48536\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__48582\,
            I => \N__48536\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__48577\,
            I => \N__48536\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48576\,
            I => \N__48531\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48575\,
            I => \N__48531\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__48572\,
            I => \N__48528\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48571\,
            I => \N__48521\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48570\,
            I => \N__48521\
        );

    \I__11459\ : InMux
    port map (
            O => \N__48569\,
            I => \N__48521\
        );

    \I__11458\ : InMux
    port map (
            O => \N__48568\,
            I => \N__48516\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48516\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__48564\,
            I => \N__48506\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__48561\,
            I => \N__48500\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__48554\,
            I => \N__48500\
        );

    \I__11453\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48497\
        );

    \I__11452\ : Span4Mux_s3_v
    port map (
            O => \N__48550\,
            I => \N__48490\
        );

    \I__11451\ : Span4Mux_v
    port map (
            O => \N__48545\,
            I => \N__48490\
        );

    \I__11450\ : Span4Mux_h
    port map (
            O => \N__48536\,
            I => \N__48490\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__48531\,
            I => \N__48487\
        );

    \I__11448\ : Span4Mux_h
    port map (
            O => \N__48528\,
            I => \N__48484\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__48521\,
            I => \N__48479\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__48516\,
            I => \N__48479\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48515\,
            I => \N__48474\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48514\,
            I => \N__48474\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48513\,
            I => \N__48469\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48512\,
            I => \N__48464\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48511\,
            I => \N__48464\
        );

    \I__11440\ : InMux
    port map (
            O => \N__48510\,
            I => \N__48461\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48509\,
            I => \N__48458\
        );

    \I__11438\ : Span4Mux_s3_v
    port map (
            O => \N__48506\,
            I => \N__48455\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48452\
        );

    \I__11436\ : Span4Mux_v
    port map (
            O => \N__48500\,
            I => \N__48443\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48443\
        );

    \I__11434\ : Span4Mux_h
    port map (
            O => \N__48490\,
            I => \N__48443\
        );

    \I__11433\ : Span4Mux_s3_v
    port map (
            O => \N__48487\,
            I => \N__48443\
        );

    \I__11432\ : Span4Mux_v
    port map (
            O => \N__48484\,
            I => \N__48436\
        );

    \I__11431\ : Span4Mux_h
    port map (
            O => \N__48479\,
            I => \N__48436\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__48474\,
            I => \N__48436\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48473\,
            I => \N__48431\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48472\,
            I => \N__48431\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48426\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48426\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__48461\,
            I => \ALU.a_1\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__48458\,
            I => \ALU.a_1\
        );

    \I__11423\ : Odrv4
    port map (
            O => \N__48455\,
            I => \ALU.a_1\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__48452\,
            I => \ALU.a_1\
        );

    \I__11421\ : Odrv4
    port map (
            O => \N__48443\,
            I => \ALU.a_1\
        );

    \I__11420\ : Odrv4
    port map (
            O => \N__48436\,
            I => \ALU.a_1\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48431\,
            I => \ALU.a_1\
        );

    \I__11418\ : Odrv4
    port map (
            O => \N__48426\,
            I => \ALU.a_1\
        );

    \I__11417\ : CascadeMux
    port map (
            O => \N__48409\,
            I => \N__48396\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48408\,
            I => \N__48392\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48407\,
            I => \N__48387\
        );

    \I__11414\ : InMux
    port map (
            O => \N__48406\,
            I => \N__48384\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48405\,
            I => \N__48381\
        );

    \I__11412\ : InMux
    port map (
            O => \N__48404\,
            I => \N__48378\
        );

    \I__11411\ : InMux
    port map (
            O => \N__48403\,
            I => \N__48373\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48373\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48401\,
            I => \N__48370\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48400\,
            I => \N__48367\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48399\,
            I => \N__48358\
        );

    \I__11406\ : InMux
    port map (
            O => \N__48396\,
            I => \N__48355\
        );

    \I__11405\ : InMux
    port map (
            O => \N__48395\,
            I => \N__48352\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48392\,
            I => \N__48348\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48391\,
            I => \N__48343\
        );

    \I__11402\ : InMux
    port map (
            O => \N__48390\,
            I => \N__48343\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__48387\,
            I => \N__48339\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__48384\,
            I => \N__48336\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__48381\,
            I => \N__48330\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48330\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48327\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__48370\,
            I => \N__48324\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48320\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48366\,
            I => \N__48315\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48365\,
            I => \N__48315\
        );

    \I__11392\ : InMux
    port map (
            O => \N__48364\,
            I => \N__48308\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48308\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48362\,
            I => \N__48308\
        );

    \I__11389\ : InMux
    port map (
            O => \N__48361\,
            I => \N__48304\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__48358\,
            I => \N__48301\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__48355\,
            I => \N__48296\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__48352\,
            I => \N__48296\
        );

    \I__11385\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48293\
        );

    \I__11384\ : Span4Mux_v
    port map (
            O => \N__48348\,
            I => \N__48285\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__48343\,
            I => \N__48282\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48279\
        );

    \I__11381\ : Span4Mux_s3_v
    port map (
            O => \N__48339\,
            I => \N__48274\
        );

    \I__11380\ : Span4Mux_s3_v
    port map (
            O => \N__48336\,
            I => \N__48274\
        );

    \I__11379\ : InMux
    port map (
            O => \N__48335\,
            I => \N__48271\
        );

    \I__11378\ : Span4Mux_s3_v
    port map (
            O => \N__48330\,
            I => \N__48264\
        );

    \I__11377\ : Span4Mux_s3_v
    port map (
            O => \N__48327\,
            I => \N__48264\
        );

    \I__11376\ : Span4Mux_v
    port map (
            O => \N__48324\,
            I => \N__48264\
        );

    \I__11375\ : InMux
    port map (
            O => \N__48323\,
            I => \N__48261\
        );

    \I__11374\ : Span4Mux_v
    port map (
            O => \N__48320\,
            I => \N__48258\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48315\,
            I => \N__48253\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__48308\,
            I => \N__48253\
        );

    \I__11371\ : InMux
    port map (
            O => \N__48307\,
            I => \N__48250\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__48304\,
            I => \N__48247\
        );

    \I__11369\ : Span4Mux_s3_v
    port map (
            O => \N__48301\,
            I => \N__48242\
        );

    \I__11368\ : Span4Mux_v
    port map (
            O => \N__48296\,
            I => \N__48242\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__48293\,
            I => \N__48239\
        );

    \I__11366\ : CascadeMux
    port map (
            O => \N__48292\,
            I => \N__48236\
        );

    \I__11365\ : InMux
    port map (
            O => \N__48291\,
            I => \N__48230\
        );

    \I__11364\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48230\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48289\,
            I => \N__48225\
        );

    \I__11362\ : InMux
    port map (
            O => \N__48288\,
            I => \N__48225\
        );

    \I__11361\ : Span4Mux_h
    port map (
            O => \N__48285\,
            I => \N__48222\
        );

    \I__11360\ : Span4Mux_v
    port map (
            O => \N__48282\,
            I => \N__48217\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__48279\,
            I => \N__48217\
        );

    \I__11358\ : Sp12to4
    port map (
            O => \N__48274\,
            I => \N__48206\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__48271\,
            I => \N__48206\
        );

    \I__11356\ : Sp12to4
    port map (
            O => \N__48264\,
            I => \N__48206\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__48261\,
            I => \N__48206\
        );

    \I__11354\ : Sp12to4
    port map (
            O => \N__48258\,
            I => \N__48206\
        );

    \I__11353\ : Span4Mux_v
    port map (
            O => \N__48253\,
            I => \N__48195\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__48250\,
            I => \N__48195\
        );

    \I__11351\ : Span4Mux_s3_v
    port map (
            O => \N__48247\,
            I => \N__48195\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__48242\,
            I => \N__48195\
        );

    \I__11349\ : Span4Mux_s3_v
    port map (
            O => \N__48239\,
            I => \N__48195\
        );

    \I__11348\ : InMux
    port map (
            O => \N__48236\,
            I => \N__48190\
        );

    \I__11347\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48190\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__48230\,
            I => \N__48185\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__48225\,
            I => \N__48185\
        );

    \I__11344\ : Span4Mux_v
    port map (
            O => \N__48222\,
            I => \N__48180\
        );

    \I__11343\ : Span4Mux_h
    port map (
            O => \N__48217\,
            I => \N__48180\
        );

    \I__11342\ : Odrv12
    port map (
            O => \N__48206\,
            I => \ALU.a_2\
        );

    \I__11341\ : Odrv4
    port map (
            O => \N__48195\,
            I => \ALU.a_2\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__48190\,
            I => \ALU.a_2\
        );

    \I__11339\ : Odrv4
    port map (
            O => \N__48185\,
            I => \ALU.a_2\
        );

    \I__11338\ : Odrv4
    port map (
            O => \N__48180\,
            I => \ALU.a_2\
        );

    \I__11337\ : CascadeMux
    port map (
            O => \N__48169\,
            I => \ALU.rshift_3_ns_1_0_cascade_\
        );

    \I__11336\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48163\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__48163\,
            I => \N__48160\
        );

    \I__11334\ : Span4Mux_s3_v
    port map (
            O => \N__48160\,
            I => \N__48157\
        );

    \I__11333\ : Span4Mux_h
    port map (
            O => \N__48157\,
            I => \N__48154\
        );

    \I__11332\ : Odrv4
    port map (
            O => \N__48154\,
            I => \ALU.r4_RNII2A0LZ0Z_2\
        );

    \I__11331\ : InMux
    port map (
            O => \N__48151\,
            I => \N__48147\
        );

    \I__11330\ : CascadeMux
    port map (
            O => \N__48150\,
            I => \N__48144\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__48147\,
            I => \N__48141\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48144\,
            I => \N__48138\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__48141\,
            I => \N__48131\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__48138\,
            I => \N__48131\
        );

    \I__11325\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48128\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48136\,
            I => \N__48125\
        );

    \I__11323\ : Odrv4
    port map (
            O => \N__48131\,
            I => \ALU.lshift_5\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__48128\,
            I => \ALU.lshift_5\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__48125\,
            I => \ALU.lshift_5\
        );

    \I__11320\ : CascadeMux
    port map (
            O => \N__48118\,
            I => \N__48115\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48112\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__48112\,
            I => \N__48109\
        );

    \I__11317\ : Span4Mux_h
    port map (
            O => \N__48109\,
            I => \N__48106\
        );

    \I__11316\ : Span4Mux_v
    port map (
            O => \N__48106\,
            I => \N__48103\
        );

    \I__11315\ : Odrv4
    port map (
            O => \N__48103\,
            I => \ALU.r0_12_prm_8_5_s0_c_RNOZ0\
        );

    \I__11314\ : CascadeMux
    port map (
            O => \N__48100\,
            I => \N__48097\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48097\,
            I => \N__48094\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__48094\,
            I => \N__48091\
        );

    \I__11311\ : Span4Mux_v
    port map (
            O => \N__48091\,
            I => \N__48088\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__48088\,
            I => \N__48085\
        );

    \I__11309\ : Span4Mux_h
    port map (
            O => \N__48085\,
            I => \N__48082\
        );

    \I__11308\ : Odrv4
    port map (
            O => \N__48082\,
            I => \ALU.r4_RNI0C236Z0Z_9\
        );

    \I__11307\ : InMux
    port map (
            O => \N__48079\,
            I => \N__48073\
        );

    \I__11306\ : InMux
    port map (
            O => \N__48078\,
            I => \N__48070\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48077\,
            I => \N__48065\
        );

    \I__11304\ : InMux
    port map (
            O => \N__48076\,
            I => \N__48065\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__48073\,
            I => \N__48062\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__48070\,
            I => \N__48058\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__48065\,
            I => \N__48055\
        );

    \I__11300\ : Span4Mux_h
    port map (
            O => \N__48062\,
            I => \N__48052\
        );

    \I__11299\ : CascadeMux
    port map (
            O => \N__48061\,
            I => \N__48049\
        );

    \I__11298\ : Span4Mux_v
    port map (
            O => \N__48058\,
            I => \N__48046\
        );

    \I__11297\ : Span4Mux_v
    port map (
            O => \N__48055\,
            I => \N__48043\
        );

    \I__11296\ : Span4Mux_h
    port map (
            O => \N__48052\,
            I => \N__48040\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48037\
        );

    \I__11294\ : Span4Mux_h
    port map (
            O => \N__48046\,
            I => \N__48034\
        );

    \I__11293\ : Span4Mux_h
    port map (
            O => \N__48043\,
            I => \N__48031\
        );

    \I__11292\ : Span4Mux_h
    port map (
            O => \N__48040\,
            I => \N__48026\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__48037\,
            I => \N__48026\
        );

    \I__11290\ : Span4Mux_h
    port map (
            O => \N__48034\,
            I => \N__48021\
        );

    \I__11289\ : Span4Mux_h
    port map (
            O => \N__48031\,
            I => \N__48021\
        );

    \I__11288\ : Span4Mux_v
    port map (
            O => \N__48026\,
            I => \N__48018\
        );

    \I__11287\ : Span4Mux_v
    port map (
            O => \N__48021\,
            I => \N__48015\
        );

    \I__11286\ : Span4Mux_s2_h
    port map (
            O => \N__48018\,
            I => \N__48012\
        );

    \I__11285\ : Span4Mux_h
    port map (
            O => \N__48015\,
            I => \N__48009\
        );

    \I__11284\ : Odrv4
    port map (
            O => \N__48012\,
            I => \ALU.a7_b_7\
        );

    \I__11283\ : Odrv4
    port map (
            O => \N__48009\,
            I => \ALU.a7_b_7\
        );

    \I__11282\ : CascadeMux
    port map (
            O => \N__48004\,
            I => \N__48001\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48001\,
            I => \N__47998\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__47998\,
            I => \N__47995\
        );

    \I__11279\ : Span4Mux_h
    port map (
            O => \N__47995\,
            I => \N__47992\
        );

    \I__11278\ : Span4Mux_v
    port map (
            O => \N__47992\,
            I => \N__47989\
        );

    \I__11277\ : Odrv4
    port map (
            O => \N__47989\,
            I => \ALU.r0_12_prm_7_7_s0_c_RNOZ0\
        );

    \I__11276\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47983\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__47983\,
            I => \ALU.r0_12_prm_8_14_s1_c_RNOZ0\
        );

    \I__11274\ : InMux
    port map (
            O => \N__47980\,
            I => \N__47977\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__47977\,
            I => \N__47973\
        );

    \I__11272\ : CascadeMux
    port map (
            O => \N__47976\,
            I => \N__47970\
        );

    \I__11271\ : Span4Mux_h
    port map (
            O => \N__47973\,
            I => \N__47966\
        );

    \I__11270\ : InMux
    port map (
            O => \N__47970\,
            I => \N__47963\
        );

    \I__11269\ : InMux
    port map (
            O => \N__47969\,
            I => \N__47960\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__47966\,
            I => \N__47956\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__47963\,
            I => \N__47953\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__47960\,
            I => \N__47950\
        );

    \I__11265\ : InMux
    port map (
            O => \N__47959\,
            I => \N__47947\
        );

    \I__11264\ : Odrv4
    port map (
            O => \N__47956\,
            I => \ALU.lshift_14\
        );

    \I__11263\ : Odrv4
    port map (
            O => \N__47953\,
            I => \ALU.lshift_14\
        );

    \I__11262\ : Odrv4
    port map (
            O => \N__47950\,
            I => \ALU.lshift_14\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__47947\,
            I => \ALU.lshift_14\
        );

    \I__11260\ : InMux
    port map (
            O => \N__47938\,
            I => \N__47935\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__47935\,
            I => \N__47932\
        );

    \I__11258\ : Odrv4
    port map (
            O => \N__47932\,
            I => \ALU.r0_12_prm_7_14_s1_c_RNOZ0\
        );

    \I__11257\ : CascadeMux
    port map (
            O => \N__47929\,
            I => \N__47925\
        );

    \I__11256\ : InMux
    port map (
            O => \N__47928\,
            I => \N__47922\
        );

    \I__11255\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47919\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__47922\,
            I => \N__47916\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__47919\,
            I => \N__47913\
        );

    \I__11252\ : Odrv12
    port map (
            O => \N__47916\,
            I => \ALU.r2_RNINPPC9_0Z0Z_14\
        );

    \I__11251\ : Odrv4
    port map (
            O => \N__47913\,
            I => \ALU.r2_RNINPPC9_0Z0Z_14\
        );

    \I__11250\ : InMux
    port map (
            O => \N__47908\,
            I => \N__47905\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__47905\,
            I => \N__47902\
        );

    \I__11248\ : Span4Mux_h
    port map (
            O => \N__47902\,
            I => \N__47899\
        );

    \I__11247\ : Odrv4
    port map (
            O => \N__47899\,
            I => \ALU.r0_12_prm_6_14_s1_c_RNOZ0\
        );

    \I__11246\ : CascadeMux
    port map (
            O => \N__47896\,
            I => \N__47892\
        );

    \I__11245\ : InMux
    port map (
            O => \N__47895\,
            I => \N__47889\
        );

    \I__11244\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47886\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__47889\,
            I => \N__47883\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__47886\,
            I => \N__47880\
        );

    \I__11241\ : Span4Mux_h
    port map (
            O => \N__47883\,
            I => \N__47875\
        );

    \I__11240\ : Span4Mux_h
    port map (
            O => \N__47880\,
            I => \N__47875\
        );

    \I__11239\ : Odrv4
    port map (
            O => \N__47875\,
            I => \ALU.un14_log_0_i_14\
        );

    \I__11238\ : InMux
    port map (
            O => \N__47872\,
            I => \N__47869\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__47869\,
            I => \ALU.r0_12_prm_5_14_s1_c_RNOZ0\
        );

    \I__11236\ : CascadeMux
    port map (
            O => \N__47866\,
            I => \N__47863\
        );

    \I__11235\ : InMux
    port map (
            O => \N__47863\,
            I => \N__47860\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__47860\,
            I => \N__47856\
        );

    \I__11233\ : CascadeMux
    port map (
            O => \N__47859\,
            I => \N__47853\
        );

    \I__11232\ : Span4Mux_h
    port map (
            O => \N__47856\,
            I => \N__47850\
        );

    \I__11231\ : InMux
    port map (
            O => \N__47853\,
            I => \N__47847\
        );

    \I__11230\ : Odrv4
    port map (
            O => \N__47850\,
            I => \ALU.r2_RNINPPC9_1Z0Z_14\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__47847\,
            I => \ALU.r2_RNINPPC9_1Z0Z_14\
        );

    \I__11228\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47839\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__47839\,
            I => \N__47836\
        );

    \I__11226\ : Odrv4
    port map (
            O => \N__47836\,
            I => \ALU.r0_12_prm_4_14_s1_c_RNOZ0\
        );

    \I__11225\ : CascadeMux
    port map (
            O => \N__47833\,
            I => \N__47830\
        );

    \I__11224\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47827\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__47827\,
            I => \N__47824\
        );

    \I__11222\ : Span4Mux_h
    port map (
            O => \N__47824\,
            I => \N__47820\
        );

    \I__11221\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47817\
        );

    \I__11220\ : Span4Mux_h
    port map (
            O => \N__47820\,
            I => \N__47814\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__47817\,
            I => \ALU.a_i_14\
        );

    \I__11218\ : Odrv4
    port map (
            O => \N__47814\,
            I => \ALU.a_i_14\
        );

    \I__11217\ : CEMux
    port map (
            O => \N__47809\,
            I => \N__47806\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__47806\,
            I => \N__47803\
        );

    \I__11215\ : Span4Mux_v
    port map (
            O => \N__47803\,
            I => \N__47799\
        );

    \I__11214\ : CEMux
    port map (
            O => \N__47802\,
            I => \N__47796\
        );

    \I__11213\ : Span4Mux_h
    port map (
            O => \N__47799\,
            I => \N__47791\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__47796\,
            I => \N__47791\
        );

    \I__11211\ : Span4Mux_v
    port map (
            O => \N__47791\,
            I => \N__47788\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__47788\,
            I => \N__47784\
        );

    \I__11209\ : CEMux
    port map (
            O => \N__47787\,
            I => \N__47781\
        );

    \I__11208\ : Span4Mux_h
    port map (
            O => \N__47784\,
            I => \N__47778\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__47781\,
            I => \N__47775\
        );

    \I__11206\ : Span4Mux_h
    port map (
            O => \N__47778\,
            I => \N__47772\
        );

    \I__11205\ : Sp12to4
    port map (
            O => \N__47775\,
            I => \N__47769\
        );

    \I__11204\ : Odrv4
    port map (
            O => \N__47772\,
            I => \ALU.un1_yindexZ0Z_4\
        );

    \I__11203\ : Odrv12
    port map (
            O => \N__47769\,
            I => \ALU.un1_yindexZ0Z_4\
        );

    \I__11202\ : CEMux
    port map (
            O => \N__47764\,
            I => \N__47759\
        );

    \I__11201\ : CEMux
    port map (
            O => \N__47763\,
            I => \N__47756\
        );

    \I__11200\ : CEMux
    port map (
            O => \N__47762\,
            I => \N__47752\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47749\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__47756\,
            I => \N__47746\
        );

    \I__11197\ : CEMux
    port map (
            O => \N__47755\,
            I => \N__47743\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__47752\,
            I => \N__47736\
        );

    \I__11195\ : Span4Mux_v
    port map (
            O => \N__47749\,
            I => \N__47736\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__47746\,
            I => \N__47736\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__47743\,
            I => \N__47733\
        );

    \I__11192\ : Span4Mux_h
    port map (
            O => \N__47736\,
            I => \N__47730\
        );

    \I__11191\ : Sp12to4
    port map (
            O => \N__47733\,
            I => \N__47727\
        );

    \I__11190\ : Sp12to4
    port map (
            O => \N__47730\,
            I => \N__47724\
        );

    \I__11189\ : Span12Mux_s5_h
    port map (
            O => \N__47727\,
            I => \N__47719\
        );

    \I__11188\ : Span12Mux_v
    port map (
            O => \N__47724\,
            I => \N__47719\
        );

    \I__11187\ : Odrv12
    port map (
            O => \N__47719\,
            I => \ALU.un1_yindexZ0Z_5\
        );

    \I__11186\ : CEMux
    port map (
            O => \N__47716\,
            I => \N__47713\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__47713\,
            I => \N__47709\
        );

    \I__11184\ : CEMux
    port map (
            O => \N__47712\,
            I => \N__47703\
        );

    \I__11183\ : IoSpan4Mux
    port map (
            O => \N__47709\,
            I => \N__47700\
        );

    \I__11182\ : CEMux
    port map (
            O => \N__47708\,
            I => \N__47697\
        );

    \I__11181\ : CEMux
    port map (
            O => \N__47707\,
            I => \N__47694\
        );

    \I__11180\ : CEMux
    port map (
            O => \N__47706\,
            I => \N__47691\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__47703\,
            I => \N__47687\
        );

    \I__11178\ : Span4Mux_s1_h
    port map (
            O => \N__47700\,
            I => \N__47681\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47681\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__47694\,
            I => \N__47678\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__47691\,
            I => \N__47675\
        );

    \I__11174\ : CEMux
    port map (
            O => \N__47690\,
            I => \N__47672\
        );

    \I__11173\ : Span4Mux_s2_h
    port map (
            O => \N__47687\,
            I => \N__47668\
        );

    \I__11172\ : CEMux
    port map (
            O => \N__47686\,
            I => \N__47665\
        );

    \I__11171\ : Span4Mux_h
    port map (
            O => \N__47681\,
            I => \N__47661\
        );

    \I__11170\ : Span4Mux_s3_h
    port map (
            O => \N__47678\,
            I => \N__47656\
        );

    \I__11169\ : Span4Mux_s3_h
    port map (
            O => \N__47675\,
            I => \N__47656\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__47672\,
            I => \N__47653\
        );

    \I__11167\ : CEMux
    port map (
            O => \N__47671\,
            I => \N__47650\
        );

    \I__11166\ : Span4Mux_v
    port map (
            O => \N__47668\,
            I => \N__47645\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__47665\,
            I => \N__47645\
        );

    \I__11164\ : CEMux
    port map (
            O => \N__47664\,
            I => \N__47642\
        );

    \I__11163\ : Span4Mux_h
    port map (
            O => \N__47661\,
            I => \N__47639\
        );

    \I__11162\ : Span4Mux_h
    port map (
            O => \N__47656\,
            I => \N__47634\
        );

    \I__11161\ : Span4Mux_h
    port map (
            O => \N__47653\,
            I => \N__47634\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__47650\,
            I => \N__47631\
        );

    \I__11159\ : Span4Mux_h
    port map (
            O => \N__47645\,
            I => \N__47628\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__47642\,
            I => \N__47625\
        );

    \I__11157\ : Span4Mux_v
    port map (
            O => \N__47639\,
            I => \N__47622\
        );

    \I__11156\ : Span4Mux_v
    port map (
            O => \N__47634\,
            I => \N__47619\
        );

    \I__11155\ : Span4Mux_h
    port map (
            O => \N__47631\,
            I => \N__47616\
        );

    \I__11154\ : Span4Mux_v
    port map (
            O => \N__47628\,
            I => \N__47611\
        );

    \I__11153\ : Span4Mux_v
    port map (
            O => \N__47625\,
            I => \N__47611\
        );

    \I__11152\ : Sp12to4
    port map (
            O => \N__47622\,
            I => \N__47608\
        );

    \I__11151\ : Span4Mux_h
    port map (
            O => \N__47619\,
            I => \N__47605\
        );

    \I__11150\ : Span4Mux_h
    port map (
            O => \N__47616\,
            I => \N__47602\
        );

    \I__11149\ : Span4Mux_h
    port map (
            O => \N__47611\,
            I => \N__47599\
        );

    \I__11148\ : Span12Mux_h
    port map (
            O => \N__47608\,
            I => \N__47596\
        );

    \I__11147\ : Span4Mux_h
    port map (
            O => \N__47605\,
            I => \N__47593\
        );

    \I__11146\ : Span4Mux_v
    port map (
            O => \N__47602\,
            I => \N__47588\
        );

    \I__11145\ : Span4Mux_h
    port map (
            O => \N__47599\,
            I => \N__47588\
        );

    \I__11144\ : Odrv12
    port map (
            O => \N__47596\,
            I => \ALU.un1_yindexZ0Z_6\
        );

    \I__11143\ : Odrv4
    port map (
            O => \N__47593\,
            I => \ALU.un1_yindexZ0Z_6\
        );

    \I__11142\ : Odrv4
    port map (
            O => \N__47588\,
            I => \ALU.un1_yindexZ0Z_6\
        );

    \I__11141\ : CEMux
    port map (
            O => \N__47581\,
            I => \N__47578\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__47578\,
            I => \N__47573\
        );

    \I__11139\ : CEMux
    port map (
            O => \N__47577\,
            I => \N__47570\
        );

    \I__11138\ : CEMux
    port map (
            O => \N__47576\,
            I => \N__47566\
        );

    \I__11137\ : Span4Mux_h
    port map (
            O => \N__47573\,
            I => \N__47561\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__47570\,
            I => \N__47561\
        );

    \I__11135\ : CEMux
    port map (
            O => \N__47569\,
            I => \N__47556\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__47566\,
            I => \N__47553\
        );

    \I__11133\ : Span4Mux_v
    port map (
            O => \N__47561\,
            I => \N__47550\
        );

    \I__11132\ : CEMux
    port map (
            O => \N__47560\,
            I => \N__47547\
        );

    \I__11131\ : CEMux
    port map (
            O => \N__47559\,
            I => \N__47544\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47556\,
            I => \N__47540\
        );

    \I__11129\ : Span4Mux_h
    port map (
            O => \N__47553\,
            I => \N__47537\
        );

    \I__11128\ : Span4Mux_h
    port map (
            O => \N__47550\,
            I => \N__47534\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__47547\,
            I => \N__47531\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__47544\,
            I => \N__47528\
        );

    \I__11125\ : CEMux
    port map (
            O => \N__47543\,
            I => \N__47525\
        );

    \I__11124\ : Span4Mux_h
    port map (
            O => \N__47540\,
            I => \N__47522\
        );

    \I__11123\ : Span4Mux_h
    port map (
            O => \N__47537\,
            I => \N__47519\
        );

    \I__11122\ : Sp12to4
    port map (
            O => \N__47534\,
            I => \N__47516\
        );

    \I__11121\ : Span4Mux_h
    port map (
            O => \N__47531\,
            I => \N__47513\
        );

    \I__11120\ : Span4Mux_h
    port map (
            O => \N__47528\,
            I => \N__47508\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__47525\,
            I => \N__47508\
        );

    \I__11118\ : Span4Mux_h
    port map (
            O => \N__47522\,
            I => \N__47505\
        );

    \I__11117\ : Span4Mux_v
    port map (
            O => \N__47519\,
            I => \N__47502\
        );

    \I__11116\ : Span12Mux_h
    port map (
            O => \N__47516\,
            I => \N__47499\
        );

    \I__11115\ : Span4Mux_h
    port map (
            O => \N__47513\,
            I => \N__47496\
        );

    \I__11114\ : Span4Mux_v
    port map (
            O => \N__47508\,
            I => \N__47493\
        );

    \I__11113\ : Odrv4
    port map (
            O => \N__47505\,
            I => \ALU.un1_yindexZ0Z_7\
        );

    \I__11112\ : Odrv4
    port map (
            O => \N__47502\,
            I => \ALU.un1_yindexZ0Z_7\
        );

    \I__11111\ : Odrv12
    port map (
            O => \N__47499\,
            I => \ALU.un1_yindexZ0Z_7\
        );

    \I__11110\ : Odrv4
    port map (
            O => \N__47496\,
            I => \ALU.un1_yindexZ0Z_7\
        );

    \I__11109\ : Odrv4
    port map (
            O => \N__47493\,
            I => \ALU.un1_yindexZ0Z_7\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47479\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47479\,
            I => \N__47467\
        );

    \I__11106\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47464\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47461\
        );

    \I__11104\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47458\
        );

    \I__11103\ : CascadeMux
    port map (
            O => \N__47475\,
            I => \N__47452\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47474\,
            I => \N__47449\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47473\,
            I => \N__47446\
        );

    \I__11100\ : InMux
    port map (
            O => \N__47472\,
            I => \N__47443\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47440\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47437\
        );

    \I__11097\ : Span4Mux_h
    port map (
            O => \N__47467\,
            I => \N__47426\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__47464\,
            I => \N__47426\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__47461\,
            I => \N__47426\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47458\,
            I => \N__47426\
        );

    \I__11093\ : CascadeMux
    port map (
            O => \N__47457\,
            I => \N__47420\
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__47456\,
            I => \N__47417\
        );

    \I__11091\ : CascadeMux
    port map (
            O => \N__47455\,
            I => \N__47414\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47410\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__47449\,
            I => \N__47407\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__47446\,
            I => \N__47398\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__47443\,
            I => \N__47398\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__47440\,
            I => \N__47398\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47437\,
            I => \N__47398\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47436\,
            I => \N__47395\
        );

    \I__11083\ : CascadeMux
    port map (
            O => \N__47435\,
            I => \N__47391\
        );

    \I__11082\ : Span4Mux_h
    port map (
            O => \N__47426\,
            I => \N__47388\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47425\,
            I => \N__47385\
        );

    \I__11080\ : InMux
    port map (
            O => \N__47424\,
            I => \N__47382\
        );

    \I__11079\ : InMux
    port map (
            O => \N__47423\,
            I => \N__47377\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47420\,
            I => \N__47377\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47417\,
            I => \N__47374\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47414\,
            I => \N__47369\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47369\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47410\,
            I => \N__47366\
        );

    \I__11073\ : Span4Mux_v
    port map (
            O => \N__47407\,
            I => \N__47361\
        );

    \I__11072\ : Span4Mux_v
    port map (
            O => \N__47398\,
            I => \N__47361\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__47395\,
            I => \N__47358\
        );

    \I__11070\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47353\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47391\,
            I => \N__47353\
        );

    \I__11068\ : Span4Mux_h
    port map (
            O => \N__47388\,
            I => \N__47349\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__47385\,
            I => \N__47346\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47382\,
            I => \N__47343\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__47377\,
            I => \N__47335\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__47374\,
            I => \N__47335\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__47369\,
            I => \N__47335\
        );

    \I__11062\ : Span4Mux_v
    port map (
            O => \N__47366\,
            I => \N__47330\
        );

    \I__11061\ : Span4Mux_h
    port map (
            O => \N__47361\,
            I => \N__47330\
        );

    \I__11060\ : Span4Mux_v
    port map (
            O => \N__47358\,
            I => \N__47325\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__47353\,
            I => \N__47325\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47352\,
            I => \N__47322\
        );

    \I__11057\ : Span4Mux_v
    port map (
            O => \N__47349\,
            I => \N__47317\
        );

    \I__11056\ : Span4Mux_v
    port map (
            O => \N__47346\,
            I => \N__47317\
        );

    \I__11055\ : Span4Mux_s3_v
    port map (
            O => \N__47343\,
            I => \N__47314\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47342\,
            I => \N__47311\
        );

    \I__11053\ : Span4Mux_v
    port map (
            O => \N__47335\,
            I => \N__47308\
        );

    \I__11052\ : Sp12to4
    port map (
            O => \N__47330\,
            I => \N__47305\
        );

    \I__11051\ : Span4Mux_h
    port map (
            O => \N__47325\,
            I => \N__47302\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47322\,
            I => \ALU.b_9\
        );

    \I__11049\ : Odrv4
    port map (
            O => \N__47317\,
            I => \ALU.b_9\
        );

    \I__11048\ : Odrv4
    port map (
            O => \N__47314\,
            I => \ALU.b_9\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__47311\,
            I => \ALU.b_9\
        );

    \I__11046\ : Odrv4
    port map (
            O => \N__47308\,
            I => \ALU.b_9\
        );

    \I__11045\ : Odrv12
    port map (
            O => \N__47305\,
            I => \ALU.b_9\
        );

    \I__11044\ : Odrv4
    port map (
            O => \N__47302\,
            I => \ALU.b_9\
        );

    \I__11043\ : CascadeMux
    port map (
            O => \N__47287\,
            I => \N__47284\
        );

    \I__11042\ : InMux
    port map (
            O => \N__47284\,
            I => \N__47281\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__47281\,
            I => \N__47278\
        );

    \I__11040\ : Span4Mux_h
    port map (
            O => \N__47278\,
            I => \N__47275\
        );

    \I__11039\ : Span4Mux_h
    port map (
            O => \N__47275\,
            I => \N__47272\
        );

    \I__11038\ : Odrv4
    port map (
            O => \N__47272\,
            I => \ALU.r4_RNISU5D9_2Z0Z_9\
        );

    \I__11037\ : CascadeMux
    port map (
            O => \N__47269\,
            I => \N__47262\
        );

    \I__11036\ : CascadeMux
    port map (
            O => \N__47268\,
            I => \N__47259\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47267\,
            I => \N__47256\
        );

    \I__11034\ : InMux
    port map (
            O => \N__47266\,
            I => \N__47252\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47265\,
            I => \N__47249\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47262\,
            I => \N__47244\
        );

    \I__11031\ : InMux
    port map (
            O => \N__47259\,
            I => \N__47244\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__47256\,
            I => \N__47241\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47238\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__47252\,
            I => \N__47233\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__47249\,
            I => \N__47233\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__47244\,
            I => \N__47230\
        );

    \I__11025\ : Span12Mux_h
    port map (
            O => \N__47241\,
            I => \N__47227\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__47238\,
            I => \N__47224\
        );

    \I__11023\ : Span12Mux_v
    port map (
            O => \N__47233\,
            I => \N__47221\
        );

    \I__11022\ : Span4Mux_s2_v
    port map (
            O => \N__47230\,
            I => \N__47218\
        );

    \I__11021\ : Odrv12
    port map (
            O => \N__47227\,
            I => \ALU.a5_b_5\
        );

    \I__11020\ : Odrv4
    port map (
            O => \N__47224\,
            I => \ALU.a5_b_5\
        );

    \I__11019\ : Odrv12
    port map (
            O => \N__47221\,
            I => \ALU.a5_b_5\
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__47218\,
            I => \ALU.a5_b_5\
        );

    \I__11017\ : CascadeMux
    port map (
            O => \N__47209\,
            I => \N__47206\
        );

    \I__11016\ : InMux
    port map (
            O => \N__47206\,
            I => \N__47203\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__47203\,
            I => \N__47200\
        );

    \I__11014\ : Odrv12
    port map (
            O => \N__47200\,
            I => \ALU.r0_12_prm_7_5_s1_c_RNOZ0\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47197\,
            I => \N__47191\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47186\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47186\
        );

    \I__11010\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47179\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__47191\,
            I => \N__47176\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__47186\,
            I => \N__47173\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47185\,
            I => \N__47166\
        );

    \I__11006\ : InMux
    port map (
            O => \N__47184\,
            I => \N__47166\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47183\,
            I => \N__47166\
        );

    \I__11004\ : CascadeMux
    port map (
            O => \N__47182\,
            I => \N__47163\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47179\,
            I => \N__47160\
        );

    \I__11002\ : Span4Mux_v
    port map (
            O => \N__47176\,
            I => \N__47153\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__47173\,
            I => \N__47153\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__47166\,
            I => \N__47153\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47150\
        );

    \I__10998\ : Span4Mux_h
    port map (
            O => \N__47160\,
            I => \N__47145\
        );

    \I__10997\ : Span4Mux_v
    port map (
            O => \N__47153\,
            I => \N__47140\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47150\,
            I => \N__47140\
        );

    \I__10995\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47136\
        );

    \I__10994\ : InMux
    port map (
            O => \N__47148\,
            I => \N__47133\
        );

    \I__10993\ : Span4Mux_v
    port map (
            O => \N__47145\,
            I => \N__47128\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__47140\,
            I => \N__47128\
        );

    \I__10991\ : CascadeMux
    port map (
            O => \N__47139\,
            I => \N__47125\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__47136\,
            I => \N__47122\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47133\,
            I => \N__47119\
        );

    \I__10988\ : Span4Mux_h
    port map (
            O => \N__47128\,
            I => \N__47116\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47125\,
            I => \N__47113\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__47122\,
            I => \N__47107\
        );

    \I__10985\ : Span4Mux_v
    port map (
            O => \N__47119\,
            I => \N__47107\
        );

    \I__10984\ : Span4Mux_h
    port map (
            O => \N__47116\,
            I => \N__47102\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__47113\,
            I => \N__47102\
        );

    \I__10982\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47099\
        );

    \I__10981\ : Span4Mux_h
    port map (
            O => \N__47107\,
            I => \N__47096\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__47102\,
            I => \N__47093\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47090\
        );

    \I__10978\ : Span4Mux_h
    port map (
            O => \N__47096\,
            I => \N__47087\
        );

    \I__10977\ : IoSpan4Mux
    port map (
            O => \N__47093\,
            I => \N__47084\
        );

    \I__10976\ : Span4Mux_v
    port map (
            O => \N__47090\,
            I => \N__47081\
        );

    \I__10975\ : Span4Mux_h
    port map (
            O => \N__47087\,
            I => \N__47076\
        );

    \I__10974\ : Span4Mux_s2_h
    port map (
            O => \N__47084\,
            I => \N__47076\
        );

    \I__10973\ : Odrv4
    port map (
            O => \N__47081\,
            I => \ALU.b_14\
        );

    \I__10972\ : Odrv4
    port map (
            O => \N__47076\,
            I => \ALU.b_14\
        );

    \I__10971\ : CascadeMux
    port map (
            O => \N__47071\,
            I => \N__47067\
        );

    \I__10970\ : CascadeMux
    port map (
            O => \N__47070\,
            I => \N__47063\
        );

    \I__10969\ : InMux
    port map (
            O => \N__47067\,
            I => \N__47060\
        );

    \I__10968\ : InMux
    port map (
            O => \N__47066\,
            I => \N__47057\
        );

    \I__10967\ : InMux
    port map (
            O => \N__47063\,
            I => \N__47053\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__47060\,
            I => \N__47047\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47057\,
            I => \N__47042\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47056\,
            I => \N__47037\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__47053\,
            I => \N__47034\
        );

    \I__10962\ : InMux
    port map (
            O => \N__47052\,
            I => \N__47027\
        );

    \I__10961\ : InMux
    port map (
            O => \N__47051\,
            I => \N__47024\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47050\,
            I => \N__47021\
        );

    \I__10959\ : Span4Mux_v
    port map (
            O => \N__47047\,
            I => \N__47018\
        );

    \I__10958\ : InMux
    port map (
            O => \N__47046\,
            I => \N__47015\
        );

    \I__10957\ : InMux
    port map (
            O => \N__47045\,
            I => \N__47012\
        );

    \I__10956\ : Span4Mux_h
    port map (
            O => \N__47042\,
            I => \N__47004\
        );

    \I__10955\ : CascadeMux
    port map (
            O => \N__47041\,
            I => \N__46998\
        );

    \I__10954\ : InMux
    port map (
            O => \N__47040\,
            I => \N__46995\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__47037\,
            I => \N__46992\
        );

    \I__10952\ : Span4Mux_v
    port map (
            O => \N__47034\,
            I => \N__46989\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47033\,
            I => \N__46985\
        );

    \I__10950\ : InMux
    port map (
            O => \N__47032\,
            I => \N__46982\
        );

    \I__10949\ : InMux
    port map (
            O => \N__47031\,
            I => \N__46977\
        );

    \I__10948\ : InMux
    port map (
            O => \N__47030\,
            I => \N__46977\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__47027\,
            I => \N__46974\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__47024\,
            I => \N__46969\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__47021\,
            I => \N__46969\
        );

    \I__10944\ : Span4Mux_v
    port map (
            O => \N__47018\,
            I => \N__46966\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__47015\,
            I => \N__46963\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__47012\,
            I => \N__46960\
        );

    \I__10941\ : InMux
    port map (
            O => \N__47011\,
            I => \N__46956\
        );

    \I__10940\ : InMux
    port map (
            O => \N__47010\,
            I => \N__46949\
        );

    \I__10939\ : InMux
    port map (
            O => \N__47009\,
            I => \N__46949\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47008\,
            I => \N__46949\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47007\,
            I => \N__46946\
        );

    \I__10936\ : Span4Mux_h
    port map (
            O => \N__47004\,
            I => \N__46943\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47003\,
            I => \N__46940\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47002\,
            I => \N__46933\
        );

    \I__10933\ : InMux
    port map (
            O => \N__47001\,
            I => \N__46933\
        );

    \I__10932\ : InMux
    port map (
            O => \N__46998\,
            I => \N__46933\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__46995\,
            I => \N__46930\
        );

    \I__10930\ : Span4Mux_h
    port map (
            O => \N__46992\,
            I => \N__46925\
        );

    \I__10929\ : Span4Mux_v
    port map (
            O => \N__46989\,
            I => \N__46925\
        );

    \I__10928\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46922\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__46985\,
            I => \N__46919\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__46982\,
            I => \N__46910\
        );

    \I__10925\ : LocalMux
    port map (
            O => \N__46977\,
            I => \N__46910\
        );

    \I__10924\ : Span4Mux_v
    port map (
            O => \N__46974\,
            I => \N__46910\
        );

    \I__10923\ : Span4Mux_v
    port map (
            O => \N__46969\,
            I => \N__46910\
        );

    \I__10922\ : Span4Mux_v
    port map (
            O => \N__46966\,
            I => \N__46907\
        );

    \I__10921\ : Span4Mux_s2_h
    port map (
            O => \N__46963\,
            I => \N__46904\
        );

    \I__10920\ : Span4Mux_v
    port map (
            O => \N__46960\,
            I => \N__46901\
        );

    \I__10919\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46898\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__46956\,
            I => \N__46891\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__46949\,
            I => \N__46891\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__46946\,
            I => \N__46891\
        );

    \I__10915\ : Span4Mux_h
    port map (
            O => \N__46943\,
            I => \N__46886\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__46940\,
            I => \N__46886\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__46933\,
            I => \N__46883\
        );

    \I__10912\ : Span4Mux_v
    port map (
            O => \N__46930\,
            I => \N__46870\
        );

    \I__10911\ : Span4Mux_v
    port map (
            O => \N__46925\,
            I => \N__46870\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46922\,
            I => \N__46870\
        );

    \I__10909\ : Span4Mux_h
    port map (
            O => \N__46919\,
            I => \N__46870\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__46910\,
            I => \N__46870\
        );

    \I__10907\ : Span4Mux_h
    port map (
            O => \N__46907\,
            I => \N__46870\
        );

    \I__10906\ : Span4Mux_h
    port map (
            O => \N__46904\,
            I => \N__46867\
        );

    \I__10905\ : Odrv4
    port map (
            O => \N__46901\,
            I => \ALU.a_14\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__46898\,
            I => \ALU.a_14\
        );

    \I__10903\ : Odrv12
    port map (
            O => \N__46891\,
            I => \ALU.a_14\
        );

    \I__10902\ : Odrv4
    port map (
            O => \N__46886\,
            I => \ALU.a_14\
        );

    \I__10901\ : Odrv12
    port map (
            O => \N__46883\,
            I => \ALU.a_14\
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__46870\,
            I => \ALU.a_14\
        );

    \I__10899\ : Odrv4
    port map (
            O => \N__46867\,
            I => \ALU.a_14\
        );

    \I__10898\ : CascadeMux
    port map (
            O => \N__46852\,
            I => \N__46849\
        );

    \I__10897\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46846\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__46846\,
            I => \N__46843\
        );

    \I__10895\ : Span12Mux_s3_v
    port map (
            O => \N__46843\,
            I => \N__46840\
        );

    \I__10894\ : Odrv12
    port map (
            O => \N__46840\,
            I => \ALU.r0_12_prm_7_7_s1_c_RNOZ0\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46834\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__46834\,
            I => \N__46828\
        );

    \I__10891\ : InMux
    port map (
            O => \N__46833\,
            I => \N__46825\
        );

    \I__10890\ : CascadeMux
    port map (
            O => \N__46832\,
            I => \N__46819\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46816\
        );

    \I__10888\ : Span4Mux_v
    port map (
            O => \N__46828\,
            I => \N__46811\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46825\,
            I => \N__46811\
        );

    \I__10886\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46808\
        );

    \I__10885\ : CascadeMux
    port map (
            O => \N__46823\,
            I => \N__46802\
        );

    \I__10884\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46799\
        );

    \I__10883\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46790\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__46816\,
            I => \N__46782\
        );

    \I__10881\ : Span4Mux_h
    port map (
            O => \N__46811\,
            I => \N__46782\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__46808\,
            I => \N__46782\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46807\,
            I => \N__46772\
        );

    \I__10878\ : InMux
    port map (
            O => \N__46806\,
            I => \N__46767\
        );

    \I__10877\ : InMux
    port map (
            O => \N__46805\,
            I => \N__46767\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46802\,
            I => \N__46764\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__46799\,
            I => \N__46761\
        );

    \I__10874\ : InMux
    port map (
            O => \N__46798\,
            I => \N__46758\
        );

    \I__10873\ : InMux
    port map (
            O => \N__46797\,
            I => \N__46755\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46796\,
            I => \N__46751\
        );

    \I__10871\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46737\
        );

    \I__10870\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46737\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46737\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46790\,
            I => \N__46734\
        );

    \I__10867\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46731\
        );

    \I__10866\ : Span4Mux_h
    port map (
            O => \N__46782\,
            I => \N__46728\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46781\,
            I => \N__46723\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46723\
        );

    \I__10863\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46714\
        );

    \I__10862\ : InMux
    port map (
            O => \N__46778\,
            I => \N__46714\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46714\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46714\
        );

    \I__10859\ : CascadeMux
    port map (
            O => \N__46775\,
            I => \N__46711\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__46772\,
            I => \N__46705\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46705\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46764\,
            I => \N__46702\
        );

    \I__10855\ : Span4Mux_v
    port map (
            O => \N__46761\,
            I => \N__46699\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46758\,
            I => \N__46694\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__46755\,
            I => \N__46694\
        );

    \I__10852\ : CascadeMux
    port map (
            O => \N__46754\,
            I => \N__46690\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__46751\,
            I => \N__46687\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46684\
        );

    \I__10849\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46681\
        );

    \I__10848\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46673\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46673\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46746\,
            I => \N__46663\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46663\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46663\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46737\,
            I => \N__46660\
        );

    \I__10842\ : Span4Mux_v
    port map (
            O => \N__46734\,
            I => \N__46655\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46731\,
            I => \N__46655\
        );

    \I__10840\ : Span4Mux_v
    port map (
            O => \N__46728\,
            I => \N__46652\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46723\,
            I => \N__46647\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46647\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46711\,
            I => \N__46644\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46710\,
            I => \N__46641\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__46705\,
            I => \N__46638\
        );

    \I__10834\ : Span4Mux_h
    port map (
            O => \N__46702\,
            I => \N__46631\
        );

    \I__10833\ : Span4Mux_h
    port map (
            O => \N__46699\,
            I => \N__46631\
        );

    \I__10832\ : Span4Mux_s2_v
    port map (
            O => \N__46694\,
            I => \N__46631\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46626\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46690\,
            I => \N__46626\
        );

    \I__10829\ : Span4Mux_s1_h
    port map (
            O => \N__46687\,
            I => \N__46621\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46684\,
            I => \N__46621\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46681\,
            I => \N__46618\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46680\,
            I => \N__46615\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46612\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46609\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__46673\,
            I => \N__46606\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46672\,
            I => \N__46603\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46598\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46598\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46663\,
            I => \N__46595\
        );

    \I__10818\ : Span4Mux_s3_h
    port map (
            O => \N__46660\,
            I => \N__46586\
        );

    \I__10817\ : Span4Mux_s3_h
    port map (
            O => \N__46655\,
            I => \N__46586\
        );

    \I__10816\ : Span4Mux_v
    port map (
            O => \N__46652\,
            I => \N__46586\
        );

    \I__10815\ : Span4Mux_v
    port map (
            O => \N__46647\,
            I => \N__46586\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46575\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46575\
        );

    \I__10812\ : Span4Mux_h
    port map (
            O => \N__46638\,
            I => \N__46575\
        );

    \I__10811\ : Span4Mux_h
    port map (
            O => \N__46631\,
            I => \N__46575\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46626\,
            I => \N__46575\
        );

    \I__10809\ : Span4Mux_h
    port map (
            O => \N__46621\,
            I => \N__46572\
        );

    \I__10808\ : Odrv12
    port map (
            O => \N__46618\,
            I => \ALU.b_1\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__46615\,
            I => \ALU.b_1\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46612\,
            I => \ALU.b_1\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46609\,
            I => \ALU.b_1\
        );

    \I__10804\ : Odrv4
    port map (
            O => \N__46606\,
            I => \ALU.b_1\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__46603\,
            I => \ALU.b_1\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46598\,
            I => \ALU.b_1\
        );

    \I__10801\ : Odrv4
    port map (
            O => \N__46595\,
            I => \ALU.b_1\
        );

    \I__10800\ : Odrv4
    port map (
            O => \N__46586\,
            I => \ALU.b_1\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__46575\,
            I => \ALU.b_1\
        );

    \I__10798\ : Odrv4
    port map (
            O => \N__46572\,
            I => \ALU.b_1\
        );

    \I__10797\ : CascadeMux
    port map (
            O => \N__46549\,
            I => \N__46546\
        );

    \I__10796\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46543\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__46543\,
            I => \N__46540\
        );

    \I__10794\ : Span4Mux_h
    port map (
            O => \N__46540\,
            I => \N__46537\
        );

    \I__10793\ : Odrv4
    port map (
            O => \N__46537\,
            I => \ALU.un14_log_0_i_1\
        );

    \I__10792\ : CascadeMux
    port map (
            O => \N__46534\,
            I => \N__46531\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46528\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46528\,
            I => \ALU.r0_12_prm_5_1_c_RNOZ0Z_0\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46522\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__46522\,
            I => \N__46519\
        );

    \I__10787\ : Span4Mux_v
    port map (
            O => \N__46519\,
            I => \N__46516\
        );

    \I__10786\ : Span4Mux_h
    port map (
            O => \N__46516\,
            I => \N__46513\
        );

    \I__10785\ : Odrv4
    port map (
            O => \N__46513\,
            I => \ALU.rshift_14\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46510\,
            I => \N__46506\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46509\,
            I => \N__46503\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__46506\,
            I => \N__46497\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46503\,
            I => \N__46497\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46494\
        );

    \I__10779\ : Span4Mux_v
    port map (
            O => \N__46497\,
            I => \N__46488\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46494\,
            I => \N__46488\
        );

    \I__10777\ : InMux
    port map (
            O => \N__46493\,
            I => \N__46485\
        );

    \I__10776\ : Span4Mux_v
    port map (
            O => \N__46488\,
            I => \N__46482\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46485\,
            I => \N__46479\
        );

    \I__10774\ : Span4Mux_h
    port map (
            O => \N__46482\,
            I => \N__46474\
        );

    \I__10773\ : Span4Mux_v
    port map (
            O => \N__46479\,
            I => \N__46474\
        );

    \I__10772\ : Odrv4
    port map (
            O => \N__46474\,
            I => \ALU.N_622_1\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46471\,
            I => \N__46468\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46468\,
            I => \ALU.r0_12_prm_8_1_c_RNOZ0\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46465\,
            I => \N__46457\
        );

    \I__10768\ : InMux
    port map (
            O => \N__46464\,
            I => \N__46453\
        );

    \I__10767\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46450\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46447\
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__46461\,
            I => \N__46443\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46440\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46457\,
            I => \N__46437\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46456\,
            I => \N__46434\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__46453\,
            I => \N__46426\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46426\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46447\,
            I => \N__46423\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__46446\,
            I => \N__46419\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46443\,
            I => \N__46416\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__46440\,
            I => \N__46413\
        );

    \I__10755\ : Span4Mux_h
    port map (
            O => \N__46437\,
            I => \N__46409\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__46434\,
            I => \N__46406\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46403\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46432\,
            I => \N__46400\
        );

    \I__10751\ : CascadeMux
    port map (
            O => \N__46431\,
            I => \N__46397\
        );

    \I__10750\ : Span4Mux_v
    port map (
            O => \N__46426\,
            I => \N__46392\
        );

    \I__10749\ : Span4Mux_v
    port map (
            O => \N__46423\,
            I => \N__46392\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46387\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46419\,
            I => \N__46387\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__46416\,
            I => \N__46384\
        );

    \I__10745\ : Span4Mux_v
    port map (
            O => \N__46413\,
            I => \N__46379\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46412\,
            I => \N__46376\
        );

    \I__10743\ : Span4Mux_h
    port map (
            O => \N__46409\,
            I => \N__46372\
        );

    \I__10742\ : Span4Mux_v
    port map (
            O => \N__46406\,
            I => \N__46367\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46403\,
            I => \N__46367\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__46400\,
            I => \N__46364\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46360\
        );

    \I__10738\ : Span4Mux_h
    port map (
            O => \N__46392\,
            I => \N__46355\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__46387\,
            I => \N__46355\
        );

    \I__10736\ : Span4Mux_v
    port map (
            O => \N__46384\,
            I => \N__46352\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46349\
        );

    \I__10734\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46345\
        );

    \I__10733\ : Span4Mux_h
    port map (
            O => \N__46379\,
            I => \N__46340\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__46376\,
            I => \N__46340\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46337\
        );

    \I__10730\ : Span4Mux_h
    port map (
            O => \N__46372\,
            I => \N__46327\
        );

    \I__10729\ : Span4Mux_h
    port map (
            O => \N__46367\,
            I => \N__46327\
        );

    \I__10728\ : Span4Mux_h
    port map (
            O => \N__46364\,
            I => \N__46327\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46324\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__46360\,
            I => \N__46321\
        );

    \I__10725\ : Span4Mux_v
    port map (
            O => \N__46355\,
            I => \N__46318\
        );

    \I__10724\ : Span4Mux_h
    port map (
            O => \N__46352\,
            I => \N__46312\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__46349\,
            I => \N__46309\
        );

    \I__10722\ : CascadeMux
    port map (
            O => \N__46348\,
            I => \N__46304\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46301\
        );

    \I__10720\ : Span4Mux_v
    port map (
            O => \N__46340\,
            I => \N__46298\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__46337\,
            I => \N__46295\
        );

    \I__10718\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46292\
        );

    \I__10717\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46287\
        );

    \I__10716\ : InMux
    port map (
            O => \N__46334\,
            I => \N__46287\
        );

    \I__10715\ : Span4Mux_v
    port map (
            O => \N__46327\,
            I => \N__46284\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__46324\,
            I => \N__46281\
        );

    \I__10713\ : Span4Mux_s2_v
    port map (
            O => \N__46321\,
            I => \N__46276\
        );

    \I__10712\ : Span4Mux_h
    port map (
            O => \N__46318\,
            I => \N__46276\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46317\,
            I => \N__46269\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46316\,
            I => \N__46269\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46315\,
            I => \N__46269\
        );

    \I__10708\ : Span4Mux_v
    port map (
            O => \N__46312\,
            I => \N__46264\
        );

    \I__10707\ : Span4Mux_s2_v
    port map (
            O => \N__46309\,
            I => \N__46264\
        );

    \I__10706\ : InMux
    port map (
            O => \N__46308\,
            I => \N__46261\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46307\,
            I => \N__46256\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46304\,
            I => \N__46256\
        );

    \I__10703\ : Span12Mux_v
    port map (
            O => \N__46301\,
            I => \N__46245\
        );

    \I__10702\ : Sp12to4
    port map (
            O => \N__46298\,
            I => \N__46245\
        );

    \I__10701\ : Span12Mux_s2_v
    port map (
            O => \N__46295\,
            I => \N__46245\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__46292\,
            I => \N__46245\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__46287\,
            I => \N__46245\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__46284\,
            I => \ALU.b_8\
        );

    \I__10697\ : Odrv4
    port map (
            O => \N__46281\,
            I => \ALU.b_8\
        );

    \I__10696\ : Odrv4
    port map (
            O => \N__46276\,
            I => \ALU.b_8\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__46269\,
            I => \ALU.b_8\
        );

    \I__10694\ : Odrv4
    port map (
            O => \N__46264\,
            I => \ALU.b_8\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__46261\,
            I => \ALU.b_8\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__46256\,
            I => \ALU.b_8\
        );

    \I__10691\ : Odrv12
    port map (
            O => \N__46245\,
            I => \ALU.b_8\
        );

    \I__10690\ : CascadeMux
    port map (
            O => \N__46228\,
            I => \N__46224\
        );

    \I__10689\ : CascadeMux
    port map (
            O => \N__46227\,
            I => \N__46221\
        );

    \I__10688\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46211\
        );

    \I__10687\ : InMux
    port map (
            O => \N__46221\,
            I => \N__46211\
        );

    \I__10686\ : InMux
    port map (
            O => \N__46220\,
            I => \N__46208\
        );

    \I__10685\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46205\
        );

    \I__10684\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46201\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__46217\,
            I => \N__46196\
        );

    \I__10682\ : InMux
    port map (
            O => \N__46216\,
            I => \N__46193\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46211\,
            I => \N__46183\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__46208\,
            I => \N__46183\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__46205\,
            I => \N__46174\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46204\,
            I => \N__46169\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__46201\,
            I => \N__46166\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46163\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46157\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46196\,
            I => \N__46154\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46148\
        );

    \I__10672\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46143\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46143\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46140\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__46189\,
            I => \N__46136\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46188\,
            I => \N__46132\
        );

    \I__10667\ : Span4Mux_v
    port map (
            O => \N__46183\,
            I => \N__46129\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46182\,
            I => \N__46126\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46123\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46120\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46179\,
            I => \N__46115\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46115\
        );

    \I__10661\ : InMux
    port map (
            O => \N__46177\,
            I => \N__46112\
        );

    \I__10660\ : Span4Mux_v
    port map (
            O => \N__46174\,
            I => \N__46109\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46104\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46172\,
            I => \N__46104\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__46169\,
            I => \N__46100\
        );

    \I__10656\ : Span4Mux_v
    port map (
            O => \N__46166\,
            I => \N__46097\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46163\,
            I => \N__46094\
        );

    \I__10654\ : InMux
    port map (
            O => \N__46162\,
            I => \N__46091\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46161\,
            I => \N__46086\
        );

    \I__10652\ : InMux
    port map (
            O => \N__46160\,
            I => \N__46086\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__46157\,
            I => \N__46081\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__46154\,
            I => \N__46081\
        );

    \I__10649\ : InMux
    port map (
            O => \N__46153\,
            I => \N__46075\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46075\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46070\
        );

    \I__10646\ : Span4Mux_h
    port map (
            O => \N__46148\,
            I => \N__46063\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46063\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__46140\,
            I => \N__46063\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46056\
        );

    \I__10642\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46056\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46056\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__46132\,
            I => \N__46052\
        );

    \I__10639\ : Span4Mux_h
    port map (
            O => \N__46129\,
            I => \N__46047\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__46126\,
            I => \N__46047\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46123\,
            I => \N__46036\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__46120\,
            I => \N__46036\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__46115\,
            I => \N__46036\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__46112\,
            I => \N__46036\
        );

    \I__10633\ : Sp12to4
    port map (
            O => \N__46109\,
            I => \N__46036\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46104\,
            I => \N__46033\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46103\,
            I => \N__46030\
        );

    \I__10630\ : Span4Mux_s1_v
    port map (
            O => \N__46100\,
            I => \N__46027\
        );

    \I__10629\ : Span4Mux_h
    port map (
            O => \N__46097\,
            I => \N__46016\
        );

    \I__10628\ : Span4Mux_v
    port map (
            O => \N__46094\,
            I => \N__46016\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46091\,
            I => \N__46016\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__46016\
        );

    \I__10625\ : Span4Mux_v
    port map (
            O => \N__46081\,
            I => \N__46016\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46013\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46010\
        );

    \I__10622\ : CascadeMux
    port map (
            O => \N__46074\,
            I => \N__46005\
        );

    \I__10621\ : CascadeMux
    port map (
            O => \N__46073\,
            I => \N__46002\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__46070\,
            I => \N__45999\
        );

    \I__10619\ : Span4Mux_h
    port map (
            O => \N__46063\,
            I => \N__45996\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__46056\,
            I => \N__45993\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46055\,
            I => \N__45990\
        );

    \I__10616\ : Span4Mux_h
    port map (
            O => \N__46052\,
            I => \N__45983\
        );

    \I__10615\ : Span4Mux_h
    port map (
            O => \N__46047\,
            I => \N__45983\
        );

    \I__10614\ : Span12Mux_h
    port map (
            O => \N__46036\,
            I => \N__45980\
        );

    \I__10613\ : Span4Mux_v
    port map (
            O => \N__46033\,
            I => \N__45971\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__46030\,
            I => \N__45971\
        );

    \I__10611\ : Span4Mux_v
    port map (
            O => \N__46027\,
            I => \N__45971\
        );

    \I__10610\ : Span4Mux_h
    port map (
            O => \N__46016\,
            I => \N__45971\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__46013\,
            I => \N__45966\
        );

    \I__10608\ : Span4Mux_h
    port map (
            O => \N__46010\,
            I => \N__45966\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46009\,
            I => \N__45957\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45957\
        );

    \I__10605\ : InMux
    port map (
            O => \N__46005\,
            I => \N__45957\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45957\
        );

    \I__10603\ : Span12Mux_s5_v
    port map (
            O => \N__45999\,
            I => \N__45954\
        );

    \I__10602\ : Span4Mux_h
    port map (
            O => \N__45996\,
            I => \N__45947\
        );

    \I__10601\ : Span4Mux_h
    port map (
            O => \N__45993\,
            I => \N__45947\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__45990\,
            I => \N__45947\
        );

    \I__10599\ : InMux
    port map (
            O => \N__45989\,
            I => \N__45944\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45988\,
            I => \N__45941\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__45983\,
            I => \ALU.a_8\
        );

    \I__10596\ : Odrv12
    port map (
            O => \N__45980\,
            I => \ALU.a_8\
        );

    \I__10595\ : Odrv4
    port map (
            O => \N__45971\,
            I => \ALU.a_8\
        );

    \I__10594\ : Odrv4
    port map (
            O => \N__45966\,
            I => \ALU.a_8\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__45957\,
            I => \ALU.a_8\
        );

    \I__10592\ : Odrv12
    port map (
            O => \N__45954\,
            I => \ALU.a_8\
        );

    \I__10591\ : Odrv4
    port map (
            O => \N__45947\,
            I => \ALU.a_8\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45944\,
            I => \ALU.a_8\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__45941\,
            I => \ALU.a_8\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__45922\,
            I => \N__45919\
        );

    \I__10587\ : InMux
    port map (
            O => \N__45919\,
            I => \N__45916\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__45916\,
            I => \N__45913\
        );

    \I__10585\ : Odrv4
    port map (
            O => \N__45913\,
            I => \ALU.r0_12_prm_7_8_s1_c_RNOZ0\
        );

    \I__10584\ : CascadeMux
    port map (
            O => \N__45910\,
            I => \N__45907\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45907\,
            I => \N__45904\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__45904\,
            I => \N__45901\
        );

    \I__10581\ : Span4Mux_h
    port map (
            O => \N__45901\,
            I => \N__45898\
        );

    \I__10580\ : Odrv4
    port map (
            O => \N__45898\,
            I => \ALU.r0_12_prm_7_9_s0_c_RNOZ0\
        );

    \I__10579\ : CEMux
    port map (
            O => \N__45895\,
            I => \N__45892\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__45892\,
            I => \N__45889\
        );

    \I__10577\ : Span4Mux_v
    port map (
            O => \N__45889\,
            I => \N__45885\
        );

    \I__10576\ : CEMux
    port map (
            O => \N__45888\,
            I => \N__45882\
        );

    \I__10575\ : Span4Mux_h
    port map (
            O => \N__45885\,
            I => \N__45879\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__45882\,
            I => \N__45876\
        );

    \I__10573\ : Span4Mux_h
    port map (
            O => \N__45879\,
            I => \N__45873\
        );

    \I__10572\ : Span4Mux_v
    port map (
            O => \N__45876\,
            I => \N__45870\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__45873\,
            I => \N__45867\
        );

    \I__10570\ : Span4Mux_h
    port map (
            O => \N__45870\,
            I => \N__45864\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__45867\,
            I => \N__45861\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__45864\,
            I => \N__45858\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__45861\,
            I => \ALU.un1_yindexZ0Z_1\
        );

    \I__10566\ : Odrv4
    port map (
            O => \N__45858\,
            I => \ALU.un1_yindexZ0Z_1\
        );

    \I__10565\ : CEMux
    port map (
            O => \N__45853\,
            I => \N__45850\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45850\,
            I => \N__45847\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__45847\,
            I => \N__45843\
        );

    \I__10562\ : CEMux
    port map (
            O => \N__45846\,
            I => \N__45839\
        );

    \I__10561\ : Span4Mux_v
    port map (
            O => \N__45843\,
            I => \N__45836\
        );

    \I__10560\ : CEMux
    port map (
            O => \N__45842\,
            I => \N__45833\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__45839\,
            I => \N__45830\
        );

    \I__10558\ : Span4Mux_h
    port map (
            O => \N__45836\,
            I => \N__45827\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__45833\,
            I => \N__45824\
        );

    \I__10556\ : Span4Mux_v
    port map (
            O => \N__45830\,
            I => \N__45821\
        );

    \I__10555\ : Span4Mux_h
    port map (
            O => \N__45827\,
            I => \N__45818\
        );

    \I__10554\ : Span12Mux_h
    port map (
            O => \N__45824\,
            I => \N__45815\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__45821\,
            I => \N__45812\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__45818\,
            I => \ALU.un1_yindexZ0Z_2\
        );

    \I__10551\ : Odrv12
    port map (
            O => \N__45815\,
            I => \ALU.un1_yindexZ0Z_2\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__45812\,
            I => \ALU.un1_yindexZ0Z_2\
        );

    \I__10549\ : CEMux
    port map (
            O => \N__45805\,
            I => \N__45802\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__45802\,
            I => \N__45798\
        );

    \I__10547\ : CEMux
    port map (
            O => \N__45801\,
            I => \N__45795\
        );

    \I__10546\ : Span4Mux_v
    port map (
            O => \N__45798\,
            I => \N__45792\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45789\
        );

    \I__10544\ : Span4Mux_h
    port map (
            O => \N__45792\,
            I => \N__45786\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__45789\,
            I => \N__45783\
        );

    \I__10542\ : Span4Mux_h
    port map (
            O => \N__45786\,
            I => \N__45780\
        );

    \I__10541\ : Span4Mux_h
    port map (
            O => \N__45783\,
            I => \N__45777\
        );

    \I__10540\ : Span4Mux_v
    port map (
            O => \N__45780\,
            I => \N__45774\
        );

    \I__10539\ : Span4Mux_h
    port map (
            O => \N__45777\,
            I => \N__45771\
        );

    \I__10538\ : Odrv4
    port map (
            O => \N__45774\,
            I => \ALU.un1_yindexZ0Z_3\
        );

    \I__10537\ : Odrv4
    port map (
            O => \N__45771\,
            I => \ALU.un1_yindexZ0Z_3\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45766\,
            I => \N__45762\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45765\,
            I => \N__45759\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__45762\,
            I => \N__45756\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__45759\,
            I => \N__45753\
        );

    \I__10532\ : Span4Mux_v
    port map (
            O => \N__45756\,
            I => \N__45748\
        );

    \I__10531\ : Span4Mux_h
    port map (
            O => \N__45753\,
            I => \N__45748\
        );

    \I__10530\ : Span4Mux_v
    port map (
            O => \N__45748\,
            I => \N__45745\
        );

    \I__10529\ : Odrv4
    port map (
            O => \N__45745\,
            I => \ALU.r4_RNI8B628_0Z0Z_5\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__45742\,
            I => \N__45739\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45739\,
            I => \N__45736\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__45736\,
            I => \ALU.r0_12_prm_5_5_s1_c_RNOZ0\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45733\,
            I => \N__45730\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__45730\,
            I => \N__45727\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__45727\,
            I => \N__45724\
        );

    \I__10522\ : Odrv4
    port map (
            O => \N__45724\,
            I => \ALU.r0_12_prm_4_5_s1_c_RNOZ0\
        );

    \I__10521\ : CascadeMux
    port map (
            O => \N__45721\,
            I => \N__45718\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45718\,
            I => \N__45715\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__45715\,
            I => \N__45711\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45708\
        );

    \I__10517\ : Span4Mux_h
    port map (
            O => \N__45711\,
            I => \N__45705\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__45708\,
            I => \ALU.a_i_5\
        );

    \I__10515\ : Odrv4
    port map (
            O => \N__45705\,
            I => \ALU.a_i_5\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45700\,
            I => \N__45697\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__45697\,
            I => \N__45694\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__45694\,
            I => \ALU.r0_12_prm_2_5_s1_c_RNOZ0\
        );

    \I__10511\ : CascadeMux
    port map (
            O => \N__45691\,
            I => \N__45688\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45688\,
            I => \N__45683\
        );

    \I__10509\ : InMux
    port map (
            O => \N__45687\,
            I => \N__45680\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45686\,
            I => \N__45677\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__45683\,
            I => \N__45674\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__45680\,
            I => \N__45670\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__45677\,
            I => \N__45667\
        );

    \I__10504\ : Span4Mux_v
    port map (
            O => \N__45674\,
            I => \N__45664\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45661\
        );

    \I__10502\ : Span4Mux_h
    port map (
            O => \N__45670\,
            I => \N__45658\
        );

    \I__10501\ : Span4Mux_h
    port map (
            O => \N__45667\,
            I => \N__45655\
        );

    \I__10500\ : Sp12to4
    port map (
            O => \N__45664\,
            I => \N__45650\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__45661\,
            I => \N__45650\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__45658\,
            I => \ALU.un2_addsub_cry_4_c_RNILPG3DZ0\
        );

    \I__10497\ : Odrv4
    port map (
            O => \N__45655\,
            I => \ALU.un2_addsub_cry_4_c_RNILPG3DZ0\
        );

    \I__10496\ : Odrv12
    port map (
            O => \N__45650\,
            I => \ALU.un2_addsub_cry_4_c_RNILPG3DZ0\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45640\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45640\,
            I => \ALU.r0_12_prm_1_5_s1_c_RNOZ0\
        );

    \I__10493\ : CascadeMux
    port map (
            O => \N__45637\,
            I => \N__45632\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45636\,
            I => \N__45629\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45635\,
            I => \N__45626\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45622\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__45629\,
            I => \N__45619\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__45626\,
            I => \N__45616\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45613\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__45622\,
            I => \N__45610\
        );

    \I__10485\ : Span4Mux_h
    port map (
            O => \N__45619\,
            I => \N__45607\
        );

    \I__10484\ : Span4Mux_h
    port map (
            O => \N__45616\,
            I => \N__45604\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__45613\,
            I => \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88\
        );

    \I__10482\ : Odrv12
    port map (
            O => \N__45610\,
            I => \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88\
        );

    \I__10481\ : Odrv4
    port map (
            O => \N__45607\,
            I => \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88\
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__45604\,
            I => \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45595\,
            I => \ALU.r0_12_s1_5\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45589\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45589\,
            I => \N__45586\
        );

    \I__10476\ : Span4Mux_h
    port map (
            O => \N__45586\,
            I => \N__45583\
        );

    \I__10475\ : Odrv4
    port map (
            O => \N__45583\,
            I => \ALU.r0_12_s1_5_THRU_CO\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__45580\,
            I => \N__45577\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45574\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45574\,
            I => \N__45571\
        );

    \I__10471\ : Span4Mux_h
    port map (
            O => \N__45571\,
            I => \N__45568\
        );

    \I__10470\ : Odrv4
    port map (
            O => \N__45568\,
            I => \ALU.r0_12_prm_5_8_s1_c_RNOZ0\
        );

    \I__10469\ : CascadeMux
    port map (
            O => \N__45565\,
            I => \N__45562\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45559\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45559\,
            I => \N__45556\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__45556\,
            I => \N__45553\
        );

    \I__10465\ : Span4Mux_h
    port map (
            O => \N__45553\,
            I => \N__45550\
        );

    \I__10464\ : Span4Mux_h
    port map (
            O => \N__45550\,
            I => \N__45547\
        );

    \I__10463\ : Odrv4
    port map (
            O => \N__45547\,
            I => \ALU.r0_12_prm_5_10_s0_c_RNOZ0\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45540\
        );

    \I__10461\ : CascadeMux
    port map (
            O => \N__45543\,
            I => \N__45537\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45540\,
            I => \N__45534\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45531\
        );

    \I__10458\ : Span4Mux_h
    port map (
            O => \N__45534\,
            I => \N__45528\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__45531\,
            I => \N__45525\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__45528\,
            I => \N__45520\
        );

    \I__10455\ : Span4Mux_v
    port map (
            O => \N__45525\,
            I => \N__45520\
        );

    \I__10454\ : Span4Mux_v
    port map (
            O => \N__45520\,
            I => \N__45517\
        );

    \I__10453\ : Odrv4
    port map (
            O => \N__45517\,
            I => \ALU.un14_log_0_i_9\
        );

    \I__10452\ : CascadeMux
    port map (
            O => \N__45514\,
            I => \N__45507\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__45513\,
            I => \N__45501\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45497\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45491\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45488\
        );

    \I__10447\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45485\
        );

    \I__10446\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45480\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45476\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45473\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45470\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45467\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__45497\,
            I => \N__45464\
        );

    \I__10440\ : CascadeMux
    port map (
            O => \N__45496\,
            I => \N__45458\
        );

    \I__10439\ : CascadeMux
    port map (
            O => \N__45495\,
            I => \N__45455\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45494\,
            I => \N__45448\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__45491\,
            I => \N__45445\
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__45488\,
            I => \N__45440\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__45485\,
            I => \N__45440\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45435\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45483\,
            I => \N__45435\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45480\,
            I => \N__45432\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45479\,
            I => \N__45429\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45476\,
            I => \N__45426\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45473\,
            I => \N__45419\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45470\,
            I => \N__45419\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45467\,
            I => \N__45419\
        );

    \I__10426\ : Span4Mux_h
    port map (
            O => \N__45464\,
            I => \N__45415\
        );

    \I__10425\ : InMux
    port map (
            O => \N__45463\,
            I => \N__45412\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45409\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45406\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45401\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45398\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45395\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45392\
        );

    \I__10418\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45388\
        );

    \I__10417\ : CascadeMux
    port map (
            O => \N__45451\,
            I => \N__45385\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__45448\,
            I => \N__45380\
        );

    \I__10415\ : Span4Mux_h
    port map (
            O => \N__45445\,
            I => \N__45373\
        );

    \I__10414\ : Span4Mux_v
    port map (
            O => \N__45440\,
            I => \N__45373\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__45435\,
            I => \N__45373\
        );

    \I__10412\ : Span4Mux_v
    port map (
            O => \N__45432\,
            I => \N__45370\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45429\,
            I => \N__45367\
        );

    \I__10410\ : Span4Mux_v
    port map (
            O => \N__45426\,
            I => \N__45362\
        );

    \I__10409\ : Span4Mux_s1_v
    port map (
            O => \N__45419\,
            I => \N__45362\
        );

    \I__10408\ : CascadeMux
    port map (
            O => \N__45418\,
            I => \N__45357\
        );

    \I__10407\ : Sp12to4
    port map (
            O => \N__45415\,
            I => \N__45354\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__45412\,
            I => \N__45349\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__45409\,
            I => \N__45349\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45406\,
            I => \N__45346\
        );

    \I__10403\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45341\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45404\,
            I => \N__45341\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45401\,
            I => \N__45334\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__45398\,
            I => \N__45334\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__45395\,
            I => \N__45334\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45392\,
            I => \N__45331\
        );

    \I__10397\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45328\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__45388\,
            I => \N__45325\
        );

    \I__10395\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45322\
        );

    \I__10394\ : InMux
    port map (
            O => \N__45384\,
            I => \N__45317\
        );

    \I__10393\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45317\
        );

    \I__10392\ : Span4Mux_s2_v
    port map (
            O => \N__45380\,
            I => \N__45312\
        );

    \I__10391\ : Span4Mux_v
    port map (
            O => \N__45373\,
            I => \N__45312\
        );

    \I__10390\ : Span4Mux_h
    port map (
            O => \N__45370\,
            I => \N__45305\
        );

    \I__10389\ : Span4Mux_v
    port map (
            O => \N__45367\,
            I => \N__45305\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__45362\,
            I => \N__45305\
        );

    \I__10387\ : InMux
    port map (
            O => \N__45361\,
            I => \N__45300\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45360\,
            I => \N__45300\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45357\,
            I => \N__45297\
        );

    \I__10384\ : Span12Mux_v
    port map (
            O => \N__45354\,
            I => \N__45288\
        );

    \I__10383\ : Span12Mux_v
    port map (
            O => \N__45349\,
            I => \N__45288\
        );

    \I__10382\ : Span12Mux_s2_h
    port map (
            O => \N__45346\,
            I => \N__45288\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__45341\,
            I => \N__45288\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__45334\,
            I => \N__45285\
        );

    \I__10379\ : Odrv12
    port map (
            O => \N__45331\,
            I => \ALU.a_5\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45328\,
            I => \ALU.a_5\
        );

    \I__10377\ : Odrv4
    port map (
            O => \N__45325\,
            I => \ALU.a_5\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45322\,
            I => \ALU.a_5\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__45317\,
            I => \ALU.a_5\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45312\,
            I => \ALU.a_5\
        );

    \I__10373\ : Odrv4
    port map (
            O => \N__45305\,
            I => \ALU.a_5\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45300\,
            I => \ALU.a_5\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__45297\,
            I => \ALU.a_5\
        );

    \I__10370\ : Odrv12
    port map (
            O => \N__45288\,
            I => \ALU.a_5\
        );

    \I__10369\ : Odrv4
    port map (
            O => \N__45285\,
            I => \ALU.a_5\
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__45262\,
            I => \N__45254\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45251\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45260\,
            I => \N__45246\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45259\,
            I => \N__45243\
        );

    \I__10364\ : CascadeMux
    port map (
            O => \N__45258\,
            I => \N__45240\
        );

    \I__10363\ : CascadeMux
    port map (
            O => \N__45257\,
            I => \N__45237\
        );

    \I__10362\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45234\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__45251\,
            I => \N__45226\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45223\
        );

    \I__10359\ : CascadeMux
    port map (
            O => \N__45249\,
            I => \N__45219\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__45246\,
            I => \N__45215\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__45243\,
            I => \N__45212\
        );

    \I__10356\ : InMux
    port map (
            O => \N__45240\,
            I => \N__45207\
        );

    \I__10355\ : InMux
    port map (
            O => \N__45237\,
            I => \N__45207\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__45234\,
            I => \N__45202\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45196\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45196\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45191\
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__45230\,
            I => \N__45185\
        );

    \I__10349\ : CascadeMux
    port map (
            O => \N__45229\,
            I => \N__45182\
        );

    \I__10348\ : Span4Mux_v
    port map (
            O => \N__45226\,
            I => \N__45176\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__45223\,
            I => \N__45173\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45170\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45219\,
            I => \N__45167\
        );

    \I__10344\ : InMux
    port map (
            O => \N__45218\,
            I => \N__45164\
        );

    \I__10343\ : Span4Mux_v
    port map (
            O => \N__45215\,
            I => \N__45159\
        );

    \I__10342\ : Span4Mux_h
    port map (
            O => \N__45212\,
            I => \N__45159\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__45207\,
            I => \N__45156\
        );

    \I__10340\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45151\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45205\,
            I => \N__45151\
        );

    \I__10338\ : Span4Mux_v
    port map (
            O => \N__45202\,
            I => \N__45148\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45145\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__45196\,
            I => \N__45142\
        );

    \I__10335\ : InMux
    port map (
            O => \N__45195\,
            I => \N__45137\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45137\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__45191\,
            I => \N__45134\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45129\
        );

    \I__10331\ : InMux
    port map (
            O => \N__45189\,
            I => \N__45129\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45188\,
            I => \N__45121\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45185\,
            I => \N__45121\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45121\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45181\,
            I => \N__45118\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45115\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45179\,
            I => \N__45112\
        );

    \I__10324\ : Span4Mux_h
    port map (
            O => \N__45176\,
            I => \N__45107\
        );

    \I__10323\ : Span4Mux_v
    port map (
            O => \N__45173\,
            I => \N__45107\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45170\,
            I => \N__45103\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__45167\,
            I => \N__45100\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45164\,
            I => \N__45097\
        );

    \I__10319\ : Span4Mux_h
    port map (
            O => \N__45159\,
            I => \N__45094\
        );

    \I__10318\ : Span4Mux_h
    port map (
            O => \N__45156\,
            I => \N__45089\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__45151\,
            I => \N__45089\
        );

    \I__10316\ : Span4Mux_h
    port map (
            O => \N__45148\,
            I => \N__45086\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__45145\,
            I => \N__45081\
        );

    \I__10314\ : Span4Mux_s0_v
    port map (
            O => \N__45142\,
            I => \N__45081\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45137\,
            I => \N__45078\
        );

    \I__10312\ : Span4Mux_h
    port map (
            O => \N__45134\,
            I => \N__45073\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45129\,
            I => \N__45073\
        );

    \I__10310\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45070\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__45121\,
            I => \N__45063\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__45118\,
            I => \N__45063\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__45115\,
            I => \N__45063\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__45112\,
            I => \N__45060\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__45107\,
            I => \N__45057\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45106\,
            I => \N__45054\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__45103\,
            I => \N__45047\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__45100\,
            I => \N__45047\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__45097\,
            I => \N__45047\
        );

    \I__10300\ : Span4Mux_h
    port map (
            O => \N__45094\,
            I => \N__45042\
        );

    \I__10299\ : Span4Mux_v
    port map (
            O => \N__45089\,
            I => \N__45042\
        );

    \I__10298\ : Span4Mux_h
    port map (
            O => \N__45086\,
            I => \N__45035\
        );

    \I__10297\ : Span4Mux_v
    port map (
            O => \N__45081\,
            I => \N__45035\
        );

    \I__10296\ : Span4Mux_h
    port map (
            O => \N__45078\,
            I => \N__45035\
        );

    \I__10295\ : Span4Mux_h
    port map (
            O => \N__45073\,
            I => \N__45028\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__45070\,
            I => \N__45028\
        );

    \I__10293\ : Span4Mux_s2_v
    port map (
            O => \N__45063\,
            I => \N__45028\
        );

    \I__10292\ : Odrv12
    port map (
            O => \N__45060\,
            I => \ALU.b_5\
        );

    \I__10291\ : Odrv4
    port map (
            O => \N__45057\,
            I => \ALU.b_5\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__45054\,
            I => \ALU.b_5\
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__45047\,
            I => \ALU.b_5\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__45042\,
            I => \ALU.b_5\
        );

    \I__10287\ : Odrv4
    port map (
            O => \N__45035\,
            I => \ALU.b_5\
        );

    \I__10286\ : Odrv4
    port map (
            O => \N__45028\,
            I => \ALU.b_5\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45013\,
            I => \N__45009\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45012\,
            I => \N__45006\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__45009\,
            I => \N__45002\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__45006\,
            I => \N__44998\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44995\
        );

    \I__10280\ : Span4Mux_h
    port map (
            O => \N__45002\,
            I => \N__44992\
        );

    \I__10279\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44989\
        );

    \I__10278\ : Span4Mux_h
    port map (
            O => \N__44998\,
            I => \N__44986\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__44995\,
            I => \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__44992\,
            I => \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__44989\,
            I => \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8\
        );

    \I__10274\ : Odrv4
    port map (
            O => \N__44986\,
            I => \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8\
        );

    \I__10273\ : CascadeMux
    port map (
            O => \N__44977\,
            I => \N__44974\
        );

    \I__10272\ : InMux
    port map (
            O => \N__44974\,
            I => \N__44971\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__44971\,
            I => \N__44968\
        );

    \I__10270\ : Odrv4
    port map (
            O => \N__44968\,
            I => \ALU.r0_12_prm_1_7_s1_c_RNOZ0\
        );

    \I__10269\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44962\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44962\,
            I => \ALU.r0_12_prm_8_5_s1_c_RNOZ0Z_1\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44956\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__44956\,
            I => \ALU.r0_12_prm_8_5_s1_c_RNOZ0\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44950\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__44950\,
            I => \N__44947\
        );

    \I__10263\ : Odrv12
    port map (
            O => \N__44947\,
            I => \ALU.r0_12_prm_6_5_s1_c_RNOZ0\
        );

    \I__10262\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44941\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__44941\,
            I => \N__44937\
        );

    \I__10260\ : CascadeMux
    port map (
            O => \N__44940\,
            I => \N__44934\
        );

    \I__10259\ : Span4Mux_v
    port map (
            O => \N__44937\,
            I => \N__44931\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44928\
        );

    \I__10257\ : Span4Mux_h
    port map (
            O => \N__44931\,
            I => \N__44925\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__44928\,
            I => \N__44922\
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__44925\,
            I => \ALU.un14_log_0_i_5\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__44922\,
            I => \ALU.un14_log_0_i_5\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44917\,
            I => \ALU.r0_12_s1_7\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44911\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__44911\,
            I => \N__44908\
        );

    \I__10250\ : Span4Mux_h
    port map (
            O => \N__44908\,
            I => \N__44905\
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__44905\,
            I => \ALU.r0_12_s1_7_THRU_CO\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44899\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44896\
        );

    \I__10246\ : Span4Mux_h
    port map (
            O => \N__44896\,
            I => \N__44893\
        );

    \I__10245\ : Span4Mux_h
    port map (
            O => \N__44893\,
            I => \N__44890\
        );

    \I__10244\ : Span4Mux_v
    port map (
            O => \N__44890\,
            I => \N__44885\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44882\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44879\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__44885\,
            I => \ALU.r5_RNISMSV4Z0Z_15\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__44882\,
            I => \ALU.r5_RNISMSV4Z0Z_15\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__44879\,
            I => \ALU.r5_RNISMSV4Z0Z_15\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44869\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__44869\,
            I => \N__44866\
        );

    \I__10236\ : Span4Mux_h
    port map (
            O => \N__44866\,
            I => \N__44863\
        );

    \I__10235\ : Span4Mux_h
    port map (
            O => \N__44863\,
            I => \N__44860\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__44860\,
            I => \ALU.rshift_15_ns_1_3\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44857\,
            I => \N__44854\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__44854\,
            I => \N__44851\
        );

    \I__10231\ : Span4Mux_h
    port map (
            O => \N__44851\,
            I => \N__44848\
        );

    \I__10230\ : Span4Mux_v
    port map (
            O => \N__44848\,
            I => \N__44845\
        );

    \I__10229\ : Span4Mux_v
    port map (
            O => \N__44845\,
            I => \N__44840\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44837\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44843\,
            I => \N__44834\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__44840\,
            I => \ALU.r5_RNI465TIZ0Z_13\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__44837\,
            I => \ALU.r5_RNI465TIZ0Z_13\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__44834\,
            I => \ALU.r5_RNI465TIZ0Z_13\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44824\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__44824\,
            I => \N__44820\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44823\,
            I => \N__44817\
        );

    \I__10220\ : Span4Mux_v
    port map (
            O => \N__44820\,
            I => \N__44814\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__44817\,
            I => \N__44811\
        );

    \I__10218\ : Odrv4
    port map (
            O => \N__44814\,
            I => \ALU.r4_RNIF01FKZ0Z_2\
        );

    \I__10217\ : Odrv4
    port map (
            O => \N__44811\,
            I => \ALU.r4_RNIF01FKZ0Z_2\
        );

    \I__10216\ : CascadeMux
    port map (
            O => \N__44806\,
            I => \N__44802\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44798\
        );

    \I__10214\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44794\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44801\,
            I => \N__44791\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44798\,
            I => \N__44785\
        );

    \I__10211\ : InMux
    port map (
            O => \N__44797\,
            I => \N__44780\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44794\,
            I => \N__44777\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__44791\,
            I => \N__44773\
        );

    \I__10208\ : InMux
    port map (
            O => \N__44790\,
            I => \N__44770\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44767\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44760\
        );

    \I__10205\ : Span4Mux_v
    port map (
            O => \N__44785\,
            I => \N__44757\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44784\,
            I => \N__44754\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44783\,
            I => \N__44751\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__44780\,
            I => \N__44745\
        );

    \I__10201\ : Span4Mux_v
    port map (
            O => \N__44777\,
            I => \N__44745\
        );

    \I__10200\ : InMux
    port map (
            O => \N__44776\,
            I => \N__44742\
        );

    \I__10199\ : Span4Mux_v
    port map (
            O => \N__44773\,
            I => \N__44739\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__44770\,
            I => \N__44736\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44767\,
            I => \N__44733\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44730\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44727\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44724\
        );

    \I__10193\ : CascadeMux
    port map (
            O => \N__44763\,
            I => \N__44720\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44712\
        );

    \I__10191\ : Sp12to4
    port map (
            O => \N__44757\,
            I => \N__44712\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__44754\,
            I => \N__44712\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__44751\,
            I => \N__44709\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44750\,
            I => \N__44706\
        );

    \I__10187\ : Span4Mux_v
    port map (
            O => \N__44745\,
            I => \N__44701\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__44742\,
            I => \N__44698\
        );

    \I__10185\ : Span4Mux_h
    port map (
            O => \N__44739\,
            I => \N__44691\
        );

    \I__10184\ : Span4Mux_s2_v
    port map (
            O => \N__44736\,
            I => \N__44691\
        );

    \I__10183\ : Span4Mux_h
    port map (
            O => \N__44733\,
            I => \N__44691\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44688\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__44727\,
            I => \N__44685\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__44724\,
            I => \N__44682\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44723\,
            I => \N__44679\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44670\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44670\
        );

    \I__10176\ : Span12Mux_h
    port map (
            O => \N__44712\,
            I => \N__44667\
        );

    \I__10175\ : Span4Mux_s3_h
    port map (
            O => \N__44709\,
            I => \N__44664\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44706\,
            I => \N__44661\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44705\,
            I => \N__44656\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44656\
        );

    \I__10171\ : Span4Mux_h
    port map (
            O => \N__44701\,
            I => \N__44645\
        );

    \I__10170\ : Span4Mux_v
    port map (
            O => \N__44698\,
            I => \N__44645\
        );

    \I__10169\ : Span4Mux_h
    port map (
            O => \N__44691\,
            I => \N__44645\
        );

    \I__10168\ : Span4Mux_s2_h
    port map (
            O => \N__44688\,
            I => \N__44645\
        );

    \I__10167\ : Span4Mux_s2_v
    port map (
            O => \N__44685\,
            I => \N__44645\
        );

    \I__10166\ : Span12Mux_h
    port map (
            O => \N__44682\,
            I => \N__44640\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__44679\,
            I => \N__44640\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44678\,
            I => \N__44631\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44631\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44631\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44675\,
            I => \N__44631\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__44670\,
            I => \N__44628\
        );

    \I__10159\ : Odrv12
    port map (
            O => \N__44667\,
            I => \ALU.b_7\
        );

    \I__10158\ : Odrv4
    port map (
            O => \N__44664\,
            I => \ALU.b_7\
        );

    \I__10157\ : Odrv4
    port map (
            O => \N__44661\,
            I => \ALU.b_7\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44656\,
            I => \ALU.b_7\
        );

    \I__10155\ : Odrv4
    port map (
            O => \N__44645\,
            I => \ALU.b_7\
        );

    \I__10154\ : Odrv12
    port map (
            O => \N__44640\,
            I => \ALU.b_7\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44631\,
            I => \ALU.b_7\
        );

    \I__10152\ : Odrv12
    port map (
            O => \N__44628\,
            I => \ALU.b_7\
        );

    \I__10151\ : CascadeMux
    port map (
            O => \N__44611\,
            I => \N__44607\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44604\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44607\,
            I => \N__44597\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__44604\,
            I => \N__44590\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44603\,
            I => \N__44585\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44602\,
            I => \N__44582\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44601\,
            I => \N__44579\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44576\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__44597\,
            I => \N__44573\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44570\
        );

    \I__10141\ : InMux
    port map (
            O => \N__44595\,
            I => \N__44567\
        );

    \I__10140\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44564\
        );

    \I__10139\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44561\
        );

    \I__10138\ : Span4Mux_v
    port map (
            O => \N__44590\,
            I => \N__44558\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44553\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44553\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__44585\,
            I => \N__44546\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__44582\,
            I => \N__44539\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44579\,
            I => \N__44532\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44576\,
            I => \N__44532\
        );

    \I__10131\ : Span4Mux_v
    port map (
            O => \N__44573\,
            I => \N__44526\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__44570\,
            I => \N__44523\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44567\,
            I => \N__44520\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44509\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__44561\,
            I => \N__44509\
        );

    \I__10126\ : Span4Mux_h
    port map (
            O => \N__44558\,
            I => \N__44509\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__44553\,
            I => \N__44509\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44506\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44501\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44550\,
            I => \N__44501\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44549\,
            I => \N__44498\
        );

    \I__10120\ : Span4Mux_h
    port map (
            O => \N__44546\,
            I => \N__44495\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44490\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44544\,
            I => \N__44490\
        );

    \I__10117\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44484\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44481\
        );

    \I__10115\ : Span4Mux_v
    port map (
            O => \N__44539\,
            I => \N__44478\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44473\
        );

    \I__10113\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44473\
        );

    \I__10112\ : Span4Mux_v
    port map (
            O => \N__44532\,
            I => \N__44470\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44531\,
            I => \N__44465\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44530\,
            I => \N__44465\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44529\,
            I => \N__44462\
        );

    \I__10108\ : Span4Mux_h
    port map (
            O => \N__44526\,
            I => \N__44455\
        );

    \I__10107\ : Span4Mux_v
    port map (
            O => \N__44523\,
            I => \N__44455\
        );

    \I__10106\ : Span4Mux_v
    port map (
            O => \N__44520\,
            I => \N__44455\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44519\,
            I => \N__44450\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44450\
        );

    \I__10103\ : Span4Mux_v
    port map (
            O => \N__44509\,
            I => \N__44441\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44506\,
            I => \N__44441\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__44501\,
            I => \N__44436\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44498\,
            I => \N__44436\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__44495\,
            I => \N__44430\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44490\,
            I => \N__44430\
        );

    \I__10097\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44423\
        );

    \I__10096\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44423\
        );

    \I__10095\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44423\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__44484\,
            I => \N__44406\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44406\
        );

    \I__10092\ : Sp12to4
    port map (
            O => \N__44478\,
            I => \N__44406\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__44473\,
            I => \N__44406\
        );

    \I__10090\ : Sp12to4
    port map (
            O => \N__44470\,
            I => \N__44406\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44465\,
            I => \N__44406\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__44462\,
            I => \N__44406\
        );

    \I__10087\ : Sp12to4
    port map (
            O => \N__44455\,
            I => \N__44406\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__44450\,
            I => \N__44403\
        );

    \I__10085\ : InMux
    port map (
            O => \N__44449\,
            I => \N__44394\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44448\,
            I => \N__44394\
        );

    \I__10083\ : InMux
    port map (
            O => \N__44447\,
            I => \N__44394\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44446\,
            I => \N__44394\
        );

    \I__10081\ : Span4Mux_h
    port map (
            O => \N__44441\,
            I => \N__44389\
        );

    \I__10080\ : Span4Mux_v
    port map (
            O => \N__44436\,
            I => \N__44389\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44386\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__44430\,
            I => \ALU.a_7\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44423\,
            I => \ALU.a_7\
        );

    \I__10076\ : Odrv12
    port map (
            O => \N__44406\,
            I => \ALU.a_7\
        );

    \I__10075\ : Odrv12
    port map (
            O => \N__44403\,
            I => \ALU.a_7\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__44394\,
            I => \ALU.a_7\
        );

    \I__10073\ : Odrv4
    port map (
            O => \N__44389\,
            I => \ALU.a_7\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__44386\,
            I => \ALU.a_7\
        );

    \I__10071\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44368\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__44368\,
            I => \ALU.r0_12_prm_6_7_s1_c_RNOZ0\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44365\,
            I => \N__44362\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44362\,
            I => \N__44356\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44361\,
            I => \N__44353\
        );

    \I__10066\ : InMux
    port map (
            O => \N__44360\,
            I => \N__44339\
        );

    \I__10065\ : InMux
    port map (
            O => \N__44359\,
            I => \N__44336\
        );

    \I__10064\ : Span4Mux_h
    port map (
            O => \N__44356\,
            I => \N__44332\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__44353\,
            I => \N__44329\
        );

    \I__10062\ : InMux
    port map (
            O => \N__44352\,
            I => \N__44322\
        );

    \I__10061\ : InMux
    port map (
            O => \N__44351\,
            I => \N__44322\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44350\,
            I => \N__44322\
        );

    \I__10059\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44319\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44314\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44347\,
            I => \N__44314\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44310\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44303\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44344\,
            I => \N__44303\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44343\,
            I => \N__44300\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44342\,
            I => \N__44297\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44339\,
            I => \N__44294\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__44336\,
            I => \N__44291\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44288\
        );

    \I__10048\ : Span4Mux_h
    port map (
            O => \N__44332\,
            I => \N__44283\
        );

    \I__10047\ : Span4Mux_h
    port map (
            O => \N__44329\,
            I => \N__44283\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44280\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__44319\,
            I => \N__44277\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44271\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44313\,
            I => \N__44268\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__44310\,
            I => \N__44265\
        );

    \I__10041\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44260\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44308\,
            I => \N__44260\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44253\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44300\,
            I => \N__44253\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__44297\,
            I => \N__44253\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__44294\,
            I => \N__44241\
        );

    \I__10035\ : Span4Mux_s3_v
    port map (
            O => \N__44291\,
            I => \N__44241\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44241\
        );

    \I__10033\ : Sp12to4
    port map (
            O => \N__44283\,
            I => \N__44234\
        );

    \I__10032\ : Span12Mux_h
    port map (
            O => \N__44280\,
            I => \N__44234\
        );

    \I__10031\ : Span12Mux_s5_h
    port map (
            O => \N__44277\,
            I => \N__44234\
        );

    \I__10030\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44227\
        );

    \I__10029\ : InMux
    port map (
            O => \N__44275\,
            I => \N__44227\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44274\,
            I => \N__44227\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__44271\,
            I => \N__44222\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__44268\,
            I => \N__44222\
        );

    \I__10025\ : Span12Mux_h
    port map (
            O => \N__44265\,
            I => \N__44215\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__44260\,
            I => \N__44215\
        );

    \I__10023\ : Span12Mux_s5_h
    port map (
            O => \N__44253\,
            I => \N__44215\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44210\
        );

    \I__10021\ : InMux
    port map (
            O => \N__44251\,
            I => \N__44210\
        );

    \I__10020\ : InMux
    port map (
            O => \N__44250\,
            I => \N__44203\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44249\,
            I => \N__44203\
        );

    \I__10018\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44203\
        );

    \I__10017\ : Odrv4
    port map (
            O => \N__44241\,
            I => \ALU.b_3\
        );

    \I__10016\ : Odrv12
    port map (
            O => \N__44234\,
            I => \ALU.b_3\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__44227\,
            I => \ALU.b_3\
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__44222\,
            I => \ALU.b_3\
        );

    \I__10013\ : Odrv12
    port map (
            O => \N__44215\,
            I => \ALU.b_3\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44210\,
            I => \ALU.b_3\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44203\,
            I => \ALU.b_3\
        );

    \I__10010\ : CascadeMux
    port map (
            O => \N__44188\,
            I => \N__44185\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44185\,
            I => \N__44182\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__44182\,
            I => \N__44179\
        );

    \I__10007\ : Span4Mux_h
    port map (
            O => \N__44179\,
            I => \N__44176\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__44176\,
            I => \ALU.r0_12_prm_1_5_s0_c_RNOZ0\
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__44173\,
            I => \N__44170\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44165\
        );

    \I__10003\ : InMux
    port map (
            O => \N__44169\,
            I => \N__44162\
        );

    \I__10002\ : CascadeMux
    port map (
            O => \N__44168\,
            I => \N__44159\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__44165\,
            I => \N__44155\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__44162\,
            I => \N__44152\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44149\
        );

    \I__9998\ : InMux
    port map (
            O => \N__44158\,
            I => \N__44146\
        );

    \I__9997\ : Span4Mux_h
    port map (
            O => \N__44155\,
            I => \N__44141\
        );

    \I__9996\ : Span4Mux_h
    port map (
            O => \N__44152\,
            I => \N__44141\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__44149\,
            I => \N__44136\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44146\,
            I => \N__44136\
        );

    \I__9993\ : Odrv4
    port map (
            O => \N__44141\,
            I => \ALU.rshift_7\
        );

    \I__9992\ : Odrv12
    port map (
            O => \N__44136\,
            I => \ALU.rshift_7\
        );

    \I__9991\ : InMux
    port map (
            O => \N__44131\,
            I => \N__44128\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__44128\,
            I => \ALU.r0_12_prm_8_7_s1_c_RNOZ0\
        );

    \I__9989\ : CascadeMux
    port map (
            O => \N__44125\,
            I => \N__44122\
        );

    \I__9988\ : InMux
    port map (
            O => \N__44122\,
            I => \N__44119\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__44119\,
            I => \N__44115\
        );

    \I__9986\ : CascadeMux
    port map (
            O => \N__44118\,
            I => \N__44112\
        );

    \I__9985\ : Span4Mux_h
    port map (
            O => \N__44115\,
            I => \N__44108\
        );

    \I__9984\ : InMux
    port map (
            O => \N__44112\,
            I => \N__44105\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44102\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__44108\,
            I => \ALU.lshift_7\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__44105\,
            I => \ALU.lshift_7\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__44102\,
            I => \ALU.lshift_7\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44095\,
            I => \N__44091\
        );

    \I__9978\ : CascadeMux
    port map (
            O => \N__44094\,
            I => \N__44088\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44085\
        );

    \I__9976\ : InMux
    port map (
            O => \N__44088\,
            I => \N__44082\
        );

    \I__9975\ : Span4Mux_v
    port map (
            O => \N__44085\,
            I => \N__44079\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44076\
        );

    \I__9973\ : Span4Mux_s1_v
    port map (
            O => \N__44079\,
            I => \N__44071\
        );

    \I__9972\ : Span4Mux_v
    port map (
            O => \N__44076\,
            I => \N__44071\
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__44071\,
            I => \ALU.un14_log_0_i_7\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44068\,
            I => \N__44065\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__44065\,
            I => \ALU.r0_12_prm_5_7_s1_c_RNOZ0\
        );

    \I__9968\ : CascadeMux
    port map (
            O => \N__44062\,
            I => \N__44059\
        );

    \I__9967\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44056\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__44056\,
            I => \N__44052\
        );

    \I__9965\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44049\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__44052\,
            I => \N__44046\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__44049\,
            I => \ALU.r4_RNIHENK8_0Z0Z_7\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__44046\,
            I => \ALU.r4_RNIHENK8_0Z0Z_7\
        );

    \I__9961\ : InMux
    port map (
            O => \N__44041\,
            I => \N__44038\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__44038\,
            I => \ALU.r0_12_prm_4_7_s1_c_RNOZ0\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__44035\,
            I => \N__44032\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44032\,
            I => \N__44029\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__44029\,
            I => \N__44025\
        );

    \I__9956\ : InMux
    port map (
            O => \N__44028\,
            I => \N__44022\
        );

    \I__9955\ : Span4Mux_h
    port map (
            O => \N__44025\,
            I => \N__44019\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__44022\,
            I => \ALU.a_i_7\
        );

    \I__9953\ : Odrv4
    port map (
            O => \N__44019\,
            I => \ALU.a_i_7\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44010\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44013\,
            I => \N__44005\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__44010\,
            I => \N__44002\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44009\,
            I => \N__43999\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44008\,
            I => \N__43996\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__44005\,
            I => \N__43993\
        );

    \I__9946\ : Span4Mux_h
    port map (
            O => \N__44002\,
            I => \N__43990\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__43999\,
            I => \N__43985\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__43996\,
            I => \N__43985\
        );

    \I__9943\ : Span4Mux_h
    port map (
            O => \N__43993\,
            I => \N__43982\
        );

    \I__9942\ : Sp12to4
    port map (
            O => \N__43990\,
            I => \N__43977\
        );

    \I__9941\ : Span12Mux_h
    port map (
            O => \N__43985\,
            I => \N__43977\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__43982\,
            I => \ALU.un2_addsub_cry_6_c_RNIPJK8EZ0\
        );

    \I__9939\ : Odrv12
    port map (
            O => \N__43977\,
            I => \ALU.un2_addsub_cry_6_c_RNIPJK8EZ0\
        );

    \I__9938\ : CascadeMux
    port map (
            O => \N__43972\,
            I => \N__43969\
        );

    \I__9937\ : InMux
    port map (
            O => \N__43969\,
            I => \N__43966\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__43966\,
            I => \ALU.r0_12_prm_2_7_s1_c_RNOZ0\
        );

    \I__9935\ : InMux
    port map (
            O => \N__43963\,
            I => \N__43958\
        );

    \I__9934\ : InMux
    port map (
            O => \N__43962\,
            I => \N__43955\
        );

    \I__9933\ : InMux
    port map (
            O => \N__43961\,
            I => \N__43951\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__43958\,
            I => \N__43944\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__43955\,
            I => \N__43941\
        );

    \I__9930\ : CascadeMux
    port map (
            O => \N__43954\,
            I => \N__43938\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__43951\,
            I => \N__43933\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43950\,
            I => \N__43921\
        );

    \I__9927\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43921\
        );

    \I__9926\ : InMux
    port map (
            O => \N__43948\,
            I => \N__43921\
        );

    \I__9925\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43917\
        );

    \I__9924\ : Span4Mux_v
    port map (
            O => \N__43944\,
            I => \N__43909\
        );

    \I__9923\ : Span4Mux_v
    port map (
            O => \N__43941\,
            I => \N__43909\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43938\,
            I => \N__43904\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43904\
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__43936\,
            I => \N__43901\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__43933\,
            I => \N__43893\
        );

    \I__9918\ : InMux
    port map (
            O => \N__43932\,
            I => \N__43888\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43888\
        );

    \I__9916\ : InMux
    port map (
            O => \N__43930\,
            I => \N__43883\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43880\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43928\,
            I => \N__43877\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__43921\,
            I => \N__43874\
        );

    \I__9912\ : InMux
    port map (
            O => \N__43920\,
            I => \N__43871\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__43917\,
            I => \N__43868\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43863\
        );

    \I__9909\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43863\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__43914\,
            I => \N__43857\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__43909\,
            I => \N__43854\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__43904\,
            I => \N__43851\
        );

    \I__9905\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43844\
        );

    \I__9904\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43844\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43844\
        );

    \I__9902\ : InMux
    port map (
            O => \N__43898\,
            I => \N__43841\
        );

    \I__9901\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43838\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43834\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__43893\,
            I => \N__43829\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43888\,
            I => \N__43829\
        );

    \I__9897\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43824\
        );

    \I__9896\ : InMux
    port map (
            O => \N__43886\,
            I => \N__43824\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__43883\,
            I => \N__43812\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__43880\,
            I => \N__43812\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__43877\,
            I => \N__43809\
        );

    \I__9892\ : Span4Mux_v
    port map (
            O => \N__43874\,
            I => \N__43804\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__43871\,
            I => \N__43804\
        );

    \I__9890\ : Span4Mux_v
    port map (
            O => \N__43868\,
            I => \N__43799\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__43863\,
            I => \N__43799\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43794\
        );

    \I__9887\ : InMux
    port map (
            O => \N__43861\,
            I => \N__43794\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43860\,
            I => \N__43789\
        );

    \I__9885\ : InMux
    port map (
            O => \N__43857\,
            I => \N__43789\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__43854\,
            I => \N__43782\
        );

    \I__9883\ : Span4Mux_s2_h
    port map (
            O => \N__43851\,
            I => \N__43782\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43844\,
            I => \N__43782\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43841\,
            I => \N__43777\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__43838\,
            I => \N__43777\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43774\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43767\
        );

    \I__9877\ : Span4Mux_h
    port map (
            O => \N__43829\,
            I => \N__43767\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__43824\,
            I => \N__43767\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43760\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43760\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43760\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43751\
        );

    \I__9871\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43751\
        );

    \I__9870\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43751\
        );

    \I__9869\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43751\
        );

    \I__9868\ : Span4Mux_s1_v
    port map (
            O => \N__43812\,
            I => \N__43744\
        );

    \I__9867\ : Span4Mux_h
    port map (
            O => \N__43809\,
            I => \N__43744\
        );

    \I__9866\ : Span4Mux_h
    port map (
            O => \N__43804\,
            I => \N__43744\
        );

    \I__9865\ : Odrv4
    port map (
            O => \N__43799\,
            I => \ALU.b_2\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__43794\,
            I => \ALU.b_2\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43789\,
            I => \ALU.b_2\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__43782\,
            I => \ALU.b_2\
        );

    \I__9861\ : Odrv12
    port map (
            O => \N__43777\,
            I => \ALU.b_2\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__43774\,
            I => \ALU.b_2\
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__43767\,
            I => \ALU.b_2\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__43760\,
            I => \ALU.b_2\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43751\,
            I => \ALU.b_2\
        );

    \I__9856\ : Odrv4
    port map (
            O => \N__43744\,
            I => \ALU.b_2\
        );

    \I__9855\ : CascadeMux
    port map (
            O => \N__43723\,
            I => \N__43720\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43720\,
            I => \N__43717\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__43717\,
            I => \N__43714\
        );

    \I__9852\ : Span4Mux_s0_v
    port map (
            O => \N__43714\,
            I => \N__43711\
        );

    \I__9851\ : Odrv4
    port map (
            O => \N__43711\,
            I => \ALU.r0_12_prm_5_2_c_RNOZ0Z_0\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43704\
        );

    \I__9849\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43701\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__43704\,
            I => \N__43698\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43701\,
            I => \N__43695\
        );

    \I__9846\ : Span4Mux_s3_v
    port map (
            O => \N__43698\,
            I => \N__43692\
        );

    \I__9845\ : Span4Mux_s3_v
    port map (
            O => \N__43695\,
            I => \N__43689\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__43692\,
            I => \N__43686\
        );

    \I__9843\ : Span4Mux_h
    port map (
            O => \N__43689\,
            I => \N__43683\
        );

    \I__9842\ : Odrv4
    port map (
            O => \N__43686\,
            I => \ALU.un9_addsub_cry_1_c_RNIKO6AJZ0\
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__43683\,
            I => \ALU.un9_addsub_cry_1_c_RNIKO6AJZ0\
        );

    \I__9840\ : CascadeMux
    port map (
            O => \N__43678\,
            I => \N__43675\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43675\,
            I => \N__43672\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43672\,
            I => \ALU.r0_12_prm_1_2_c_RNOZ0\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43669\,
            I => \N__43661\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43658\
        );

    \I__9835\ : CascadeMux
    port map (
            O => \N__43667\,
            I => \N__43652\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__43666\,
            I => \N__43645\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__43665\,
            I => \N__43640\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__43664\,
            I => \N__43632\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__43661\,
            I => \N__43628\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__43658\,
            I => \N__43625\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43657\,
            I => \N__43622\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43656\,
            I => \N__43619\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43655\,
            I => \N__43616\
        );

    \I__9826\ : InMux
    port map (
            O => \N__43652\,
            I => \N__43613\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43651\,
            I => \N__43608\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43650\,
            I => \N__43608\
        );

    \I__9823\ : CascadeMux
    port map (
            O => \N__43649\,
            I => \N__43603\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43600\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43597\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43594\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__43643\,
            I => \N__43591\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43640\,
            I => \N__43586\
        );

    \I__9817\ : InMux
    port map (
            O => \N__43639\,
            I => \N__43581\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43638\,
            I => \N__43581\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43637\,
            I => \N__43576\
        );

    \I__9814\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43576\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43635\,
            I => \N__43571\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43632\,
            I => \N__43571\
        );

    \I__9811\ : InMux
    port map (
            O => \N__43631\,
            I => \N__43567\
        );

    \I__9810\ : Span4Mux_s3_v
    port map (
            O => \N__43628\,
            I => \N__43562\
        );

    \I__9809\ : Span4Mux_v
    port map (
            O => \N__43625\,
            I => \N__43562\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__43622\,
            I => \N__43559\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43619\,
            I => \N__43554\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__43616\,
            I => \N__43554\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43551\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43608\,
            I => \N__43548\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43545\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43542\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43539\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__43600\,
            I => \N__43536\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43533\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43594\,
            I => \N__43530\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43527\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43590\,
            I => \N__43522\
        );

    \I__9795\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43522\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__43586\,
            I => \N__43517\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43581\,
            I => \N__43510\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__43576\,
            I => \N__43510\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__43571\,
            I => \N__43510\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43570\,
            I => \N__43507\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43567\,
            I => \N__43504\
        );

    \I__9788\ : Span4Mux_h
    port map (
            O => \N__43562\,
            I => \N__43495\
        );

    \I__9787\ : Span4Mux_s3_v
    port map (
            O => \N__43559\,
            I => \N__43495\
        );

    \I__9786\ : Span4Mux_s3_v
    port map (
            O => \N__43554\,
            I => \N__43495\
        );

    \I__9785\ : Span4Mux_v
    port map (
            O => \N__43551\,
            I => \N__43495\
        );

    \I__9784\ : Span4Mux_s2_h
    port map (
            O => \N__43548\,
            I => \N__43492\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43545\,
            I => \N__43487\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__43542\,
            I => \N__43487\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43539\,
            I => \N__43484\
        );

    \I__9780\ : Span4Mux_h
    port map (
            O => \N__43536\,
            I => \N__43473\
        );

    \I__9779\ : Span4Mux_h
    port map (
            O => \N__43533\,
            I => \N__43473\
        );

    \I__9778\ : Span4Mux_s0_v
    port map (
            O => \N__43530\,
            I => \N__43473\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__43527\,
            I => \N__43473\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43522\,
            I => \N__43473\
        );

    \I__9775\ : InMux
    port map (
            O => \N__43521\,
            I => \N__43468\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43468\
        );

    \I__9773\ : Span4Mux_h
    port map (
            O => \N__43517\,
            I => \N__43463\
        );

    \I__9772\ : Span4Mux_s3_h
    port map (
            O => \N__43510\,
            I => \N__43463\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__43507\,
            I => \N__43460\
        );

    \I__9770\ : Span4Mux_s2_h
    port map (
            O => \N__43504\,
            I => \N__43449\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__43495\,
            I => \N__43449\
        );

    \I__9768\ : Span4Mux_v
    port map (
            O => \N__43492\,
            I => \N__43449\
        );

    \I__9767\ : Span4Mux_s3_v
    port map (
            O => \N__43487\,
            I => \N__43449\
        );

    \I__9766\ : Span4Mux_s3_v
    port map (
            O => \N__43484\,
            I => \N__43449\
        );

    \I__9765\ : Odrv4
    port map (
            O => \N__43473\,
            I => \ALU.b_6\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__43468\,
            I => \ALU.b_6\
        );

    \I__9763\ : Odrv4
    port map (
            O => \N__43463\,
            I => \ALU.b_6\
        );

    \I__9762\ : Odrv4
    port map (
            O => \N__43460\,
            I => \ALU.b_6\
        );

    \I__9761\ : Odrv4
    port map (
            O => \N__43449\,
            I => \ALU.b_6\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43432\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__43437\,
            I => \N__43426\
        );

    \I__9758\ : InMux
    port map (
            O => \N__43436\,
            I => \N__43421\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43417\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43432\,
            I => \N__43412\
        );

    \I__9755\ : CascadeMux
    port map (
            O => \N__43431\,
            I => \N__43409\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43430\,
            I => \N__43405\
        );

    \I__9753\ : InMux
    port map (
            O => \N__43429\,
            I => \N__43400\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43426\,
            I => \N__43397\
        );

    \I__9751\ : CascadeMux
    port map (
            O => \N__43425\,
            I => \N__43390\
        );

    \I__9750\ : CascadeMux
    port map (
            O => \N__43424\,
            I => \N__43387\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43421\,
            I => \N__43384\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43420\,
            I => \N__43381\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43372\
        );

    \I__9746\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43369\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43366\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__43412\,
            I => \N__43362\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43359\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43356\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__43405\,
            I => \N__43352\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43404\,
            I => \N__43347\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43347\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__43400\,
            I => \N__43344\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43397\,
            I => \N__43341\
        );

    \I__9736\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43338\
        );

    \I__9735\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43333\
        );

    \I__9734\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43333\
        );

    \I__9733\ : InMux
    port map (
            O => \N__43393\,
            I => \N__43330\
        );

    \I__9732\ : InMux
    port map (
            O => \N__43390\,
            I => \N__43325\
        );

    \I__9731\ : InMux
    port map (
            O => \N__43387\,
            I => \N__43325\
        );

    \I__9730\ : Span4Mux_h
    port map (
            O => \N__43384\,
            I => \N__43320\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43320\
        );

    \I__9728\ : InMux
    port map (
            O => \N__43380\,
            I => \N__43315\
        );

    \I__9727\ : InMux
    port map (
            O => \N__43379\,
            I => \N__43315\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43378\,
            I => \N__43310\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43377\,
            I => \N__43310\
        );

    \I__9724\ : InMux
    port map (
            O => \N__43376\,
            I => \N__43303\
        );

    \I__9723\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43303\
        );

    \I__9722\ : Span4Mux_v
    port map (
            O => \N__43372\,
            I => \N__43300\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__43369\,
            I => \N__43297\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43366\,
            I => \N__43294\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43365\,
            I => \N__43291\
        );

    \I__9718\ : Span4Mux_h
    port map (
            O => \N__43362\,
            I => \N__43284\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43359\,
            I => \N__43284\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__43356\,
            I => \N__43284\
        );

    \I__9715\ : CascadeMux
    port map (
            O => \N__43355\,
            I => \N__43276\
        );

    \I__9714\ : Span4Mux_h
    port map (
            O => \N__43352\,
            I => \N__43269\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__43347\,
            I => \N__43269\
        );

    \I__9712\ : Span4Mux_s1_v
    port map (
            O => \N__43344\,
            I => \N__43269\
        );

    \I__9711\ : Span4Mux_h
    port map (
            O => \N__43341\,
            I => \N__43266\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__43338\,
            I => \N__43261\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43261\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43258\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__43325\,
            I => \N__43255\
        );

    \I__9706\ : Span4Mux_h
    port map (
            O => \N__43320\,
            I => \N__43252\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__43315\,
            I => \N__43247\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__43310\,
            I => \N__43247\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43242\
        );

    \I__9702\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43242\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__43303\,
            I => \N__43239\
        );

    \I__9700\ : Span4Mux_h
    port map (
            O => \N__43300\,
            I => \N__43228\
        );

    \I__9699\ : Span4Mux_s1_v
    port map (
            O => \N__43297\,
            I => \N__43228\
        );

    \I__9698\ : Span4Mux_v
    port map (
            O => \N__43294\,
            I => \N__43228\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__43291\,
            I => \N__43228\
        );

    \I__9696\ : Span4Mux_v
    port map (
            O => \N__43284\,
            I => \N__43228\
        );

    \I__9695\ : InMux
    port map (
            O => \N__43283\,
            I => \N__43221\
        );

    \I__9694\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43221\
        );

    \I__9693\ : InMux
    port map (
            O => \N__43281\,
            I => \N__43221\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43280\,
            I => \N__43218\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43279\,
            I => \N__43213\
        );

    \I__9690\ : InMux
    port map (
            O => \N__43276\,
            I => \N__43213\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__43269\,
            I => \N__43202\
        );

    \I__9688\ : Span4Mux_v
    port map (
            O => \N__43266\,
            I => \N__43202\
        );

    \I__9687\ : Span4Mux_v
    port map (
            O => \N__43261\,
            I => \N__43202\
        );

    \I__9686\ : Span4Mux_s3_h
    port map (
            O => \N__43258\,
            I => \N__43202\
        );

    \I__9685\ : Span4Mux_v
    port map (
            O => \N__43255\,
            I => \N__43202\
        );

    \I__9684\ : Span4Mux_h
    port map (
            O => \N__43252\,
            I => \N__43199\
        );

    \I__9683\ : Span12Mux_v
    port map (
            O => \N__43247\,
            I => \N__43194\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43242\,
            I => \N__43194\
        );

    \I__9681\ : Span4Mux_v
    port map (
            O => \N__43239\,
            I => \N__43189\
        );

    \I__9680\ : Span4Mux_h
    port map (
            O => \N__43228\,
            I => \N__43189\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__43221\,
            I => \ALU.a_6\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43218\,
            I => \ALU.a_6\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__43213\,
            I => \ALU.a_6\
        );

    \I__9676\ : Odrv4
    port map (
            O => \N__43202\,
            I => \ALU.a_6\
        );

    \I__9675\ : Odrv4
    port map (
            O => \N__43199\,
            I => \ALU.a_6\
        );

    \I__9674\ : Odrv12
    port map (
            O => \N__43194\,
            I => \ALU.a_6\
        );

    \I__9673\ : Odrv4
    port map (
            O => \N__43189\,
            I => \ALU.a_6\
        );

    \I__9672\ : CascadeMux
    port map (
            O => \N__43174\,
            I => \N__43171\
        );

    \I__9671\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43168\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43168\,
            I => \N__43165\
        );

    \I__9669\ : Span4Mux_h
    port map (
            O => \N__43165\,
            I => \N__43162\
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__43162\,
            I => \ALU.r0_12_prm_5_6_s0_c_RNOZ0\
        );

    \I__9667\ : CascadeMux
    port map (
            O => \N__43159\,
            I => \N__43156\
        );

    \I__9666\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43153\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43153\,
            I => \N__43150\
        );

    \I__9664\ : Span12Mux_v
    port map (
            O => \N__43150\,
            I => \N__43147\
        );

    \I__9663\ : Odrv12
    port map (
            O => \N__43147\,
            I => \ALU.r0_12_prm_5_7_s0_c_RNOZ0\
        );

    \I__9662\ : InMux
    port map (
            O => \N__43144\,
            I => \N__43141\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__43141\,
            I => \N__43135\
        );

    \I__9660\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43132\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43129\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43124\
        );

    \I__9657\ : Span4Mux_h
    port map (
            O => \N__43135\,
            I => \N__43118\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__43132\,
            I => \N__43118\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__43129\,
            I => \N__43115\
        );

    \I__9654\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43112\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43127\,
            I => \N__43109\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43124\,
            I => \N__43106\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43123\,
            I => \N__43103\
        );

    \I__9650\ : Span4Mux_v
    port map (
            O => \N__43118\,
            I => \N__43100\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__43115\,
            I => \N__43097\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__43112\,
            I => \N__43092\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__43109\,
            I => \N__43092\
        );

    \I__9646\ : Span12Mux_h
    port map (
            O => \N__43106\,
            I => \N__43089\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__43103\,
            I => \N__43086\
        );

    \I__9644\ : Span4Mux_v
    port map (
            O => \N__43100\,
            I => \N__43079\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__43097\,
            I => \N__43079\
        );

    \I__9642\ : Span4Mux_v
    port map (
            O => \N__43092\,
            I => \N__43079\
        );

    \I__9641\ : Span12Mux_v
    port map (
            O => \N__43089\,
            I => \N__43076\
        );

    \I__9640\ : Span12Mux_v
    port map (
            O => \N__43086\,
            I => \N__43071\
        );

    \I__9639\ : Sp12to4
    port map (
            O => \N__43079\,
            I => \N__43071\
        );

    \I__9638\ : Odrv12
    port map (
            O => \N__43076\,
            I => \ALU.r5_RNILM5AEZ0Z_15\
        );

    \I__9637\ : Odrv12
    port map (
            O => \N__43071\,
            I => \ALU.r5_RNILM5AEZ0Z_15\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43062\
        );

    \I__9635\ : InMux
    port map (
            O => \N__43065\,
            I => \N__43059\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__43056\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__43059\,
            I => \N__43049\
        );

    \I__9632\ : Span4Mux_v
    port map (
            O => \N__43056\,
            I => \N__43049\
        );

    \I__9631\ : InMux
    port map (
            O => \N__43055\,
            I => \N__43046\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43043\
        );

    \I__9629\ : Span4Mux_v
    port map (
            O => \N__43049\,
            I => \N__43038\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__43046\,
            I => \N__43038\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43043\,
            I => \ALU.r5_RNILV3HJZ0Z_12\
        );

    \I__9626\ : Odrv4
    port map (
            O => \N__43038\,
            I => \ALU.r5_RNILV3HJZ0Z_12\
        );

    \I__9625\ : InMux
    port map (
            O => \N__43033\,
            I => \N__43030\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__43030\,
            I => \N__43027\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__43027\,
            I => \N__43024\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__43024\,
            I => \N__43021\
        );

    \I__9621\ : Span4Mux_s2_v
    port map (
            O => \N__43021\,
            I => \N__43018\
        );

    \I__9620\ : Span4Mux_h
    port map (
            O => \N__43018\,
            I => \N__43015\
        );

    \I__9619\ : Odrv4
    port map (
            O => \N__43015\,
            I => \ALU.rshift_9\
        );

    \I__9618\ : InMux
    port map (
            O => \N__43012\,
            I => \N__43007\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43011\,
            I => \N__43004\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43010\,
            I => \N__43001\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__43007\,
            I => \N__42998\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__43004\,
            I => \N__42993\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43001\,
            I => \N__42993\
        );

    \I__9612\ : Odrv12
    port map (
            O => \N__42998\,
            I => \ALU.r4_RNI9H7SJZ0Z_5\
        );

    \I__9611\ : Odrv12
    port map (
            O => \N__42993\,
            I => \ALU.r4_RNI9H7SJZ0Z_5\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__42988\,
            I => \ALU.lshift_7_cascade_\
        );

    \I__9609\ : InMux
    port map (
            O => \N__42985\,
            I => \N__42982\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__42982\,
            I => \N__42979\
        );

    \I__9607\ : Span4Mux_h
    port map (
            O => \N__42979\,
            I => \N__42976\
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__42976\,
            I => \ALU.r0_12_prm_8_7_s0_c_RNOZ0\
        );

    \I__9605\ : InMux
    port map (
            O => \N__42973\,
            I => \ALU.r0_12_s1_9\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42970\,
            I => \N__42967\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__42967\,
            I => \N__42964\
        );

    \I__9602\ : Span4Mux_h
    port map (
            O => \N__42964\,
            I => \N__42961\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__42961\,
            I => \N__42958\
        );

    \I__9600\ : Odrv4
    port map (
            O => \N__42958\,
            I => \ALU.r0_12_s1_9_THRU_CO\
        );

    \I__9599\ : CascadeMux
    port map (
            O => \N__42955\,
            I => \N__42952\
        );

    \I__9598\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42949\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__42949\,
            I => \N__42946\
        );

    \I__9596\ : Span4Mux_v
    port map (
            O => \N__42946\,
            I => \N__42943\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__42943\,
            I => \N__42940\
        );

    \I__9594\ : Odrv4
    port map (
            O => \N__42940\,
            I => \ALU.r0_12_prm_7_14_s0_c_RNOZ0\
        );

    \I__9593\ : CascadeMux
    port map (
            O => \N__42937\,
            I => \N__42934\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42934\,
            I => \N__42931\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__42931\,
            I => \N__42928\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__42928\,
            I => \ALU.un14_log_0_i_2\
        );

    \I__9589\ : CascadeMux
    port map (
            O => \N__42925\,
            I => \N__42922\
        );

    \I__9588\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42919\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__42919\,
            I => \ALU.mult_2\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42916\,
            I => \N__42910\
        );

    \I__9585\ : InMux
    port map (
            O => \N__42915\,
            I => \N__42910\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__42910\,
            I => \N__42907\
        );

    \I__9583\ : Span4Mux_h
    port map (
            O => \N__42907\,
            I => \N__42904\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__42904\,
            I => \N__42901\
        );

    \I__9581\ : Odrv4
    port map (
            O => \N__42901\,
            I => \ALU.madd_cry_0_THRU_CO\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42898\,
            I => \N__42893\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42897\,
            I => \N__42888\
        );

    \I__9578\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42888\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__42893\,
            I => \N__42885\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__42888\,
            I => \N__42882\
        );

    \I__9575\ : Span4Mux_v
    port map (
            O => \N__42885\,
            I => \N__42879\
        );

    \I__9574\ : Odrv12
    port map (
            O => \N__42882\,
            I => \ALU.madd_axb_1\
        );

    \I__9573\ : Odrv4
    port map (
            O => \N__42879\,
            I => \ALU.madd_axb_1\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42871\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__42871\,
            I => \ALU.r0_12_prm_3_2_c_RNOZ0\
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__42868\,
            I => \N__42863\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42867\,
            I => \N__42858\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42866\,
            I => \N__42855\
        );

    \I__9567\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42852\
        );

    \I__9566\ : CascadeMux
    port map (
            O => \N__42862\,
            I => \N__42845\
        );

    \I__9565\ : InMux
    port map (
            O => \N__42861\,
            I => \N__42839\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__42858\,
            I => \N__42834\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__42855\,
            I => \N__42831\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__42852\,
            I => \N__42828\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42851\,
            I => \N__42822\
        );

    \I__9560\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42819\
        );

    \I__9559\ : InMux
    port map (
            O => \N__42849\,
            I => \N__42812\
        );

    \I__9558\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42809\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42804\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42804\
        );

    \I__9555\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42801\
        );

    \I__9554\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42798\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__42839\,
            I => \N__42795\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42792\
        );

    \I__9551\ : InMux
    port map (
            O => \N__42837\,
            I => \N__42789\
        );

    \I__9550\ : Span4Mux_v
    port map (
            O => \N__42834\,
            I => \N__42782\
        );

    \I__9549\ : Span4Mux_s2_v
    port map (
            O => \N__42831\,
            I => \N__42782\
        );

    \I__9548\ : Span4Mux_v
    port map (
            O => \N__42828\,
            I => \N__42779\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42827\,
            I => \N__42774\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42774\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42771\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42822\,
            I => \N__42766\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__42819\,
            I => \N__42766\
        );

    \I__9542\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42759\
        );

    \I__9541\ : InMux
    port map (
            O => \N__42817\,
            I => \N__42759\
        );

    \I__9540\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42759\
        );

    \I__9539\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42756\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__42812\,
            I => \N__42747\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42747\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__42804\,
            I => \N__42744\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__42801\,
            I => \N__42739\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__42798\,
            I => \N__42739\
        );

    \I__9533\ : Span4Mux_h
    port map (
            O => \N__42795\,
            I => \N__42734\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__42792\,
            I => \N__42734\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42789\,
            I => \N__42731\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42728\
        );

    \I__9529\ : CascadeMux
    port map (
            O => \N__42787\,
            I => \N__42720\
        );

    \I__9528\ : Span4Mux_h
    port map (
            O => \N__42782\,
            I => \N__42715\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__42779\,
            I => \N__42715\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__42774\,
            I => \N__42712\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__42771\,
            I => \N__42705\
        );

    \I__9524\ : Span4Mux_v
    port map (
            O => \N__42766\,
            I => \N__42705\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__42759\,
            I => \N__42705\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__42756\,
            I => \N__42702\
        );

    \I__9521\ : CascadeMux
    port map (
            O => \N__42755\,
            I => \N__42699\
        );

    \I__9520\ : CascadeMux
    port map (
            O => \N__42754\,
            I => \N__42696\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42691\
        );

    \I__9518\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42691\
        );

    \I__9517\ : Span4Mux_h
    port map (
            O => \N__42747\,
            I => \N__42686\
        );

    \I__9516\ : Span4Mux_v
    port map (
            O => \N__42744\,
            I => \N__42686\
        );

    \I__9515\ : Span4Mux_v
    port map (
            O => \N__42739\,
            I => \N__42683\
        );

    \I__9514\ : Span4Mux_v
    port map (
            O => \N__42734\,
            I => \N__42678\
        );

    \I__9513\ : Span4Mux_h
    port map (
            O => \N__42731\,
            I => \N__42678\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42728\,
            I => \N__42675\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42670\
        );

    \I__9510\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42670\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42663\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42663\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42663\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42720\,
            I => \N__42660\
        );

    \I__9505\ : Span4Mux_h
    port map (
            O => \N__42715\,
            I => \N__42655\
        );

    \I__9504\ : Span4Mux_s2_h
    port map (
            O => \N__42712\,
            I => \N__42655\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__42705\,
            I => \N__42650\
        );

    \I__9502\ : Span4Mux_s2_v
    port map (
            O => \N__42702\,
            I => \N__42650\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42699\,
            I => \N__42645\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42696\,
            I => \N__42645\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__42691\,
            I => \N__42642\
        );

    \I__9498\ : Span4Mux_h
    port map (
            O => \N__42686\,
            I => \N__42635\
        );

    \I__9497\ : Span4Mux_h
    port map (
            O => \N__42683\,
            I => \N__42635\
        );

    \I__9496\ : Span4Mux_h
    port map (
            O => \N__42678\,
            I => \N__42635\
        );

    \I__9495\ : Odrv4
    port map (
            O => \N__42675\,
            I => \ALU.a_4\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42670\,
            I => \ALU.a_4\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__42663\,
            I => \ALU.a_4\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__42660\,
            I => \ALU.a_4\
        );

    \I__9491\ : Odrv4
    port map (
            O => \N__42655\,
            I => \ALU.a_4\
        );

    \I__9490\ : Odrv4
    port map (
            O => \N__42650\,
            I => \ALU.a_4\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42645\,
            I => \ALU.a_4\
        );

    \I__9488\ : Odrv12
    port map (
            O => \N__42642\,
            I => \ALU.a_4\
        );

    \I__9487\ : Odrv4
    port map (
            O => \N__42635\,
            I => \ALU.a_4\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__42616\,
            I => \N__42613\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42610\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__42610\,
            I => \N__42607\
        );

    \I__9483\ : Span4Mux_v
    port map (
            O => \N__42607\,
            I => \N__42604\
        );

    \I__9482\ : Odrv4
    port map (
            O => \N__42604\,
            I => \ALU.r4_RNI87HO5Z0Z_4\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42598\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42595\
        );

    \I__9479\ : Span4Mux_h
    port map (
            O => \N__42595\,
            I => \N__42592\
        );

    \I__9478\ : Span4Mux_v
    port map (
            O => \N__42592\,
            I => \N__42589\
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__42589\,
            I => \ALU.r0_12_prm_8_9_s1_c_RNOZ0\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42586\,
            I => \N__42582\
        );

    \I__9475\ : CascadeMux
    port map (
            O => \N__42585\,
            I => \N__42579\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42582\,
            I => \N__42576\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42579\,
            I => \N__42573\
        );

    \I__9472\ : Span4Mux_v
    port map (
            O => \N__42576\,
            I => \N__42570\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42573\,
            I => \N__42567\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__42570\,
            I => \N__42562\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__42567\,
            I => \N__42562\
        );

    \I__9468\ : Span4Mux_v
    port map (
            O => \N__42562\,
            I => \N__42558\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42555\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__42558\,
            I => \ALU.lshift_9\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42555\,
            I => \ALU.lshift_9\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42547\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__42547\,
            I => \N__42544\
        );

    \I__9462\ : Odrv4
    port map (
            O => \N__42544\,
            I => \ALU.r0_12_prm_7_9_s1_c_RNOZ0\
        );

    \I__9461\ : InMux
    port map (
            O => \N__42541\,
            I => \N__42537\
        );

    \I__9460\ : CascadeMux
    port map (
            O => \N__42540\,
            I => \N__42534\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42537\,
            I => \N__42531\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42534\,
            I => \N__42528\
        );

    \I__9457\ : Span4Mux_h
    port map (
            O => \N__42531\,
            I => \N__42525\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42528\,
            I => \N__42522\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__42525\,
            I => \ALU.r4_RNISU5D9_0Z0Z_9\
        );

    \I__9454\ : Odrv4
    port map (
            O => \N__42522\,
            I => \ALU.r4_RNISU5D9_0Z0Z_9\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42514\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42514\,
            I => \N__42511\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__42511\,
            I => \ALU.r0_12_prm_6_9_s1_c_RNOZ0\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42504\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42501\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42504\,
            I => \N__42498\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42501\,
            I => \N__42495\
        );

    \I__9446\ : Span4Mux_h
    port map (
            O => \N__42498\,
            I => \N__42492\
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__42495\,
            I => \ALU.r4_RNISU5D9_1Z0Z_9\
        );

    \I__9444\ : Odrv4
    port map (
            O => \N__42492\,
            I => \ALU.r4_RNISU5D9_1Z0Z_9\
        );

    \I__9443\ : CascadeMux
    port map (
            O => \N__42487\,
            I => \N__42484\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42484\,
            I => \N__42481\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__42481\,
            I => \ALU.r0_12_prm_5_9_s1_c_RNOZ0\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__42478\,
            I => \N__42475\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42475\,
            I => \N__42472\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42472\,
            I => \N__42469\
        );

    \I__9437\ : Span4Mux_v
    port map (
            O => \N__42469\,
            I => \N__42465\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42462\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__42465\,
            I => \N__42459\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42462\,
            I => \ALU.a_i_9\
        );

    \I__9433\ : Odrv4
    port map (
            O => \N__42459\,
            I => \ALU.a_i_9\
        );

    \I__9432\ : InMux
    port map (
            O => \N__42454\,
            I => \N__42451\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__42451\,
            I => \ALU.r0_12_prm_2_9_s1_c_RNOZ0\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42448\,
            I => \N__42444\
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__42447\,
            I => \N__42441\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__42444\,
            I => \N__42437\
        );

    \I__9427\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42434\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42440\,
            I => \N__42431\
        );

    \I__9425\ : Span4Mux_h
    port map (
            O => \N__42437\,
            I => \N__42427\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__42434\,
            I => \N__42422\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__42431\,
            I => \N__42422\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42430\,
            I => \N__42419\
        );

    \I__9421\ : Span4Mux_h
    port map (
            O => \N__42427\,
            I => \N__42416\
        );

    \I__9420\ : Span4Mux_h
    port map (
            O => \N__42422\,
            I => \N__42413\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__42419\,
            I => \ALU.un2_addsub_cry_8_c_RNINO51FZ0\
        );

    \I__9418\ : Odrv4
    port map (
            O => \N__42416\,
            I => \ALU.un2_addsub_cry_8_c_RNINO51FZ0\
        );

    \I__9417\ : Odrv4
    port map (
            O => \N__42413\,
            I => \ALU.un2_addsub_cry_8_c_RNINO51FZ0\
        );

    \I__9416\ : InMux
    port map (
            O => \N__42406\,
            I => \N__42403\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__42403\,
            I => \ALU.r0_12_prm_1_9_s1_c_RNOZ0\
        );

    \I__9414\ : CascadeMux
    port map (
            O => \N__42400\,
            I => \N__42396\
        );

    \I__9413\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42392\
        );

    \I__9412\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42388\
        );

    \I__9411\ : InMux
    port map (
            O => \N__42395\,
            I => \N__42385\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__42392\,
            I => \N__42382\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42379\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42388\,
            I => \N__42374\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42385\,
            I => \N__42374\
        );

    \I__9406\ : Span4Mux_h
    port map (
            O => \N__42382\,
            I => \N__42369\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__42379\,
            I => \N__42369\
        );

    \I__9404\ : Span4Mux_v
    port map (
            O => \N__42374\,
            I => \N__42366\
        );

    \I__9403\ : Odrv4
    port map (
            O => \N__42369\,
            I => \ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9\
        );

    \I__9402\ : Odrv4
    port map (
            O => \N__42366\,
            I => \ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9\
        );

    \I__9401\ : InMux
    port map (
            O => \N__42361\,
            I => \N__42358\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__42358\,
            I => \N__42355\
        );

    \I__9399\ : Span4Mux_v
    port map (
            O => \N__42355\,
            I => \N__42352\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__42352\,
            I => \ALU.lshift_3_ns_1_10\
        );

    \I__9397\ : CascadeMux
    port map (
            O => \N__42349\,
            I => \ALU.r4_RNI67NNKZ0Z_7_cascade_\
        );

    \I__9396\ : CascadeMux
    port map (
            O => \N__42346\,
            I => \N__42343\
        );

    \I__9395\ : InMux
    port map (
            O => \N__42343\,
            I => \N__42339\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42342\,
            I => \N__42336\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__42339\,
            I => \N__42333\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__42336\,
            I => \N__42330\
        );

    \I__9391\ : Span4Mux_v
    port map (
            O => \N__42333\,
            I => \N__42327\
        );

    \I__9390\ : Odrv12
    port map (
            O => \N__42330\,
            I => \ALU.lshift_10\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__42327\,
            I => \ALU.lshift_10\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42322\,
            I => \N__42318\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42321\,
            I => \N__42313\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__42318\,
            I => \N__42310\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42305\
        );

    \I__9384\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42305\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42313\,
            I => \ALU.N_610_1\
        );

    \I__9382\ : Odrv12
    port map (
            O => \N__42310\,
            I => \ALU.N_610_1\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__42305\,
            I => \ALU.N_610_1\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42298\,
            I => \N__42295\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42295\,
            I => \N__42291\
        );

    \I__9378\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42288\
        );

    \I__9377\ : Odrv12
    port map (
            O => \N__42291\,
            I => \ALU.r4_RNIAHIIAZ0Z_2\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__42288\,
            I => \ALU.r4_RNIAHIIAZ0Z_2\
        );

    \I__9375\ : CascadeMux
    port map (
            O => \N__42283\,
            I => \N__42280\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42280\,
            I => \N__42274\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42279\,
            I => \N__42274\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__42274\,
            I => \ALU.r4_RNI38O1GZ0Z_2\
        );

    \I__9371\ : CascadeMux
    port map (
            O => \N__42271\,
            I => \ALU.r4_RNI38O1GZ0Z_2_cascade_\
        );

    \I__9370\ : InMux
    port map (
            O => \N__42268\,
            I => \N__42259\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42259\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42259\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42259\,
            I => \ALU.r4_RNICN8R81Z0Z_7\
        );

    \I__9366\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42253\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__42253\,
            I => \N__42250\
        );

    \I__9364\ : Span4Mux_v
    port map (
            O => \N__42250\,
            I => \N__42247\
        );

    \I__9363\ : Odrv4
    port map (
            O => \N__42247\,
            I => \ALU.r0_12_prm_8_10_s1_c_RNOZ0\
        );

    \I__9362\ : InMux
    port map (
            O => \N__42244\,
            I => \N__42241\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__42241\,
            I => \ALU.r4_RNI67NNKZ0Z_7\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42238\,
            I => \N__42235\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__42235\,
            I => \ALU.r5_RNI355TIZ0Z_13\
        );

    \I__9358\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42226\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42226\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__42226\,
            I => \N__42223\
        );

    \I__9355\ : Span4Mux_v
    port map (
            O => \N__42223\,
            I => \N__42219\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42216\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__42219\,
            I => \N__42213\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42216\,
            I => \ALU.r4_RNIO7CSJZ0Z_4\
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__42213\,
            I => \ALU.r4_RNIO7CSJZ0Z_4\
        );

    \I__9350\ : CascadeMux
    port map (
            O => \N__42208\,
            I => \ALU.lshift_15_ns_1_14_cascade_\
        );

    \I__9349\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42200\
        );

    \I__9348\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42194\
        );

    \I__9347\ : InMux
    port map (
            O => \N__42203\,
            I => \N__42194\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__42200\,
            I => \N__42191\
        );

    \I__9345\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42188\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__42194\,
            I => \N__42185\
        );

    \I__9343\ : Span4Mux_h
    port map (
            O => \N__42191\,
            I => \N__42182\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__42188\,
            I => \N__42179\
        );

    \I__9341\ : Odrv12
    port map (
            O => \N__42185\,
            I => \ALU.r4_RNILVIQFZ0Z_2\
        );

    \I__9340\ : Odrv4
    port map (
            O => \N__42182\,
            I => \ALU.r4_RNILVIQFZ0Z_2\
        );

    \I__9339\ : Odrv12
    port map (
            O => \N__42179\,
            I => \ALU.r4_RNILVIQFZ0Z_2\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42172\,
            I => \N__42169\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__42169\,
            I => \ALU.r0_12_prm_8_9_s1_c_RNOZ0Z_1\
        );

    \I__9336\ : InMux
    port map (
            O => \N__42166\,
            I => \ALU.r0_12_1\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42163\,
            I => \N__42160\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__42160\,
            I => \N__42157\
        );

    \I__9333\ : Span4Mux_v
    port map (
            O => \N__42157\,
            I => \N__42151\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42156\,
            I => \N__42148\
        );

    \I__9331\ : InMux
    port map (
            O => \N__42155\,
            I => \N__42144\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42154\,
            I => \N__42140\
        );

    \I__9329\ : Span4Mux_h
    port map (
            O => \N__42151\,
            I => \N__42136\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__42148\,
            I => \N__42133\
        );

    \I__9327\ : InMux
    port map (
            O => \N__42147\,
            I => \N__42130\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__42144\,
            I => \N__42126\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42123\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42140\,
            I => \N__42120\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42139\,
            I => \N__42117\
        );

    \I__9322\ : Span4Mux_v
    port map (
            O => \N__42136\,
            I => \N__42112\
        );

    \I__9321\ : Span4Mux_h
    port map (
            O => \N__42133\,
            I => \N__42112\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__42130\,
            I => \N__42109\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42106\
        );

    \I__9318\ : Span4Mux_h
    port map (
            O => \N__42126\,
            I => \N__42103\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__42123\,
            I => \N__42096\
        );

    \I__9316\ : Span4Mux_v
    port map (
            O => \N__42120\,
            I => \N__42096\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__42117\,
            I => \N__42096\
        );

    \I__9314\ : Span4Mux_h
    port map (
            O => \N__42112\,
            I => \N__42093\
        );

    \I__9313\ : Span4Mux_h
    port map (
            O => \N__42109\,
            I => \N__42090\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42106\,
            I => \N__42087\
        );

    \I__9311\ : Span4Mux_h
    port map (
            O => \N__42103\,
            I => \N__42082\
        );

    \I__9310\ : Span4Mux_v
    port map (
            O => \N__42096\,
            I => \N__42082\
        );

    \I__9309\ : Span4Mux_v
    port map (
            O => \N__42093\,
            I => \N__42079\
        );

    \I__9308\ : Span4Mux_h
    port map (
            O => \N__42090\,
            I => \N__42076\
        );

    \I__9307\ : Span12Mux_h
    port map (
            O => \N__42087\,
            I => \N__42073\
        );

    \I__9306\ : Span4Mux_h
    port map (
            O => \N__42082\,
            I => \N__42070\
        );

    \I__9305\ : Odrv4
    port map (
            O => \N__42079\,
            I => \ALU.r0_12_1_THRU_CO\
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__42076\,
            I => \ALU.r0_12_1_THRU_CO\
        );

    \I__9303\ : Odrv12
    port map (
            O => \N__42073\,
            I => \ALU.r0_12_1_THRU_CO\
        );

    \I__9302\ : Odrv4
    port map (
            O => \N__42070\,
            I => \ALU.r0_12_1_THRU_CO\
        );

    \I__9301\ : CascadeMux
    port map (
            O => \N__42061\,
            I => \N__42058\
        );

    \I__9300\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42052\
        );

    \I__9299\ : InMux
    port map (
            O => \N__42057\,
            I => \N__42052\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__42052\,
            I => \N__42049\
        );

    \I__9297\ : Span4Mux_v
    port map (
            O => \N__42049\,
            I => \N__42046\
        );

    \I__9296\ : Odrv4
    port map (
            O => \N__42046\,
            I => \ALU.un9_addsub_cry_0_c_RNIG8GLJZ0\
        );

    \I__9295\ : InMux
    port map (
            O => \N__42043\,
            I => \N__42040\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__42040\,
            I => \ALU.r0_12_prm_1_1_c_RNOZ0\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__42037\,
            I => \N__42034\
        );

    \I__9292\ : InMux
    port map (
            O => \N__42034\,
            I => \N__42031\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__42031\,
            I => \N__42028\
        );

    \I__9290\ : Odrv12
    port map (
            O => \N__42028\,
            I => \ALU.r0_12_prm_5_9_s0_c_RNOZ0\
        );

    \I__9289\ : CascadeMux
    port map (
            O => \N__42025\,
            I => \N__42022\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42022\,
            I => \N__42018\
        );

    \I__9287\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42015\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__42018\,
            I => \N__42012\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__42015\,
            I => \ALU.r4_RNIKUMQ8_0Z0Z_8\
        );

    \I__9284\ : Odrv12
    port map (
            O => \N__42012\,
            I => \ALU.r4_RNIKUMQ8_0Z0Z_8\
        );

    \I__9283\ : CascadeMux
    port map (
            O => \N__42007\,
            I => \N__42004\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42004\,
            I => \N__42001\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42001\,
            I => \ALU.r0_12_prm_6_8_s1_c_RNOZ0\
        );

    \I__9280\ : CascadeMux
    port map (
            O => \N__41998\,
            I => \N__41995\
        );

    \I__9279\ : InMux
    port map (
            O => \N__41995\,
            I => \N__41992\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41989\
        );

    \I__9277\ : Span12Mux_s9_h
    port map (
            O => \N__41989\,
            I => \N__41986\
        );

    \I__9276\ : Odrv12
    port map (
            O => \N__41986\,
            I => \ALU.r0_12_prm_8_10_s0_c_RNOZ0\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__41983\,
            I => \N__41980\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41980\,
            I => \N__41976\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41973\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41976\,
            I => \ALU.rshift_1\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41973\,
            I => \ALU.rshift_1\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__41968\,
            I => \N__41965\
        );

    \I__9269\ : InMux
    port map (
            O => \N__41965\,
            I => \N__41962\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__41962\,
            I => \N__41959\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__41959\,
            I => \ALU.lshift_1\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41956\,
            I => \N__41953\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__41953\,
            I => \N__41948\
        );

    \I__9264\ : InMux
    port map (
            O => \N__41952\,
            I => \N__41943\
        );

    \I__9263\ : InMux
    port map (
            O => \N__41951\,
            I => \N__41943\
        );

    \I__9262\ : Span4Mux_v
    port map (
            O => \N__41948\,
            I => \N__41939\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__41943\,
            I => \N__41936\
        );

    \I__9260\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41933\
        );

    \I__9259\ : Span4Mux_h
    port map (
            O => \N__41939\,
            I => \N__41928\
        );

    \I__9258\ : Span4Mux_h
    port map (
            O => \N__41936\,
            I => \N__41928\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__41933\,
            I => \ALU.a1_b_1\
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__41928\,
            I => \ALU.a1_b_1\
        );

    \I__9255\ : CascadeMux
    port map (
            O => \N__41923\,
            I => \N__41920\
        );

    \I__9254\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41917\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__41917\,
            I => \N__41914\
        );

    \I__9252\ : Span4Mux_h
    port map (
            O => \N__41914\,
            I => \N__41911\
        );

    \I__9251\ : Span4Mux_h
    port map (
            O => \N__41911\,
            I => \N__41908\
        );

    \I__9250\ : Odrv4
    port map (
            O => \N__41908\,
            I => \ALU.r0_12_prm_7_1_c_RNOZ0\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41905\,
            I => \N__41902\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__41902\,
            I => \N__41899\
        );

    \I__9247\ : Span4Mux_v
    port map (
            O => \N__41899\,
            I => \N__41896\
        );

    \I__9246\ : Odrv4
    port map (
            O => \N__41896\,
            I => \ALU.r0_12_prm_6_1_c_RNOZ0\
        );

    \I__9245\ : InMux
    port map (
            O => \N__41893\,
            I => \N__41890\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__41890\,
            I => \N__41887\
        );

    \I__9243\ : Span4Mux_h
    port map (
            O => \N__41887\,
            I => \N__41884\
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__41884\,
            I => \ALU.r0_12_prm_5_1_c_RNOZ0\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41881\,
            I => \N__41878\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41878\,
            I => \N__41875\
        );

    \I__9239\ : Span4Mux_v
    port map (
            O => \N__41875\,
            I => \N__41872\
        );

    \I__9238\ : Odrv4
    port map (
            O => \N__41872\,
            I => \ALU.r4_RNID1636Z0Z_1\
        );

    \I__9237\ : CascadeMux
    port map (
            O => \N__41869\,
            I => \N__41866\
        );

    \I__9236\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41863\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__41863\,
            I => \ALU.a_i_1\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41857\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__41857\,
            I => \N__41854\
        );

    \I__9232\ : Span4Mux_v
    port map (
            O => \N__41854\,
            I => \N__41851\
        );

    \I__9231\ : Sp12to4
    port map (
            O => \N__41851\,
            I => \N__41848\
        );

    \I__9230\ : Span12Mux_h
    port map (
            O => \N__41848\,
            I => \N__41845\
        );

    \I__9229\ : Odrv12
    port map (
            O => \N__41845\,
            I => \ALU.r0_12_prm_3_1_c_RNOZ0\
        );

    \I__9228\ : CascadeMux
    port map (
            O => \N__41842\,
            I => \N__41839\
        );

    \I__9227\ : InMux
    port map (
            O => \N__41839\,
            I => \N__41836\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41836\,
            I => \N__41833\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__41833\,
            I => \N__41830\
        );

    \I__9224\ : Span4Mux_h
    port map (
            O => \N__41830\,
            I => \N__41827\
        );

    \I__9223\ : Span4Mux_h
    port map (
            O => \N__41827\,
            I => \N__41824\
        );

    \I__9222\ : Span4Mux_h
    port map (
            O => \N__41824\,
            I => \N__41820\
        );

    \I__9221\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41817\
        );

    \I__9220\ : Span4Mux_s1_h
    port map (
            O => \N__41820\,
            I => \N__41812\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__41817\,
            I => \N__41812\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__41812\,
            I => \ALU.mult_1\
        );

    \I__9217\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41806\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__41806\,
            I => \ALU.r4_RNIVFRGQ_0Z0Z_2\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41803\,
            I => \N__41800\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__41800\,
            I => \ALU.r0_12_prm_8_4_c_RNOZ0\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41793\
        );

    \I__9212\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41790\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41787\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41790\,
            I => \N__41784\
        );

    \I__9209\ : Span4Mux_h
    port map (
            O => \N__41787\,
            I => \N__41781\
        );

    \I__9208\ : Span4Mux_v
    port map (
            O => \N__41784\,
            I => \N__41778\
        );

    \I__9207\ : Sp12to4
    port map (
            O => \N__41781\,
            I => \N__41775\
        );

    \I__9206\ : Odrv4
    port map (
            O => \N__41778\,
            I => \ALU.r4_RNIODO6KZ0Z_7\
        );

    \I__9205\ : Odrv12
    port map (
            O => \N__41775\,
            I => \ALU.r4_RNIODO6KZ0Z_7\
        );

    \I__9204\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41767\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__41767\,
            I => \N__41764\
        );

    \I__9202\ : Odrv4
    port map (
            O => \N__41764\,
            I => \ALU.r0_12_prm_8_4_c_RNOZ0Z_3\
        );

    \I__9201\ : InMux
    port map (
            O => \N__41761\,
            I => \N__41757\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41760\,
            I => \N__41754\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__41757\,
            I => \N__41751\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__41754\,
            I => \N__41748\
        );

    \I__9197\ : Span4Mux_h
    port map (
            O => \N__41751\,
            I => \N__41745\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__41748\,
            I => \N__41742\
        );

    \I__9195\ : Odrv4
    port map (
            O => \N__41745\,
            I => \ALU.un9_addsub_cry_3_c_RNIV8DFIZ0\
        );

    \I__9194\ : Odrv4
    port map (
            O => \N__41742\,
            I => \ALU.un9_addsub_cry_3_c_RNIV8DFIZ0\
        );

    \I__9193\ : CascadeMux
    port map (
            O => \N__41737\,
            I => \N__41734\
        );

    \I__9192\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41731\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__41731\,
            I => \ALU.r0_12_prm_1_4_c_RNOZ0\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41728\,
            I => \N__41723\
        );

    \I__9189\ : InMux
    port map (
            O => \N__41727\,
            I => \N__41718\
        );

    \I__9188\ : InMux
    port map (
            O => \N__41726\,
            I => \N__41718\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__41723\,
            I => \N__41715\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__41718\,
            I => \N__41712\
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__41715\,
            I => \ALU.r5_RNI7NOB9Z0Z_13\
        );

    \I__9184\ : Odrv12
    port map (
            O => \N__41712\,
            I => \ALU.r5_RNI7NOB9Z0Z_13\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41707\,
            I => \N__41703\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41700\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41703\,
            I => \N__41697\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41700\,
            I => \N__41694\
        );

    \I__9179\ : Span4Mux_s2_v
    port map (
            O => \N__41697\,
            I => \N__41691\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__41694\,
            I => \N__41688\
        );

    \I__9177\ : Span4Mux_h
    port map (
            O => \N__41691\,
            I => \N__41682\
        );

    \I__9176\ : Span4Mux_v
    port map (
            O => \N__41688\,
            I => \N__41679\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41687\,
            I => \N__41674\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41686\,
            I => \N__41674\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41685\,
            I => \N__41671\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__41682\,
            I => \ALU.r5_RNIUE7TIZ0Z_13\
        );

    \I__9171\ : Odrv4
    port map (
            O => \N__41679\,
            I => \ALU.r5_RNIUE7TIZ0Z_13\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41674\,
            I => \ALU.r5_RNIUE7TIZ0Z_13\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__41671\,
            I => \ALU.r5_RNIUE7TIZ0Z_13\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41658\
        );

    \I__9167\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41655\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41658\,
            I => \ALU.r4_RNIRL1V71Z0Z_7\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__41655\,
            I => \ALU.r4_RNIRL1V71Z0Z_7\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41650\,
            I => \N__41646\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41649\,
            I => \N__41643\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41646\,
            I => \N__41639\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41636\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41633\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__41639\,
            I => \N__41630\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__41636\,
            I => \N__41626\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41633\,
            I => \N__41623\
        );

    \I__9156\ : Span4Mux_h
    port map (
            O => \N__41630\,
            I => \N__41620\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41617\
        );

    \I__9154\ : Span4Mux_h
    port map (
            O => \N__41626\,
            I => \N__41614\
        );

    \I__9153\ : Span4Mux_h
    port map (
            O => \N__41623\,
            I => \N__41607\
        );

    \I__9152\ : Span4Mux_v
    port map (
            O => \N__41620\,
            I => \N__41607\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__41617\,
            I => \N__41607\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__41614\,
            I => \ALU.a6_b_6\
        );

    \I__9149\ : Odrv4
    port map (
            O => \N__41607\,
            I => \ALU.a6_b_6\
        );

    \I__9148\ : CascadeMux
    port map (
            O => \N__41602\,
            I => \N__41599\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41599\,
            I => \N__41596\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41596\,
            I => \N__41593\
        );

    \I__9145\ : Span4Mux_s2_v
    port map (
            O => \N__41593\,
            I => \N__41590\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__41590\,
            I => \ALU.r0_12_prm_7_6_s0_c_RNOZ0\
        );

    \I__9143\ : CascadeMux
    port map (
            O => \N__41587\,
            I => \N__41584\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41581\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__41581\,
            I => \N__41578\
        );

    \I__9140\ : Span12Mux_s4_v
    port map (
            O => \N__41578\,
            I => \N__41575\
        );

    \I__9139\ : Odrv12
    port map (
            O => \N__41575\,
            I => \ALU.r0_12_prm_6_6_s0_c_RNOZ0\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41567\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41571\,
            I => \N__41562\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41570\,
            I => \N__41558\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41567\,
            I => \N__41552\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41549\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__41565\,
            I => \N__41545\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__41562\,
            I => \N__41539\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41536\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41558\,
            I => \N__41533\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41557\,
            I => \N__41530\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41556\,
            I => \N__41527\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41555\,
            I => \N__41524\
        );

    \I__9126\ : Span4Mux_v
    port map (
            O => \N__41552\,
            I => \N__41521\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41549\,
            I => \N__41517\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41512\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41545\,
            I => \N__41512\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41544\,
            I => \N__41505\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41543\,
            I => \N__41505\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41505\
        );

    \I__9119\ : Span4Mux_h
    port map (
            O => \N__41539\,
            I => \N__41493\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__41536\,
            I => \N__41493\
        );

    \I__9117\ : Span4Mux_v
    port map (
            O => \N__41533\,
            I => \N__41490\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__41530\,
            I => \N__41485\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41527\,
            I => \N__41485\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41524\,
            I => \N__41482\
        );

    \I__9113\ : Span4Mux_v
    port map (
            O => \N__41521\,
            I => \N__41479\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41475\
        );

    \I__9111\ : Span4Mux_h
    port map (
            O => \N__41517\,
            I => \N__41472\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41512\,
            I => \N__41469\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__41505\,
            I => \N__41465\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41449\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41449\
        );

    \I__9106\ : InMux
    port map (
            O => \N__41502\,
            I => \N__41449\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41449\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41500\,
            I => \N__41449\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41449\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41449\
        );

    \I__9101\ : Span4Mux_v
    port map (
            O => \N__41493\,
            I => \N__41446\
        );

    \I__9100\ : Span4Mux_v
    port map (
            O => \N__41490\,
            I => \N__41442\
        );

    \I__9099\ : Span4Mux_v
    port map (
            O => \N__41485\,
            I => \N__41437\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__41482\,
            I => \N__41437\
        );

    \I__9097\ : Span4Mux_v
    port map (
            O => \N__41479\,
            I => \N__41434\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41478\,
            I => \N__41431\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41475\,
            I => \N__41428\
        );

    \I__9094\ : Span4Mux_v
    port map (
            O => \N__41472\,
            I => \N__41425\
        );

    \I__9093\ : Span4Mux_v
    port map (
            O => \N__41469\,
            I => \N__41422\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41419\
        );

    \I__9091\ : Span4Mux_v
    port map (
            O => \N__41465\,
            I => \N__41416\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41413\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41449\,
            I => \N__41408\
        );

    \I__9088\ : Span4Mux_h
    port map (
            O => \N__41446\,
            I => \N__41408\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41405\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__41442\,
            I => \N__41400\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__41437\,
            I => \N__41400\
        );

    \I__9084\ : Sp12to4
    port map (
            O => \N__41434\,
            I => \N__41395\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__41431\,
            I => \N__41395\
        );

    \I__9082\ : Span4Mux_h
    port map (
            O => \N__41428\,
            I => \N__41390\
        );

    \I__9081\ : Span4Mux_v
    port map (
            O => \N__41425\,
            I => \N__41390\
        );

    \I__9080\ : Span4Mux_v
    port map (
            O => \N__41422\,
            I => \N__41387\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__41419\,
            I => \ALU.a_13\
        );

    \I__9078\ : Odrv4
    port map (
            O => \N__41416\,
            I => \ALU.a_13\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__41413\,
            I => \ALU.a_13\
        );

    \I__9076\ : Odrv4
    port map (
            O => \N__41408\,
            I => \ALU.a_13\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41405\,
            I => \ALU.a_13\
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__41400\,
            I => \ALU.a_13\
        );

    \I__9073\ : Odrv12
    port map (
            O => \N__41395\,
            I => \ALU.a_13\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__41390\,
            I => \ALU.a_13\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__41387\,
            I => \ALU.a_13\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__41368\,
            I => \N__41359\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41367\,
            I => \N__41346\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41366\,
            I => \N__41343\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__41365\,
            I => \N__41340\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__41364\,
            I => \N__41336\
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__41363\,
            I => \N__41333\
        );

    \I__9064\ : CascadeMux
    port map (
            O => \N__41362\,
            I => \N__41330\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41324\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41324\
        );

    \I__9061\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41321\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41318\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41355\,
            I => \N__41311\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41354\,
            I => \N__41306\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41306\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41352\,
            I => \N__41303\
        );

    \I__9055\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41298\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41295\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41349\,
            I => \N__41290\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41346\,
            I => \N__41285\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41343\,
            I => \N__41285\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41282\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41277\
        );

    \I__9048\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41277\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41271\
        );

    \I__9046\ : InMux
    port map (
            O => \N__41330\,
            I => \N__41271\
        );

    \I__9045\ : InMux
    port map (
            O => \N__41329\,
            I => \N__41268\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__41324\,
            I => \N__41265\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41262\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__41318\,
            I => \N__41259\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41256\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41253\
        );

    \I__9039\ : InMux
    port map (
            O => \N__41315\,
            I => \N__41248\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41314\,
            I => \N__41248\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41311\,
            I => \N__41243\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__41306\,
            I => \N__41243\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__41303\,
            I => \N__41240\
        );

    \I__9034\ : InMux
    port map (
            O => \N__41302\,
            I => \N__41235\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41235\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__41298\,
            I => \N__41232\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41295\,
            I => \N__41229\
        );

    \I__9030\ : InMux
    port map (
            O => \N__41294\,
            I => \N__41224\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41224\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__41290\,
            I => \N__41221\
        );

    \I__9027\ : Span4Mux_v
    port map (
            O => \N__41285\,
            I => \N__41218\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41282\,
            I => \N__41213\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41277\,
            I => \N__41213\
        );

    \I__9024\ : InMux
    port map (
            O => \N__41276\,
            I => \N__41210\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__41271\,
            I => \N__41207\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__41268\,
            I => \N__41204\
        );

    \I__9021\ : Span4Mux_v
    port map (
            O => \N__41265\,
            I => \N__41199\
        );

    \I__9020\ : Span4Mux_h
    port map (
            O => \N__41262\,
            I => \N__41199\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__41259\,
            I => \N__41196\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__41256\,
            I => \N__41193\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41190\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__41248\,
            I => \N__41187\
        );

    \I__9015\ : Span4Mux_v
    port map (
            O => \N__41243\,
            I => \N__41180\
        );

    \I__9014\ : Span4Mux_v
    port map (
            O => \N__41240\,
            I => \N__41180\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41235\,
            I => \N__41180\
        );

    \I__9012\ : Span4Mux_h
    port map (
            O => \N__41232\,
            I => \N__41173\
        );

    \I__9011\ : Span4Mux_h
    port map (
            O => \N__41229\,
            I => \N__41173\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41173\
        );

    \I__9009\ : Span4Mux_v
    port map (
            O => \N__41221\,
            I => \N__41170\
        );

    \I__9008\ : Span4Mux_h
    port map (
            O => \N__41218\,
            I => \N__41167\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__41213\,
            I => \N__41162\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__41210\,
            I => \N__41162\
        );

    \I__9005\ : Span4Mux_h
    port map (
            O => \N__41207\,
            I => \N__41155\
        );

    \I__9004\ : Span4Mux_v
    port map (
            O => \N__41204\,
            I => \N__41155\
        );

    \I__9003\ : Span4Mux_h
    port map (
            O => \N__41199\,
            I => \N__41155\
        );

    \I__9002\ : Span4Mux_h
    port map (
            O => \N__41196\,
            I => \N__41150\
        );

    \I__9001\ : Span4Mux_h
    port map (
            O => \N__41193\,
            I => \N__41150\
        );

    \I__9000\ : Span4Mux_v
    port map (
            O => \N__41190\,
            I => \N__41145\
        );

    \I__8999\ : Span4Mux_v
    port map (
            O => \N__41187\,
            I => \N__41145\
        );

    \I__8998\ : Span4Mux_h
    port map (
            O => \N__41180\,
            I => \N__41140\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__41173\,
            I => \N__41140\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__41170\,
            I => \N__41135\
        );

    \I__8995\ : Span4Mux_h
    port map (
            O => \N__41167\,
            I => \N__41135\
        );

    \I__8994\ : Span4Mux_h
    port map (
            O => \N__41162\,
            I => \N__41132\
        );

    \I__8993\ : Odrv4
    port map (
            O => \N__41155\,
            I => \ALU.a_12\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__41150\,
            I => \ALU.a_12\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__41145\,
            I => \ALU.a_12\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__41140\,
            I => \ALU.a_12\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__41135\,
            I => \ALU.a_12\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__41132\,
            I => \ALU.a_12\
        );

    \I__8987\ : InMux
    port map (
            O => \N__41119\,
            I => \N__41115\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41112\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__41115\,
            I => \N__41109\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__41112\,
            I => \N__41104\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__41109\,
            I => \N__41104\
        );

    \I__8982\ : Span4Mux_v
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__8981\ : Odrv4
    port map (
            O => \N__41101\,
            I => \ALU.r4_RNI9H7SJZ0Z_6\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41098\,
            I => \N__41095\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__41095\,
            I => \N__41092\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__41092\,
            I => \N__41087\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41084\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41090\,
            I => \N__41081\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__41087\,
            I => \ALU.r5_RNI0QK3KZ0Z_11\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41084\,
            I => \ALU.r5_RNI0QK3KZ0Z_11\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__41081\,
            I => \ALU.r5_RNI0QK3KZ0Z_11\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__41074\,
            I => \ALU.r0_12_prm_8_4_c_RNOZ0Z_2_cascade_\
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__41071\,
            I => \N__41068\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41064\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41061\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__41064\,
            I => \ALU.rshift_4\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__41061\,
            I => \ALU.rshift_4\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41056\,
            I => \N__41053\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__41053\,
            I => \ALU.lshift_15_ns_1_8\
        );

    \I__8964\ : InMux
    port map (
            O => \N__41050\,
            I => \N__41047\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__41047\,
            I => \ALU.lshift_3_ns_1_4\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41044\,
            I => \N__41040\
        );

    \I__8961\ : InMux
    port map (
            O => \N__41043\,
            I => \N__41037\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__41040\,
            I => \ALU.r4_RNI6PL1LZ0Z_2\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__41037\,
            I => \ALU.r4_RNI6PL1LZ0Z_2\
        );

    \I__8958\ : CascadeMux
    port map (
            O => \N__41032\,
            I => \ALU.r4_RNI6PL1LZ0Z_2_cascade_\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41029\,
            I => \N__41026\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__41026\,
            I => \N__41021\
        );

    \I__8955\ : InMux
    port map (
            O => \N__41025\,
            I => \N__41018\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41024\,
            I => \N__41015\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__41021\,
            I => \N__41008\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41018\,
            I => \N__41008\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41008\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__41008\,
            I => \N__41005\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__41005\,
            I => \N__41002\
        );

    \I__8948\ : Odrv4
    port map (
            O => \N__41002\,
            I => \ALU.r4_RNIVFRGQZ0Z_2\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__40999\,
            I => \ALU.rshift_3_ns_1_9_cascade_\
        );

    \I__8946\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40993\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__40993\,
            I => \N__40983\
        );

    \I__8944\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40974\
        );

    \I__8943\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40974\
        );

    \I__8942\ : InMux
    port map (
            O => \N__40990\,
            I => \N__40974\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__40989\,
            I => \N__40971\
        );

    \I__8940\ : InMux
    port map (
            O => \N__40988\,
            I => \N__40951\
        );

    \I__8939\ : InMux
    port map (
            O => \N__40987\,
            I => \N__40951\
        );

    \I__8938\ : InMux
    port map (
            O => \N__40986\,
            I => \N__40948\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__40983\,
            I => \N__40945\
        );

    \I__8936\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40942\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40939\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40936\
        );

    \I__8933\ : InMux
    port map (
            O => \N__40971\,
            I => \N__40933\
        );

    \I__8932\ : CascadeMux
    port map (
            O => \N__40970\,
            I => \N__40928\
        );

    \I__8931\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40925\
        );

    \I__8930\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40912\
        );

    \I__8929\ : InMux
    port map (
            O => \N__40967\,
            I => \N__40912\
        );

    \I__8928\ : InMux
    port map (
            O => \N__40966\,
            I => \N__40912\
        );

    \I__8927\ : InMux
    port map (
            O => \N__40965\,
            I => \N__40912\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40964\,
            I => \N__40912\
        );

    \I__8925\ : InMux
    port map (
            O => \N__40963\,
            I => \N__40912\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40962\,
            I => \N__40908\
        );

    \I__8923\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40901\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40960\,
            I => \N__40901\
        );

    \I__8921\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40901\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40898\
        );

    \I__8919\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40893\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40893\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__40951\,
            I => \N__40889\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__40948\,
            I => \N__40886\
        );

    \I__8915\ : Span4Mux_v
    port map (
            O => \N__40945\,
            I => \N__40883\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__40942\,
            I => \N__40878\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40878\
        );

    \I__8912\ : Span4Mux_v
    port map (
            O => \N__40936\,
            I => \N__40871\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__40933\,
            I => \N__40871\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40932\,
            I => \N__40868\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40931\,
            I => \N__40865\
        );

    \I__8908\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40862\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__40925\,
            I => \N__40857\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__40912\,
            I => \N__40857\
        );

    \I__8905\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40854\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__40908\,
            I => \N__40851\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__40901\,
            I => \N__40846\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40898\,
            I => \N__40846\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__40893\,
            I => \N__40843\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40840\
        );

    \I__8899\ : Span4Mux_s1_h
    port map (
            O => \N__40889\,
            I => \N__40837\
        );

    \I__8898\ : Span4Mux_h
    port map (
            O => \N__40886\,
            I => \N__40834\
        );

    \I__8897\ : Span4Mux_h
    port map (
            O => \N__40883\,
            I => \N__40829\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__40878\,
            I => \N__40829\
        );

    \I__8895\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40824\
        );

    \I__8894\ : InMux
    port map (
            O => \N__40876\,
            I => \N__40824\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__40871\,
            I => \N__40817\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__40868\,
            I => \N__40817\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40865\,
            I => \N__40817\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__40862\,
            I => \N__40814\
        );

    \I__8889\ : Span4Mux_v
    port map (
            O => \N__40857\,
            I => \N__40811\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__40854\,
            I => \N__40806\
        );

    \I__8887\ : Span12Mux_v
    port map (
            O => \N__40851\,
            I => \N__40806\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__40846\,
            I => \N__40793\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__40843\,
            I => \N__40793\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__40840\,
            I => \N__40793\
        );

    \I__8883\ : Span4Mux_v
    port map (
            O => \N__40837\,
            I => \N__40793\
        );

    \I__8882\ : Span4Mux_v
    port map (
            O => \N__40834\,
            I => \N__40793\
        );

    \I__8881\ : Span4Mux_h
    port map (
            O => \N__40829\,
            I => \N__40793\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__40824\,
            I => \N__40788\
        );

    \I__8879\ : Span4Mux_h
    port map (
            O => \N__40817\,
            I => \N__40788\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__40814\,
            I => \N__40785\
        );

    \I__8877\ : Odrv4
    port map (
            O => \N__40811\,
            I => \ALU.a_11\
        );

    \I__8876\ : Odrv12
    port map (
            O => \N__40806\,
            I => \ALU.a_11\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__40793\,
            I => \ALU.a_11\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__40788\,
            I => \ALU.a_11\
        );

    \I__8873\ : Odrv4
    port map (
            O => \N__40785\,
            I => \ALU.a_11\
        );

    \I__8872\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40771\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__40771\,
            I => \N__40768\
        );

    \I__8870\ : Span12Mux_v
    port map (
            O => \N__40768\,
            I => \N__40765\
        );

    \I__8869\ : Odrv12
    port map (
            O => \N__40765\,
            I => \ALU.r0_12_prm_5_8_s0_c_RNOZ0\
        );

    \I__8868\ : CascadeMux
    port map (
            O => \N__40762\,
            I => \ALU.N_610_1_cascade_\
        );

    \I__8867\ : CascadeMux
    port map (
            O => \N__40759\,
            I => \ALU.r4_RNIVFRGQ_0Z0Z_2_cascade_\
        );

    \I__8866\ : CascadeMux
    port map (
            O => \N__40756\,
            I => \N__40753\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40750\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__40750\,
            I => \ALU.lshift_4\
        );

    \I__8863\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40743\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40740\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40737\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40740\,
            I => \N__40732\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__40737\,
            I => \N__40732\
        );

    \I__8858\ : Span4Mux_h
    port map (
            O => \N__40732\,
            I => \N__40727\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40731\,
            I => \N__40722\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40730\,
            I => \N__40722\
        );

    \I__8855\ : Span4Mux_h
    port map (
            O => \N__40727\,
            I => \N__40717\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40722\,
            I => \N__40717\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__40717\,
            I => \ALU.a2_b_2\
        );

    \I__8852\ : CascadeMux
    port map (
            O => \N__40714\,
            I => \N__40711\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40711\,
            I => \N__40708\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__40708\,
            I => \ALU.r0_12_prm_7_2_c_RNOZ0\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__40705\,
            I => \N__40701\
        );

    \I__8848\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40698\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40695\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__40698\,
            I => \N__40691\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40695\,
            I => \N__40688\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40694\,
            I => \N__40684\
        );

    \I__8843\ : Span4Mux_h
    port map (
            O => \N__40691\,
            I => \N__40679\
        );

    \I__8842\ : Span4Mux_s2_v
    port map (
            O => \N__40688\,
            I => \N__40679\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40676\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40684\,
            I => \N__40673\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__40679\,
            I => \ALU.lshift_0\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__40676\,
            I => \ALU.lshift_0\
        );

    \I__8837\ : Odrv4
    port map (
            O => \N__40673\,
            I => \ALU.lshift_0\
        );

    \I__8836\ : CascadeMux
    port map (
            O => \N__40666\,
            I => \N__40663\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40660\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__40660\,
            I => \N__40657\
        );

    \I__8833\ : Span4Mux_h
    port map (
            O => \N__40657\,
            I => \N__40654\
        );

    \I__8832\ : Span4Mux_v
    port map (
            O => \N__40654\,
            I => \N__40651\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__40651\,
            I => \ALU.r4_RNIHENK8_1Z0Z_7\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40648\,
            I => \N__40644\
        );

    \I__8829\ : CascadeMux
    port map (
            O => \N__40647\,
            I => \N__40641\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40644\,
            I => \N__40638\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40641\,
            I => \N__40635\
        );

    \I__8826\ : Span4Mux_v
    port map (
            O => \N__40638\,
            I => \N__40632\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__40635\,
            I => \N__40629\
        );

    \I__8824\ : Span4Mux_h
    port map (
            O => \N__40632\,
            I => \N__40624\
        );

    \I__8823\ : Span4Mux_h
    port map (
            O => \N__40629\,
            I => \N__40624\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__40624\,
            I => \N__40621\
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__40621\,
            I => \ALU.b_i_0\
        );

    \I__8820\ : CascadeMux
    port map (
            O => \N__40618\,
            I => \N__40614\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40611\
        );

    \I__8818\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40608\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__40611\,
            I => \N__40603\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__40608\,
            I => \N__40600\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40597\
        );

    \I__8814\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40594\
        );

    \I__8813\ : Span4Mux_s2_v
    port map (
            O => \N__40603\,
            I => \N__40587\
        );

    \I__8812\ : Span4Mux_s2_v
    port map (
            O => \N__40600\,
            I => \N__40587\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__40597\,
            I => \N__40587\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__40594\,
            I => \N__40584\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__40587\,
            I => \ALU.un2_addsub_axb_0_i\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__40584\,
            I => \ALU.un2_addsub_axb_0_i\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__40573\,
            I => \N__40569\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40572\,
            I => \N__40566\
        );

    \I__8803\ : Span4Mux_s1_v
    port map (
            O => \N__40569\,
            I => \N__40561\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40566\,
            I => \N__40561\
        );

    \I__8801\ : Span4Mux_v
    port map (
            O => \N__40561\,
            I => \N__40558\
        );

    \I__8800\ : Span4Mux_h
    port map (
            O => \N__40558\,
            I => \N__40555\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__40555\,
            I => \ALU.un2_addsub_cry_1_c_RNI1H7SGZ0\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40549\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40549\,
            I => \N__40546\
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__40546\,
            I => \ALU.r0_12_prm_2_2_c_RNOZ0\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40540\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40537\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__40537\,
            I => \ALU.r0_12_prm_6_2_c_RNOZ0\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40534\,
            I => \N__40527\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40524\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40532\,
            I => \N__40513\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40531\,
            I => \N__40513\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40530\,
            I => \N__40505\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__40527\,
            I => \N__40501\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40524\,
            I => \N__40498\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40495\
        );

    \I__8784\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40492\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40521\,
            I => \N__40489\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40482\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40477\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40477\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40513\,
            I => \N__40474\
        );

    \I__8778\ : InMux
    port map (
            O => \N__40512\,
            I => \N__40469\
        );

    \I__8777\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40469\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40510\,
            I => \N__40466\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40509\,
            I => \N__40461\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40508\,
            I => \N__40461\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__40505\,
            I => \N__40458\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40504\,
            I => \N__40455\
        );

    \I__8771\ : Span4Mux_h
    port map (
            O => \N__40501\,
            I => \N__40448\
        );

    \I__8770\ : Span4Mux_s2_v
    port map (
            O => \N__40498\,
            I => \N__40448\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40495\,
            I => \N__40448\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40492\,
            I => \N__40445\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40489\,
            I => \N__40442\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40488\,
            I => \N__40439\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40487\,
            I => \N__40434\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40434\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40425\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__40482\,
            I => \N__40420\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40477\,
            I => \N__40420\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__40474\,
            I => \N__40415\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40469\,
            I => \N__40415\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__40466\,
            I => \N__40410\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__40461\,
            I => \N__40410\
        );

    \I__8756\ : Span4Mux_s2_h
    port map (
            O => \N__40458\,
            I => \N__40407\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__40455\,
            I => \N__40404\
        );

    \I__8754\ : Span4Mux_h
    port map (
            O => \N__40448\,
            I => \N__40401\
        );

    \I__8753\ : Span12Mux_s4_v
    port map (
            O => \N__40445\,
            I => \N__40394\
        );

    \I__8752\ : Span12Mux_v
    port map (
            O => \N__40442\,
            I => \N__40394\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__40439\,
            I => \N__40394\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__40434\,
            I => \N__40391\
        );

    \I__8749\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40386\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40432\,
            I => \N__40386\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40431\,
            I => \N__40381\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40381\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40429\,
            I => \N__40376\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40428\,
            I => \N__40376\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40425\,
            I => \N__40371\
        );

    \I__8742\ : Span4Mux_h
    port map (
            O => \N__40420\,
            I => \N__40371\
        );

    \I__8741\ : Span4Mux_h
    port map (
            O => \N__40415\,
            I => \N__40366\
        );

    \I__8740\ : Span4Mux_v
    port map (
            O => \N__40410\,
            I => \N__40366\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__40407\,
            I => \N__40361\
        );

    \I__8738\ : Span4Mux_h
    port map (
            O => \N__40404\,
            I => \N__40361\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__40401\,
            I => \ALU.b_4\
        );

    \I__8736\ : Odrv12
    port map (
            O => \N__40394\,
            I => \ALU.b_4\
        );

    \I__8735\ : Odrv12
    port map (
            O => \N__40391\,
            I => \ALU.b_4\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40386\,
            I => \ALU.b_4\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40381\,
            I => \ALU.b_4\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40376\,
            I => \ALU.b_4\
        );

    \I__8731\ : Odrv4
    port map (
            O => \N__40371\,
            I => \ALU.b_4\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__40366\,
            I => \ALU.b_4\
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__40361\,
            I => \ALU.b_4\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40339\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40339\,
            I => \ALU.r0_12_prm_5_4_c_RNOZ0\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40336\,
            I => \N__40333\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40333\,
            I => \N__40330\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__40330\,
            I => \N__40327\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__40327\,
            I => \ALU.r0_12_prm_5_2_c_RNOZ0\
        );

    \I__8722\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40321\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40318\
        );

    \I__8720\ : Span4Mux_h
    port map (
            O => \N__40318\,
            I => \N__40315\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__40315\,
            I => \ALU.r4_RNIL9636Z0Z_2\
        );

    \I__8718\ : CascadeMux
    port map (
            O => \N__40312\,
            I => \N__40309\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40306\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__40306\,
            I => \ALU.a_i_2\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40303\,
            I => \ALU.r0_12_2\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40297\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__40297\,
            I => \N__40293\
        );

    \I__8712\ : InMux
    port map (
            O => \N__40296\,
            I => \N__40290\
        );

    \I__8711\ : Span4Mux_v
    port map (
            O => \N__40293\,
            I => \N__40282\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__40290\,
            I => \N__40282\
        );

    \I__8709\ : InMux
    port map (
            O => \N__40289\,
            I => \N__40279\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40276\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40287\,
            I => \N__40271\
        );

    \I__8706\ : Span4Mux_v
    port map (
            O => \N__40282\,
            I => \N__40268\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__40279\,
            I => \N__40263\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__40276\,
            I => \N__40263\
        );

    \I__8703\ : InMux
    port map (
            O => \N__40275\,
            I => \N__40260\
        );

    \I__8702\ : InMux
    port map (
            O => \N__40274\,
            I => \N__40257\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__40271\,
            I => \N__40254\
        );

    \I__8700\ : Span4Mux_h
    port map (
            O => \N__40268\,
            I => \N__40251\
        );

    \I__8699\ : Span4Mux_v
    port map (
            O => \N__40263\,
            I => \N__40244\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40260\,
            I => \N__40244\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__40257\,
            I => \N__40244\
        );

    \I__8696\ : Span4Mux_v
    port map (
            O => \N__40254\,
            I => \N__40240\
        );

    \I__8695\ : Span4Mux_h
    port map (
            O => \N__40251\,
            I => \N__40235\
        );

    \I__8694\ : Span4Mux_v
    port map (
            O => \N__40244\,
            I => \N__40235\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40232\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__40240\,
            I => \N__40229\
        );

    \I__8691\ : Span4Mux_h
    port map (
            O => \N__40235\,
            I => \N__40224\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__40232\,
            I => \N__40224\
        );

    \I__8689\ : Span4Mux_h
    port map (
            O => \N__40229\,
            I => \N__40221\
        );

    \I__8688\ : Span4Mux_v
    port map (
            O => \N__40224\,
            I => \N__40218\
        );

    \I__8687\ : Odrv4
    port map (
            O => \N__40221\,
            I => \ALU.r0_12_2_THRU_CO\
        );

    \I__8686\ : Odrv4
    port map (
            O => \N__40218\,
            I => \ALU.r0_12_2_THRU_CO\
        );

    \I__8685\ : CascadeMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__8684\ : InMux
    port map (
            O => \N__40210\,
            I => \N__40207\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__40207\,
            I => \ALU.lshift_2\
        );

    \I__8682\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40201\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__40201\,
            I => \ALU.r0_12_prm_8_2_c_RNOZ0\
        );

    \I__8680\ : CascadeMux
    port map (
            O => \N__40198\,
            I => \N__40195\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40195\,
            I => \N__40192\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40192\,
            I => \N__40189\
        );

    \I__8677\ : Span4Mux_h
    port map (
            O => \N__40189\,
            I => \N__40186\
        );

    \I__8676\ : Odrv4
    port map (
            O => \N__40186\,
            I => \ALU.r0_12_prm_8_0_s0_c_RNOZ0\
        );

    \I__8675\ : InMux
    port map (
            O => \N__40183\,
            I => \N__40177\
        );

    \I__8674\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40177\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__40177\,
            I => \N__40170\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40167\
        );

    \I__8671\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40164\
        );

    \I__8670\ : CascadeMux
    port map (
            O => \N__40174\,
            I => \N__40161\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40173\,
            I => \N__40151\
        );

    \I__8668\ : Span4Mux_h
    port map (
            O => \N__40170\,
            I => \N__40146\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__40167\,
            I => \N__40146\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40164\,
            I => \N__40143\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40135\
        );

    \I__8664\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40135\
        );

    \I__8663\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40135\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40158\,
            I => \N__40132\
        );

    \I__8661\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40129\
        );

    \I__8660\ : InMux
    port map (
            O => \N__40156\,
            I => \N__40126\
        );

    \I__8659\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40123\
        );

    \I__8658\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40120\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__40151\,
            I => \N__40115\
        );

    \I__8656\ : Span4Mux_v
    port map (
            O => \N__40146\,
            I => \N__40115\
        );

    \I__8655\ : Span4Mux_h
    port map (
            O => \N__40143\,
            I => \N__40110\
        );

    \I__8654\ : InMux
    port map (
            O => \N__40142\,
            I => \N__40107\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40103\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__40132\,
            I => \N__40098\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__40129\,
            I => \N__40098\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__40126\,
            I => \N__40092\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__40123\,
            I => \N__40092\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__40120\,
            I => \N__40087\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__40115\,
            I => \N__40087\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40081\
        );

    \I__8645\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40078\
        );

    \I__8644\ : Span4Mux_v
    port map (
            O => \N__40110\,
            I => \N__40075\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__40107\,
            I => \N__40072\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40106\,
            I => \N__40069\
        );

    \I__8641\ : Span4Mux_v
    port map (
            O => \N__40103\,
            I => \N__40066\
        );

    \I__8640\ : Span4Mux_v
    port map (
            O => \N__40098\,
            I => \N__40063\
        );

    \I__8639\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40060\
        );

    \I__8638\ : Span4Mux_v
    port map (
            O => \N__40092\,
            I => \N__40055\
        );

    \I__8637\ : Span4Mux_v
    port map (
            O => \N__40087\,
            I => \N__40055\
        );

    \I__8636\ : InMux
    port map (
            O => \N__40086\,
            I => \N__40049\
        );

    \I__8635\ : InMux
    port map (
            O => \N__40085\,
            I => \N__40049\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40084\,
            I => \N__40046\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__40081\,
            I => \N__40039\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__40078\,
            I => \N__40039\
        );

    \I__8631\ : Span4Mux_h
    port map (
            O => \N__40075\,
            I => \N__40039\
        );

    \I__8630\ : Span4Mux_h
    port map (
            O => \N__40072\,
            I => \N__40036\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40025\
        );

    \I__8628\ : Sp12to4
    port map (
            O => \N__40066\,
            I => \N__40025\
        );

    \I__8627\ : Sp12to4
    port map (
            O => \N__40063\,
            I => \N__40025\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__40060\,
            I => \N__40025\
        );

    \I__8625\ : Sp12to4
    port map (
            O => \N__40055\,
            I => \N__40025\
        );

    \I__8624\ : InMux
    port map (
            O => \N__40054\,
            I => \N__40022\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40049\,
            I => \ALU.a_15\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__40046\,
            I => \ALU.a_15\
        );

    \I__8621\ : Odrv4
    port map (
            O => \N__40039\,
            I => \ALU.a_15\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__40036\,
            I => \ALU.a_15\
        );

    \I__8619\ : Odrv12
    port map (
            O => \N__40025\,
            I => \ALU.a_15\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__40022\,
            I => \ALU.a_15\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40009\,
            I => \N__40004\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40008\,
            I => \N__40001\
        );

    \I__8615\ : InMux
    port map (
            O => \N__40007\,
            I => \N__39998\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__40004\,
            I => \N__39995\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__40001\,
            I => \N__39989\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__39998\,
            I => \N__39985\
        );

    \I__8611\ : Span4Mux_h
    port map (
            O => \N__39995\,
            I => \N__39982\
        );

    \I__8610\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39974\
        );

    \I__8609\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39974\
        );

    \I__8608\ : InMux
    port map (
            O => \N__39992\,
            I => \N__39974\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__39989\,
            I => \N__39970\
        );

    \I__8606\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39967\
        );

    \I__8605\ : Span4Mux_h
    port map (
            O => \N__39985\,
            I => \N__39964\
        );

    \I__8604\ : Span4Mux_v
    port map (
            O => \N__39982\,
            I => \N__39961\
        );

    \I__8603\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39958\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__39974\,
            I => \N__39954\
        );

    \I__8601\ : InMux
    port map (
            O => \N__39973\,
            I => \N__39951\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__39970\,
            I => \N__39946\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__39967\,
            I => \N__39946\
        );

    \I__8598\ : Span4Mux_h
    port map (
            O => \N__39964\,
            I => \N__39943\
        );

    \I__8597\ : Sp12to4
    port map (
            O => \N__39961\,
            I => \N__39938\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39958\,
            I => \N__39938\
        );

    \I__8595\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39935\
        );

    \I__8594\ : Span4Mux_h
    port map (
            O => \N__39954\,
            I => \N__39932\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__39951\,
            I => \N__39929\
        );

    \I__8592\ : Span4Mux_h
    port map (
            O => \N__39946\,
            I => \N__39926\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__39943\,
            I => \N__39922\
        );

    \I__8590\ : Span12Mux_h
    port map (
            O => \N__39938\,
            I => \N__39919\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39935\,
            I => \N__39910\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__39932\,
            I => \N__39910\
        );

    \I__8587\ : Span4Mux_s2_h
    port map (
            O => \N__39929\,
            I => \N__39910\
        );

    \I__8586\ : Span4Mux_h
    port map (
            O => \N__39926\,
            I => \N__39910\
        );

    \I__8585\ : InMux
    port map (
            O => \N__39925\,
            I => \N__39907\
        );

    \I__8584\ : Odrv4
    port map (
            O => \N__39922\,
            I => \ALU.b_15\
        );

    \I__8583\ : Odrv12
    port map (
            O => \N__39919\,
            I => \ALU.b_15\
        );

    \I__8582\ : Odrv4
    port map (
            O => \N__39910\,
            I => \ALU.b_15\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__39907\,
            I => \ALU.b_15\
        );

    \I__8580\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39895\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__39895\,
            I => \N__39892\
        );

    \I__8578\ : Odrv4
    port map (
            O => \N__39892\,
            I => \ALU.r0_12_prm_7_15_s0_c_RNOZ0\
        );

    \I__8577\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39886\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__39886\,
            I => \N__39883\
        );

    \I__8575\ : Span4Mux_h
    port map (
            O => \N__39883\,
            I => \N__39880\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__39880\,
            I => \ALU.r0_12_prm_8_13_s1_c_RNOZ0Z_1\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39877\,
            I => \N__39867\
        );

    \I__8572\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39867\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__39875\,
            I => \N__39864\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39854\
        );

    \I__8569\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39854\
        );

    \I__8568\ : InMux
    port map (
            O => \N__39872\,
            I => \N__39851\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__39867\,
            I => \N__39846\
        );

    \I__8566\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39843\
        );

    \I__8565\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39838\
        );

    \I__8564\ : InMux
    port map (
            O => \N__39862\,
            I => \N__39838\
        );

    \I__8563\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39834\
        );

    \I__8562\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39831\
        );

    \I__8561\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39827\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39854\,
            I => \N__39823\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__39851\,
            I => \N__39820\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__39850\,
            I => \N__39817\
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__39849\,
            I => \N__39814\
        );

    \I__8556\ : Span4Mux_v
    port map (
            O => \N__39846\,
            I => \N__39808\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39843\,
            I => \N__39808\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39805\
        );

    \I__8553\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39802\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__39834\,
            I => \N__39797\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__39831\,
            I => \N__39797\
        );

    \I__8550\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39794\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__39827\,
            I => \N__39791\
        );

    \I__8548\ : InMux
    port map (
            O => \N__39826\,
            I => \N__39788\
        );

    \I__8547\ : Span4Mux_v
    port map (
            O => \N__39823\,
            I => \N__39783\
        );

    \I__8546\ : Span4Mux_v
    port map (
            O => \N__39820\,
            I => \N__39783\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39780\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39814\,
            I => \N__39775\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39775\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__39808\,
            I => \N__39772\
        );

    \I__8541\ : Span4Mux_s2_h
    port map (
            O => \N__39805\,
            I => \N__39769\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__39802\,
            I => \N__39766\
        );

    \I__8539\ : Span4Mux_h
    port map (
            O => \N__39797\,
            I => \N__39763\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39758\
        );

    \I__8537\ : Span4Mux_v
    port map (
            O => \N__39791\,
            I => \N__39758\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__39788\,
            I => \N__39755\
        );

    \I__8535\ : Sp12to4
    port map (
            O => \N__39783\,
            I => \N__39752\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__39780\,
            I => \N__39747\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__39775\,
            I => \N__39747\
        );

    \I__8532\ : Span4Mux_h
    port map (
            O => \N__39772\,
            I => \N__39744\
        );

    \I__8531\ : Span4Mux_v
    port map (
            O => \N__39769\,
            I => \N__39739\
        );

    \I__8530\ : Span4Mux_s2_h
    port map (
            O => \N__39766\,
            I => \N__39739\
        );

    \I__8529\ : Span4Mux_h
    port map (
            O => \N__39763\,
            I => \N__39732\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__39758\,
            I => \N__39732\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__39755\,
            I => \N__39732\
        );

    \I__8526\ : Span12Mux_h
    port map (
            O => \N__39752\,
            I => \N__39727\
        );

    \I__8525\ : Sp12to4
    port map (
            O => \N__39747\,
            I => \N__39727\
        );

    \I__8524\ : Odrv4
    port map (
            O => \N__39744\,
            I => \ALU.b_12\
        );

    \I__8523\ : Odrv4
    port map (
            O => \N__39739\,
            I => \ALU.b_12\
        );

    \I__8522\ : Odrv4
    port map (
            O => \N__39732\,
            I => \ALU.b_12\
        );

    \I__8521\ : Odrv12
    port map (
            O => \N__39727\,
            I => \ALU.b_12\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__39718\,
            I => \N__39715\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39715\,
            I => \N__39712\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__39712\,
            I => \ALU.r0_12_prm_6_12_s1_c_RNOZ0\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39709\,
            I => \N__39706\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__39706\,
            I => \N__39703\
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__39703\,
            I => \ALU.r5_RNIPV8A9_0Z0Z_13\
        );

    \I__8514\ : CascadeMux
    port map (
            O => \N__39700\,
            I => \N__39697\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39697\,
            I => \N__39693\
        );

    \I__8512\ : InMux
    port map (
            O => \N__39696\,
            I => \N__39690\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__39693\,
            I => \ALU.rshift_2\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__39690\,
            I => \ALU.rshift_2\
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__39685\,
            I => \N__39682\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39682\,
            I => \N__39679\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39679\,
            I => \N__39676\
        );

    \I__8506\ : Span4Mux_h
    port map (
            O => \N__39676\,
            I => \N__39673\
        );

    \I__8505\ : Span4Mux_h
    port map (
            O => \N__39673\,
            I => \N__39670\
        );

    \I__8504\ : Odrv4
    port map (
            O => \N__39670\,
            I => \ALU.r5_RNITG1F5Z0Z_14\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39667\,
            I => \N__39664\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__39664\,
            I => \N__39661\
        );

    \I__8501\ : Odrv12
    port map (
            O => \N__39661\,
            I => \ALU.r0_12_prm_5_14_s0_c_RNOZ0\
        );

    \I__8500\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39655\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__39655\,
            I => \N__39652\
        );

    \I__8498\ : Span12Mux_v
    port map (
            O => \N__39652\,
            I => \N__39649\
        );

    \I__8497\ : Odrv12
    port map (
            O => \N__39649\,
            I => \ALU.rshift_13\
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__39646\,
            I => \N__39643\
        );

    \I__8495\ : InMux
    port map (
            O => \N__39643\,
            I => \N__39640\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__39640\,
            I => \N__39637\
        );

    \I__8493\ : Odrv12
    port map (
            O => \N__39637\,
            I => \ALU.r0_12_prm_6_14_s0_c_RNOZ0\
        );

    \I__8492\ : CascadeMux
    port map (
            O => \N__39634\,
            I => \N__39631\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39628\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__39628\,
            I => \N__39625\
        );

    \I__8489\ : Odrv12
    port map (
            O => \N__39625\,
            I => \ALU.r0_12_prm_8_14_s0_c_RNOZ0\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39622\,
            I => \N__39619\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39619\,
            I => \N__39613\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39618\,
            I => \N__39606\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39617\,
            I => \N__39606\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39616\,
            I => \N__39606\
        );

    \I__8483\ : Span4Mux_v
    port map (
            O => \N__39613\,
            I => \N__39603\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39606\,
            I => \N__39600\
        );

    \I__8481\ : Sp12to4
    port map (
            O => \N__39603\,
            I => \N__39597\
        );

    \I__8480\ : Span4Mux_v
    port map (
            O => \N__39600\,
            I => \N__39594\
        );

    \I__8479\ : Odrv12
    port map (
            O => \N__39597\,
            I => \ALU.un9_addsub_cry_7_c_RNINZ0Z3519\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__39594\,
            I => \ALU.un9_addsub_cry_7_c_RNINZ0Z3519\
        );

    \I__8477\ : CascadeMux
    port map (
            O => \N__39589\,
            I => \N__39586\
        );

    \I__8476\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39583\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__39583\,
            I => \ALU.r0_12_prm_1_8_s1_c_RNOZ0\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39580\,
            I => \N__39577\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__39577\,
            I => \N__39574\
        );

    \I__8472\ : Span4Mux_h
    port map (
            O => \N__39574\,
            I => \N__39571\
        );

    \I__8471\ : Span4Mux_h
    port map (
            O => \N__39571\,
            I => \N__39568\
        );

    \I__8470\ : Span4Mux_v
    port map (
            O => \N__39568\,
            I => \N__39565\
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__39565\,
            I => \ALU.madd_cry_6_THRU_CO\
        );

    \I__8468\ : InMux
    port map (
            O => \N__39562\,
            I => \N__39558\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39555\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__39558\,
            I => \N__39552\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39555\,
            I => \N__39549\
        );

    \I__8464\ : Span12Mux_v
    port map (
            O => \N__39552\,
            I => \N__39546\
        );

    \I__8463\ : Span4Mux_v
    port map (
            O => \N__39549\,
            I => \N__39543\
        );

    \I__8462\ : Odrv12
    port map (
            O => \N__39546\,
            I => \ALU.madd_axb_7\
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__39543\,
            I => \ALU.madd_axb_7\
        );

    \I__8460\ : CascadeMux
    port map (
            O => \N__39538\,
            I => \N__39535\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39532\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__39532\,
            I => \ALU.r0_12_s0_8_THRU_CO\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39529\,
            I => \ALU.r0_12_s1_8\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39520\
        );

    \I__8455\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39517\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39524\,
            I => \N__39514\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39510\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39520\,
            I => \N__39507\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39504\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__39514\,
            I => \N__39501\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39498\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39510\,
            I => \N__39495\
        );

    \I__8447\ : Span4Mux_h
    port map (
            O => \N__39507\,
            I => \N__39490\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__39504\,
            I => \N__39485\
        );

    \I__8445\ : Span4Mux_v
    port map (
            O => \N__39501\,
            I => \N__39485\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__39498\,
            I => \N__39482\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__39495\,
            I => \N__39479\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39494\,
            I => \N__39476\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39493\,
            I => \N__39473\
        );

    \I__8440\ : Span4Mux_h
    port map (
            O => \N__39490\,
            I => \N__39469\
        );

    \I__8439\ : Span4Mux_h
    port map (
            O => \N__39485\,
            I => \N__39466\
        );

    \I__8438\ : Span4Mux_h
    port map (
            O => \N__39482\,
            I => \N__39463\
        );

    \I__8437\ : Span4Mux_h
    port map (
            O => \N__39479\,
            I => \N__39458\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39476\,
            I => \N__39458\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__39473\,
            I => \N__39455\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39452\
        );

    \I__8433\ : Odrv4
    port map (
            O => \N__39469\,
            I => \ALU.r0_12_8\
        );

    \I__8432\ : Odrv4
    port map (
            O => \N__39466\,
            I => \ALU.r0_12_8\
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__39463\,
            I => \ALU.r0_12_8\
        );

    \I__8430\ : Odrv4
    port map (
            O => \N__39458\,
            I => \ALU.r0_12_8\
        );

    \I__8429\ : Odrv12
    port map (
            O => \N__39455\,
            I => \ALU.r0_12_8\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39452\,
            I => \ALU.r0_12_8\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39439\,
            I => \N__39435\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39438\,
            I => \N__39432\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39435\,
            I => \N__39428\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39432\,
            I => \N__39425\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39431\,
            I => \N__39422\
        );

    \I__8422\ : Span4Mux_h
    port map (
            O => \N__39428\,
            I => \N__39419\
        );

    \I__8421\ : Span4Mux_h
    port map (
            O => \N__39425\,
            I => \N__39414\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__39422\,
            I => \N__39414\
        );

    \I__8419\ : Span4Mux_h
    port map (
            O => \N__39419\,
            I => \N__39411\
        );

    \I__8418\ : Span4Mux_h
    port map (
            O => \N__39414\,
            I => \N__39408\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__39411\,
            I => r0_8
        );

    \I__8416\ : Odrv4
    port map (
            O => \N__39408\,
            I => r0_8
        );

    \I__8415\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39398\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39395\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39392\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39398\,
            I => \N__39388\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__39395\,
            I => \N__39383\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__39392\,
            I => \N__39383\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39380\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__39388\,
            I => \N__39377\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__39383\,
            I => \ALU.un2_addsub_cry_7_c_RNI5ELEEZ0\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39380\,
            I => \ALU.un2_addsub_cry_7_c_RNI5ELEEZ0\
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__39377\,
            I => \ALU.un2_addsub_cry_7_c_RNI5ELEEZ0\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__39370\,
            I => \N__39367\
        );

    \I__8403\ : InMux
    port map (
            O => \N__39367\,
            I => \N__39364\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__39364\,
            I => \N__39361\
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__39361\,
            I => \ALU.r0_12_prm_2_8_s0_c_RNOZ0\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39358\,
            I => \N__39355\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__39355\,
            I => \N__39352\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__39352\,
            I => \ALU.r5_RNITTMB9Z0Z_12\
        );

    \I__8397\ : CascadeMux
    port map (
            O => \N__39349\,
            I => \ALU.r5_RNITTMB9Z0Z_12_cascade_\
        );

    \I__8396\ : CascadeMux
    port map (
            O => \N__39346\,
            I => \ALU.rshift_15_ns_1_1_cascade_\
        );

    \I__8395\ : CascadeMux
    port map (
            O => \N__39343\,
            I => \N__39340\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39337\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__39337\,
            I => \N__39334\
        );

    \I__8392\ : Odrv12
    port map (
            O => \N__39334\,
            I => \ALU.r0_12_prm_8_8_s1_c_RNOZ0Z_1\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__39331\,
            I => \N__39328\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39328\,
            I => \N__39324\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39321\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__39324\,
            I => \N__39318\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39321\,
            I => \N__39312\
        );

    \I__8386\ : Span4Mux_h
    port map (
            O => \N__39318\,
            I => \N__39312\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39309\
        );

    \I__8384\ : Odrv4
    port map (
            O => \N__39312\,
            I => \ALU.lshift_8\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__39309\,
            I => \ALU.lshift_8\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__39304\,
            I => \N__39301\
        );

    \I__8381\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39298\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__39298\,
            I => \N__39295\
        );

    \I__8379\ : Odrv12
    port map (
            O => \N__39295\,
            I => \ALU.r0_12_prm_8_8_s1_c_RNOZ0\
        );

    \I__8378\ : CascadeMux
    port map (
            O => \N__39292\,
            I => \N__39288\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39285\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39282\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__39285\,
            I => \N__39277\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__39282\,
            I => \N__39277\
        );

    \I__8373\ : Span4Mux_v
    port map (
            O => \N__39277\,
            I => \N__39274\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__39274\,
            I => \N__39271\
        );

    \I__8371\ : Sp12to4
    port map (
            O => \N__39271\,
            I => \N__39268\
        );

    \I__8370\ : Odrv12
    port map (
            O => \N__39268\,
            I => \ALU.a8_b_8\
        );

    \I__8369\ : InMux
    port map (
            O => \N__39265\,
            I => \N__39261\
        );

    \I__8368\ : CascadeMux
    port map (
            O => \N__39264\,
            I => \N__39258\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__39261\,
            I => \N__39255\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39258\,
            I => \N__39252\
        );

    \I__8365\ : Span4Mux_h
    port map (
            O => \N__39255\,
            I => \N__39247\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__39252\,
            I => \N__39247\
        );

    \I__8363\ : Span4Mux_v
    port map (
            O => \N__39247\,
            I => \N__39244\
        );

    \I__8362\ : Odrv4
    port map (
            O => \N__39244\,
            I => \ALU.un14_log_0_i_8\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39238\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39238\,
            I => \ALU.r0_12_prm_4_8_s1_c_RNOZ0\
        );

    \I__8359\ : CascadeMux
    port map (
            O => \N__39235\,
            I => \N__39231\
        );

    \I__8358\ : CascadeMux
    port map (
            O => \N__39234\,
            I => \N__39228\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39231\,
            I => \N__39225\
        );

    \I__8356\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39222\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39225\,
            I => \ALU.a_i_8\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__39222\,
            I => \ALU.a_i_8\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__39217\,
            I => \N__39214\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39211\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39211\,
            I => \N__39208\
        );

    \I__8350\ : Odrv4
    port map (
            O => \N__39208\,
            I => \ALU.r0_12_prm_2_8_s1_c_RNOZ0\
        );

    \I__8349\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39202\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__39202\,
            I => \N__39197\
        );

    \I__8347\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39192\
        );

    \I__8346\ : InMux
    port map (
            O => \N__39200\,
            I => \N__39192\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__39197\,
            I => \N__39189\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__39192\,
            I => \N__39186\
        );

    \I__8343\ : Sp12to4
    port map (
            O => \N__39189\,
            I => \N__39183\
        );

    \I__8342\ : Span4Mux_h
    port map (
            O => \N__39186\,
            I => \N__39180\
        );

    \I__8341\ : Span12Mux_v
    port map (
            O => \N__39183\,
            I => \N__39177\
        );

    \I__8340\ : Span4Mux_h
    port map (
            O => \N__39180\,
            I => \N__39174\
        );

    \I__8339\ : Odrv12
    port map (
            O => \N__39177\,
            I => r6_8
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__39174\,
            I => r6_8
        );

    \I__8337\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39164\
        );

    \I__8336\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39159\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39159\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__39164\,
            I => \N__39156\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__39159\,
            I => \N__39153\
        );

    \I__8332\ : Span4Mux_h
    port map (
            O => \N__39156\,
            I => \N__39150\
        );

    \I__8331\ : Span12Mux_s5_h
    port map (
            O => \N__39153\,
            I => \N__39147\
        );

    \I__8330\ : Span4Mux_h
    port map (
            O => \N__39150\,
            I => \N__39144\
        );

    \I__8329\ : Odrv12
    port map (
            O => \N__39147\,
            I => r6_2
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__39144\,
            I => r6_2
        );

    \I__8327\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39136\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__39136\,
            I => \N__39133\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__39133\,
            I => \N__39129\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39125\
        );

    \I__8323\ : Span4Mux_h
    port map (
            O => \N__39129\,
            I => \N__39122\
        );

    \I__8322\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39119\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__39125\,
            I => \N__39116\
        );

    \I__8320\ : Span4Mux_h
    port map (
            O => \N__39122\,
            I => \N__39113\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39119\,
            I => \N__39110\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__39116\,
            I => \N__39107\
        );

    \I__8317\ : Span4Mux_h
    port map (
            O => \N__39113\,
            I => \N__39104\
        );

    \I__8316\ : Span12Mux_v
    port map (
            O => \N__39110\,
            I => \N__39101\
        );

    \I__8315\ : Span4Mux_h
    port map (
            O => \N__39107\,
            I => \N__39098\
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__39104\,
            I => r6_3
        );

    \I__8313\ : Odrv12
    port map (
            O => \N__39101\,
            I => r6_3
        );

    \I__8312\ : Odrv4
    port map (
            O => \N__39098\,
            I => r6_3
        );

    \I__8311\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39087\
        );

    \I__8310\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39084\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__39087\,
            I => \N__39079\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__39084\,
            I => \N__39075\
        );

    \I__8307\ : InMux
    port map (
            O => \N__39083\,
            I => \N__39072\
        );

    \I__8306\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39069\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__39079\,
            I => \N__39066\
        );

    \I__8304\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39063\
        );

    \I__8303\ : Span4Mux_v
    port map (
            O => \N__39075\,
            I => \N__39059\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__39072\,
            I => \N__39056\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__39069\,
            I => \N__39053\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__39066\,
            I => \N__39047\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__39063\,
            I => \N__39047\
        );

    \I__8298\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39044\
        );

    \I__8297\ : Span4Mux_h
    port map (
            O => \N__39059\,
            I => \N__39038\
        );

    \I__8296\ : Span4Mux_h
    port map (
            O => \N__39056\,
            I => \N__39038\
        );

    \I__8295\ : Span4Mux_h
    port map (
            O => \N__39053\,
            I => \N__39035\
        );

    \I__8294\ : InMux
    port map (
            O => \N__39052\,
            I => \N__39032\
        );

    \I__8293\ : Span4Mux_v
    port map (
            O => \N__39047\,
            I => \N__39027\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__39044\,
            I => \N__39027\
        );

    \I__8291\ : InMux
    port map (
            O => \N__39043\,
            I => \N__39024\
        );

    \I__8290\ : Span4Mux_v
    port map (
            O => \N__39038\,
            I => \N__39021\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__39035\,
            I => \N__39018\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__39032\,
            I => \N__39015\
        );

    \I__8287\ : Span4Mux_h
    port map (
            O => \N__39027\,
            I => \N__39010\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__39024\,
            I => \N__39010\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__39021\,
            I => \ALU.r0_12_4_THRU_CO\
        );

    \I__8284\ : Odrv4
    port map (
            O => \N__39018\,
            I => \ALU.r0_12_4_THRU_CO\
        );

    \I__8283\ : Odrv12
    port map (
            O => \N__39015\,
            I => \ALU.r0_12_4_THRU_CO\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__39010\,
            I => \ALU.r0_12_4_THRU_CO\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38992\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39000\,
            I => \N__38992\
        );

    \I__8279\ : InMux
    port map (
            O => \N__38999\,
            I => \N__38992\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__38992\,
            I => \N__38989\
        );

    \I__8277\ : Span4Mux_h
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__8276\ : Span4Mux_h
    port map (
            O => \N__38986\,
            I => \N__38983\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__38983\,
            I => r6_4
        );

    \I__8274\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38977\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__38977\,
            I => \ALU.r4_RNIN3236Z0Z_8\
        );

    \I__8272\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38971\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__38971\,
            I => \N__38968\
        );

    \I__8270\ : Span4Mux_v
    port map (
            O => \N__38968\,
            I => \N__38965\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__38965\,
            I => \N__38962\
        );

    \I__8268\ : Span4Mux_h
    port map (
            O => \N__38962\,
            I => \N__38959\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__38959\,
            I => \ALU.rshift_3_ns_1_1\
        );

    \I__8266\ : CascadeMux
    port map (
            O => \N__38956\,
            I => \ALU.r0_12_prm_8_1_c_RNOZ0Z_3_cascade_\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__38953\,
            I => \N__38950\
        );

    \I__8264\ : InMux
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38947\,
            I => \ALU.r0_12_prm_2_7_s0_c_RNOZ0\
        );

    \I__8262\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38940\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38943\,
            I => \N__38937\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38940\,
            I => \N__38934\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__38937\,
            I => \N__38931\
        );

    \I__8258\ : Span4Mux_h
    port map (
            O => \N__38934\,
            I => \N__38928\
        );

    \I__8257\ : Span12Mux_v
    port map (
            O => \N__38931\,
            I => \N__38925\
        );

    \I__8256\ : Odrv4
    port map (
            O => \N__38928\,
            I => \ALU.r4_RNIODO6KZ0Z_5\
        );

    \I__8255\ : Odrv12
    port map (
            O => \N__38925\,
            I => \ALU.r4_RNIODO6KZ0Z_5\
        );

    \I__8254\ : CascadeMux
    port map (
            O => \N__38920\,
            I => \ALU.lshift_8_cascade_\
        );

    \I__8253\ : InMux
    port map (
            O => \N__38917\,
            I => \N__38914\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38911\
        );

    \I__8251\ : Span4Mux_h
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__38908\,
            I => \ALU.r0_12_prm_8_8_s0_c_RNOZ0\
        );

    \I__8249\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38902\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__38902\,
            I => \N__38899\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__38899\,
            I => \N__38896\
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__38896\,
            I => \ALU.r0_12_prm_8_12_s1_c_RNOZ0Z_1\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38893\,
            I => \N__38890\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38890\,
            I => \N__38887\
        );

    \I__8243\ : Odrv4
    port map (
            O => \N__38887\,
            I => \ALU.r0_12_prm_7_8_s0_c_RNOZ0\
        );

    \I__8242\ : InMux
    port map (
            O => \N__38884\,
            I => \N__38881\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__38881\,
            I => \ALU.rshift_5\
        );

    \I__8240\ : InMux
    port map (
            O => \N__38878\,
            I => \N__38875\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__38875\,
            I => \N__38868\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38865\
        );

    \I__8237\ : InMux
    port map (
            O => \N__38873\,
            I => \N__38862\
        );

    \I__8236\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38859\
        );

    \I__8235\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38856\
        );

    \I__8234\ : Span4Mux_v
    port map (
            O => \N__38868\,
            I => \N__38850\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__38865\,
            I => \N__38850\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__38862\,
            I => \N__38845\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38859\,
            I => \N__38845\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__38856\,
            I => \N__38842\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38839\
        );

    \I__8228\ : Span4Mux_h
    port map (
            O => \N__38850\,
            I => \N__38836\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__38845\,
            I => \N__38833\
        );

    \I__8226\ : Span4Mux_h
    port map (
            O => \N__38842\,
            I => \N__38828\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__38839\,
            I => \N__38828\
        );

    \I__8224\ : Span4Mux_h
    port map (
            O => \N__38836\,
            I => \N__38824\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__38833\,
            I => \N__38819\
        );

    \I__8222\ : Span4Mux_h
    port map (
            O => \N__38828\,
            I => \N__38819\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38827\,
            I => \N__38816\
        );

    \I__8220\ : Sp12to4
    port map (
            O => \N__38824\,
            I => \N__38808\
        );

    \I__8219\ : Sp12to4
    port map (
            O => \N__38819\,
            I => \N__38808\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38816\,
            I => \N__38808\
        );

    \I__8217\ : InMux
    port map (
            O => \N__38815\,
            I => \N__38805\
        );

    \I__8216\ : Odrv12
    port map (
            O => \N__38808\,
            I => \ALU.r0_12_6\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__38805\,
            I => \ALU.r0_12_6\
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__38800\,
            I => \N__38797\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38797\,
            I => \N__38794\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__38794\,
            I => \N__38790\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38787\
        );

    \I__8210\ : Span4Mux_v
    port map (
            O => \N__38790\,
            I => \N__38783\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38787\,
            I => \N__38780\
        );

    \I__8208\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38777\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__38783\,
            I => \N__38774\
        );

    \I__8206\ : Span4Mux_h
    port map (
            O => \N__38780\,
            I => \N__38771\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__38777\,
            I => \N__38768\
        );

    \I__8204\ : Span4Mux_v
    port map (
            O => \N__38774\,
            I => \N__38761\
        );

    \I__8203\ : Span4Mux_v
    port map (
            O => \N__38771\,
            I => \N__38761\
        );

    \I__8202\ : Span4Mux_h
    port map (
            O => \N__38768\,
            I => \N__38761\
        );

    \I__8201\ : Span4Mux_h
    port map (
            O => \N__38761\,
            I => \N__38758\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__38758\,
            I => r6_6
        );

    \I__8199\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38751\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38748\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38751\,
            I => \N__38742\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__38748\,
            I => \N__38742\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38737\
        );

    \I__8194\ : Span4Mux_v
    port map (
            O => \N__38742\,
            I => \N__38734\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38741\,
            I => \N__38731\
        );

    \I__8192\ : InMux
    port map (
            O => \N__38740\,
            I => \N__38728\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__38737\,
            I => \N__38724\
        );

    \I__8190\ : Span4Mux_h
    port map (
            O => \N__38734\,
            I => \N__38719\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__38731\,
            I => \N__38719\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38728\,
            I => \N__38716\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38727\,
            I => \N__38713\
        );

    \I__8186\ : Span4Mux_v
    port map (
            O => \N__38724\,
            I => \N__38708\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__38719\,
            I => \N__38705\
        );

    \I__8184\ : Span12Mux_v
    port map (
            O => \N__38716\,
            I => \N__38700\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38700\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38697\
        );

    \I__8181\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38694\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__38708\,
            I => \ALU.r0_12_7\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__38705\,
            I => \ALU.r0_12_7\
        );

    \I__8178\ : Odrv12
    port map (
            O => \N__38700\,
            I => \ALU.r0_12_7\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38697\,
            I => \ALU.r0_12_7\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38694\,
            I => \ALU.r0_12_7\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38683\,
            I => \N__38674\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38674\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38674\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38674\,
            I => \N__38671\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__38671\,
            I => \N__38668\
        );

    \I__8170\ : Span4Mux_h
    port map (
            O => \N__38668\,
            I => \N__38665\
        );

    \I__8169\ : Span4Mux_h
    port map (
            O => \N__38665\,
            I => \N__38662\
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__38662\,
            I => r6_7
        );

    \I__8167\ : InMux
    port map (
            O => \N__38659\,
            I => \ALU.r0_12_4\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38656\,
            I => \N__38653\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__38653\,
            I => \N__38650\
        );

    \I__8164\ : Span4Mux_v
    port map (
            O => \N__38650\,
            I => \N__38646\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38643\
        );

    \I__8162\ : Sp12to4
    port map (
            O => \N__38646\,
            I => \N__38640\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38643\,
            I => \N__38637\
        );

    \I__8160\ : Odrv12
    port map (
            O => \N__38640\,
            I => \ALU.r5_RNIKS4A9Z0Z_11\
        );

    \I__8159\ : Odrv4
    port map (
            O => \N__38637\,
            I => \ALU.r5_RNIKS4A9Z0Z_11\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38632\,
            I => \N__38628\
        );

    \I__8157\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38625\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__38628\,
            I => \N__38622\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__38625\,
            I => \ALU.r4_RNIVLAIAZ0Z_9\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__38622\,
            I => \ALU.r4_RNIVLAIAZ0Z_9\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38617\,
            I => \ALU.r5_RNI0QK3KZ0Z_11_cascade_\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38614\,
            I => \N__38611\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38611\,
            I => \N__38608\
        );

    \I__8150\ : Span4Mux_v
    port map (
            O => \N__38608\,
            I => \N__38605\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__38605\,
            I => \ALU.rshift_8\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38602\,
            I => \N__38599\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__38599\,
            I => \N__38595\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38598\,
            I => \N__38592\
        );

    \I__8145\ : Span4Mux_h
    port map (
            O => \N__38595\,
            I => \N__38589\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__38592\,
            I => \N__38586\
        );

    \I__8143\ : Span4Mux_v
    port map (
            O => \N__38589\,
            I => \N__38581\
        );

    \I__8142\ : Span4Mux_v
    port map (
            O => \N__38586\,
            I => \N__38581\
        );

    \I__8141\ : Odrv4
    port map (
            O => \N__38581\,
            I => \ALU.un2_addsub_cry_3_c_RNI8MVBGZ0\
        );

    \I__8140\ : CascadeMux
    port map (
            O => \N__38578\,
            I => \N__38575\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38572\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38572\,
            I => \ALU.r0_12_prm_2_4_c_RNOZ0\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38566\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__38566\,
            I => \N__38563\
        );

    \I__8135\ : Span4Mux_v
    port map (
            O => \N__38563\,
            I => \N__38560\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__38560\,
            I => \N__38556\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38553\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__38556\,
            I => \ALU.madd_axb_3\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38553\,
            I => \ALU.madd_axb_3\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38545\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__38545\,
            I => \N__38541\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38544\,
            I => \N__38538\
        );

    \I__8127\ : Span4Mux_h
    port map (
            O => \N__38541\,
            I => \N__38535\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__38538\,
            I => \ALU.madd_cry_2_THRU_CO\
        );

    \I__8125\ : Odrv4
    port map (
            O => \N__38535\,
            I => \ALU.madd_cry_2_THRU_CO\
        );

    \I__8124\ : InMux
    port map (
            O => \N__38530\,
            I => \N__38527\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38527\,
            I => \ALU.r0_12_prm_3_4_c_RNOZ0\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38521\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38516\
        );

    \I__8120\ : CascadeMux
    port map (
            O => \N__38520\,
            I => \N__38513\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38510\
        );

    \I__8118\ : Span4Mux_v
    port map (
            O => \N__38516\,
            I => \N__38507\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38504\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__38510\,
            I => \N__38501\
        );

    \I__8115\ : Span4Mux_h
    port map (
            O => \N__38507\,
            I => \N__38498\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38504\,
            I => \N__38495\
        );

    \I__8113\ : Span4Mux_v
    port map (
            O => \N__38501\,
            I => \N__38492\
        );

    \I__8112\ : Span4Mux_h
    port map (
            O => \N__38498\,
            I => \N__38489\
        );

    \I__8111\ : Span4Mux_h
    port map (
            O => \N__38495\,
            I => \N__38486\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__38492\,
            I => \N__38483\
        );

    \I__8109\ : Sp12to4
    port map (
            O => \N__38489\,
            I => \N__38480\
        );

    \I__8108\ : Span4Mux_h
    port map (
            O => \N__38486\,
            I => \N__38477\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__38483\,
            I => \N__38474\
        );

    \I__8106\ : Odrv12
    port map (
            O => \N__38480\,
            I => r1_6
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__38477\,
            I => r1_6
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__38474\,
            I => r1_6
        );

    \I__8103\ : InMux
    port map (
            O => \N__38467\,
            I => \N__38464\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__38464\,
            I => \N__38460\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38457\
        );

    \I__8100\ : Span4Mux_h
    port map (
            O => \N__38460\,
            I => \N__38452\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38457\,
            I => \N__38452\
        );

    \I__8098\ : Span4Mux_v
    port map (
            O => \N__38452\,
            I => \N__38448\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__38451\,
            I => \N__38445\
        );

    \I__8096\ : Span4Mux_h
    port map (
            O => \N__38448\,
            I => \N__38442\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38445\,
            I => \N__38439\
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__38442\,
            I => \ALU.a4_b_4\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38439\,
            I => \ALU.a4_b_4\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__38434\,
            I => \N__38431\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38428\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38428\,
            I => \ALU.r0_12_prm_7_4_c_RNOZ0\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38422\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38422\,
            I => \N__38419\
        );

    \I__8087\ : Span4Mux_v
    port map (
            O => \N__38419\,
            I => \N__38416\
        );

    \I__8086\ : Span4Mux_h
    port map (
            O => \N__38416\,
            I => \N__38413\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__38413\,
            I => \ALU.r0_12_prm_6_4_c_RNOZ0\
        );

    \I__8084\ : CascadeMux
    port map (
            O => \N__38410\,
            I => \N__38407\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38404\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__38404\,
            I => \N__38401\
        );

    \I__8081\ : Span4Mux_h
    port map (
            O => \N__38401\,
            I => \N__38398\
        );

    \I__8080\ : Odrv4
    port map (
            O => \N__38398\,
            I => \ALU.un14_log_0_i_4\
        );

    \I__8079\ : CascadeMux
    port map (
            O => \N__38395\,
            I => \N__38392\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38392\,
            I => \N__38389\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38389\,
            I => \N__38386\
        );

    \I__8076\ : Odrv4
    port map (
            O => \N__38386\,
            I => \ALU.r0_12_prm_5_4_c_RNOZ0Z_0\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38383\,
            I => \N__38380\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__38380\,
            I => \ALU.a_i_4\
        );

    \I__8073\ : CascadeMux
    port map (
            O => \N__38377\,
            I => \N__38374\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38371\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38368\
        );

    \I__8070\ : Odrv12
    port map (
            O => \N__38368\,
            I => \ALU.mult_4\
        );

    \I__8069\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38362\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__38362\,
            I => \N__38358\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__38361\,
            I => \N__38355\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__38358\,
            I => \N__38352\
        );

    \I__8065\ : InMux
    port map (
            O => \N__38355\,
            I => \N__38349\
        );

    \I__8064\ : Sp12to4
    port map (
            O => \N__38352\,
            I => \N__38344\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__38349\,
            I => \N__38344\
        );

    \I__8062\ : Odrv12
    port map (
            O => \N__38344\,
            I => \ALU.un14_log_0_i_6\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38337\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__38340\,
            I => \N__38334\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38337\,
            I => \N__38331\
        );

    \I__8058\ : InMux
    port map (
            O => \N__38334\,
            I => \N__38328\
        );

    \I__8057\ : Span4Mux_v
    port map (
            O => \N__38331\,
            I => \N__38325\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__38328\,
            I => \N__38322\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__38325\,
            I => \ALU.r4_RNI2BKQ8_0Z0Z_6\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__38322\,
            I => \ALU.r4_RNI2BKQ8_0Z0Z_6\
        );

    \I__8053\ : CascadeMux
    port map (
            O => \N__38317\,
            I => \N__38314\
        );

    \I__8052\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38311\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__38311\,
            I => \N__38308\
        );

    \I__8050\ : Span4Mux_h
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__8049\ : IoSpan4Mux
    port map (
            O => \N__38305\,
            I => \N__38302\
        );

    \I__8048\ : Span4Mux_s0_v
    port map (
            O => \N__38302\,
            I => \N__38299\
        );

    \I__8047\ : Odrv4
    port map (
            O => \N__38299\,
            I => \ALU.r4_RNIUGHG5Z0Z_6\
        );

    \I__8046\ : CascadeMux
    port map (
            O => \N__38296\,
            I => \N__38293\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38293\,
            I => \N__38290\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__38290\,
            I => \N__38286\
        );

    \I__8043\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38283\
        );

    \I__8042\ : Span4Mux_s2_v
    port map (
            O => \N__38286\,
            I => \N__38280\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__38283\,
            I => \ALU.a_i_6\
        );

    \I__8040\ : Odrv4
    port map (
            O => \N__38280\,
            I => \ALU.a_i_6\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38272\,
            I => \N__38269\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__38269\,
            I => \ALU.r0_12_prm_3_6_s0_sf\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38266\,
            I => \N__38262\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38259\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__38262\,
            I => \N__38254\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__38259\,
            I => \N__38251\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38248\
        );

    \I__8031\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38245\
        );

    \I__8030\ : Span4Mux_s1_v
    port map (
            O => \N__38254\,
            I => \N__38242\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__38251\,
            I => \N__38239\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38236\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38233\
        );

    \I__8026\ : Span4Mux_v
    port map (
            O => \N__38242\,
            I => \N__38230\
        );

    \I__8025\ : Span4Mux_v
    port map (
            O => \N__38239\,
            I => \N__38227\
        );

    \I__8024\ : Span12Mux_h
    port map (
            O => \N__38236\,
            I => \N__38222\
        );

    \I__8023\ : Span12Mux_s2_v
    port map (
            O => \N__38233\,
            I => \N__38222\
        );

    \I__8022\ : Odrv4
    port map (
            O => \N__38230\,
            I => \ALU.un2_addsub_cry_5_c_RNIO30SDZ0\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__38227\,
            I => \ALU.un2_addsub_cry_5_c_RNIO30SDZ0\
        );

    \I__8020\ : Odrv12
    port map (
            O => \N__38222\,
            I => \ALU.un2_addsub_cry_5_c_RNIO30SDZ0\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__38215\,
            I => \N__38212\
        );

    \I__8018\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38209\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__38209\,
            I => \ALU.r0_12_prm_2_6_s0_c_RNOZ0\
        );

    \I__8016\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38201\
        );

    \I__8015\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38198\
        );

    \I__8014\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38195\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__38201\,
            I => \N__38192\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__38198\,
            I => \N__38189\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__38195\,
            I => \N__38186\
        );

    \I__8010\ : Span4Mux_s0_v
    port map (
            O => \N__38192\,
            I => \N__38182\
        );

    \I__8009\ : Span12Mux_s7_v
    port map (
            O => \N__38189\,
            I => \N__38179\
        );

    \I__8008\ : Span4Mux_v
    port map (
            O => \N__38186\,
            I => \N__38176\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38173\
        );

    \I__8006\ : Span4Mux_v
    port map (
            O => \N__38182\,
            I => \N__38170\
        );

    \I__8005\ : Odrv12
    port map (
            O => \N__38179\,
            I => \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019\
        );

    \I__8004\ : Odrv4
    port map (
            O => \N__38176\,
            I => \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38173\,
            I => \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__38170\,
            I => \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__38161\,
            I => \N__38158\
        );

    \I__8000\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38155\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__38155\,
            I => \N__38152\
        );

    \I__7998\ : Span4Mux_v
    port map (
            O => \N__38152\,
            I => \N__38149\
        );

    \I__7997\ : Odrv4
    port map (
            O => \N__38149\,
            I => \ALU.r0_12_prm_1_6_s0_c_RNOZ0\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38146\,
            I => \N__38143\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38143\,
            I => \N__38140\
        );

    \I__7994\ : Span4Mux_h
    port map (
            O => \N__38140\,
            I => \N__38137\
        );

    \I__7993\ : Odrv4
    port map (
            O => \N__38137\,
            I => \ALU.r0_12_s1_6_THRU_CO\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38134\,
            I => \N__38131\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__38131\,
            I => \N__38128\
        );

    \I__7990\ : Span4Mux_h
    port map (
            O => \N__38128\,
            I => \N__38125\
        );

    \I__7989\ : Span4Mux_h
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__7988\ : Odrv4
    port map (
            O => \N__38122\,
            I => \ALU.mult_6\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38119\,
            I => \ALU.r0_12_s0_6\
        );

    \I__7986\ : InMux
    port map (
            O => \N__38116\,
            I => \N__38113\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__38113\,
            I => \ALU.r0_12_prm_2_0_s1_c_RNOZ0\
        );

    \I__7984\ : InMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__7982\ : Span4Mux_h
    port map (
            O => \N__38104\,
            I => \N__38101\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__38101\,
            I => \ALU.r0_12_prm_8_2_c_RNOZ0Z_3\
        );

    \I__7980\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38095\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__38095\,
            I => \N__38092\
        );

    \I__7978\ : Span4Mux_h
    port map (
            O => \N__38092\,
            I => \N__38089\
        );

    \I__7977\ : Span4Mux_s1_v
    port map (
            O => \N__38089\,
            I => \N__38086\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__38086\,
            I => \ALU.r4_RNI1G9PKZ0Z_6\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38080\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__38077\
        );

    \I__7973\ : Span4Mux_s3_v
    port map (
            O => \N__38077\,
            I => \N__38072\
        );

    \I__7972\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38067\
        );

    \I__7971\ : InMux
    port map (
            O => \N__38075\,
            I => \N__38067\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__38072\,
            I => \ALU.N_845_1\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__38067\,
            I => \ALU.N_845_1\
        );

    \I__7968\ : CascadeMux
    port map (
            O => \N__38062\,
            I => \ALU.rshift_15_ns_1_2_cascade_\
        );

    \I__7967\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38056\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__38056\,
            I => \N__38053\
        );

    \I__7965\ : Span4Mux_h
    port map (
            O => \N__38053\,
            I => \N__38047\
        );

    \I__7964\ : InMux
    port map (
            O => \N__38052\,
            I => \N__38044\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38051\,
            I => \N__38039\
        );

    \I__7962\ : InMux
    port map (
            O => \N__38050\,
            I => \N__38039\
        );

    \I__7961\ : Odrv4
    port map (
            O => \N__38047\,
            I => \ALU.r5_RNI8R2TIZ0Z_11\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__38044\,
            I => \ALU.r5_RNI8R2TIZ0Z_11\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__38039\,
            I => \ALU.r5_RNI8R2TIZ0Z_11\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38032\,
            I => \N__38022\
        );

    \I__7957\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38012\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38009\
        );

    \I__7955\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38002\
        );

    \I__7954\ : InMux
    port map (
            O => \N__38028\,
            I => \N__38002\
        );

    \I__7953\ : InMux
    port map (
            O => \N__38027\,
            I => \N__37995\
        );

    \I__7952\ : InMux
    port map (
            O => \N__38026\,
            I => \N__37995\
        );

    \I__7951\ : InMux
    port map (
            O => \N__38025\,
            I => \N__37995\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__38022\,
            I => \N__37989\
        );

    \I__7949\ : InMux
    port map (
            O => \N__38021\,
            I => \N__37985\
        );

    \I__7948\ : InMux
    port map (
            O => \N__38020\,
            I => \N__37982\
        );

    \I__7947\ : InMux
    port map (
            O => \N__38019\,
            I => \N__37977\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38018\,
            I => \N__37977\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38017\,
            I => \N__37974\
        );

    \I__7944\ : InMux
    port map (
            O => \N__38016\,
            I => \N__37970\
        );

    \I__7943\ : InMux
    port map (
            O => \N__38015\,
            I => \N__37961\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__38012\,
            I => \N__37955\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__38009\,
            I => \N__37955\
        );

    \I__7940\ : InMux
    port map (
            O => \N__38008\,
            I => \N__37950\
        );

    \I__7939\ : InMux
    port map (
            O => \N__38007\,
            I => \N__37950\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__38002\,
            I => \N__37945\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__37995\,
            I => \N__37945\
        );

    \I__7936\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37938\
        );

    \I__7935\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37938\
        );

    \I__7934\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37938\
        );

    \I__7933\ : Span4Mux_s3_v
    port map (
            O => \N__37989\,
            I => \N__37935\
        );

    \I__7932\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37932\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__37985\,
            I => \N__37929\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37982\,
            I => \N__37924\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__37977\,
            I => \N__37924\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__37974\,
            I => \N__37921\
        );

    \I__7927\ : InMux
    port map (
            O => \N__37973\,
            I => \N__37918\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__37970\,
            I => \N__37915\
        );

    \I__7925\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37908\
        );

    \I__7924\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37908\
        );

    \I__7923\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37908\
        );

    \I__7922\ : InMux
    port map (
            O => \N__37966\,
            I => \N__37903\
        );

    \I__7921\ : InMux
    port map (
            O => \N__37965\,
            I => \N__37903\
        );

    \I__7920\ : InMux
    port map (
            O => \N__37964\,
            I => \N__37900\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__37961\,
            I => \N__37892\
        );

    \I__7918\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37889\
        );

    \I__7917\ : Span4Mux_h
    port map (
            O => \N__37955\,
            I => \N__37875\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37950\,
            I => \N__37875\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__37945\,
            I => \N__37875\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37875\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__37935\,
            I => \N__37870\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__37932\,
            I => \N__37870\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__37929\,
            I => \N__37867\
        );

    \I__7910\ : Span4Mux_s3_v
    port map (
            O => \N__37924\,
            I => \N__37860\
        );

    \I__7909\ : Span4Mux_s1_h
    port map (
            O => \N__37921\,
            I => \N__37860\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__37918\,
            I => \N__37860\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__37915\,
            I => \N__37855\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__37908\,
            I => \N__37855\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__37903\,
            I => \N__37852\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__37900\,
            I => \N__37849\
        );

    \I__7903\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37842\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37842\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37842\
        );

    \I__7900\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37837\
        );

    \I__7899\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37837\
        );

    \I__7898\ : Sp12to4
    port map (
            O => \N__37892\,
            I => \N__37832\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__37889\,
            I => \N__37832\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37823\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37814\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37814\
        );

    \I__7893\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37814\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37814\
        );

    \I__7891\ : Span4Mux_h
    port map (
            O => \N__37875\,
            I => \N__37811\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__37870\,
            I => \N__37804\
        );

    \I__7889\ : Span4Mux_h
    port map (
            O => \N__37867\,
            I => \N__37804\
        );

    \I__7888\ : Span4Mux_h
    port map (
            O => \N__37860\,
            I => \N__37804\
        );

    \I__7887\ : Span4Mux_h
    port map (
            O => \N__37855\,
            I => \N__37799\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__37852\,
            I => \N__37799\
        );

    \I__7885\ : Span4Mux_h
    port map (
            O => \N__37849\,
            I => \N__37794\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__37842\,
            I => \N__37794\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__37837\,
            I => \N__37789\
        );

    \I__7882\ : Span12Mux_v
    port map (
            O => \N__37832\,
            I => \N__37789\
        );

    \I__7881\ : InMux
    port map (
            O => \N__37831\,
            I => \N__37784\
        );

    \I__7880\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37784\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37775\
        );

    \I__7878\ : InMux
    port map (
            O => \N__37828\,
            I => \N__37775\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37827\,
            I => \N__37775\
        );

    \I__7876\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37775\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37823\,
            I => \ALU.bZ0Z_0\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__37814\,
            I => \ALU.bZ0Z_0\
        );

    \I__7873\ : Odrv4
    port map (
            O => \N__37811\,
            I => \ALU.bZ0Z_0\
        );

    \I__7872\ : Odrv4
    port map (
            O => \N__37804\,
            I => \ALU.bZ0Z_0\
        );

    \I__7871\ : Odrv4
    port map (
            O => \N__37799\,
            I => \ALU.bZ0Z_0\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__37794\,
            I => \ALU.bZ0Z_0\
        );

    \I__7869\ : Odrv12
    port map (
            O => \N__37789\,
            I => \ALU.bZ0Z_0\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__37784\,
            I => \ALU.bZ0Z_0\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37775\,
            I => \ALU.bZ0Z_0\
        );

    \I__7866\ : InMux
    port map (
            O => \N__37756\,
            I => \N__37753\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__37753\,
            I => \N__37749\
        );

    \I__7864\ : CascadeMux
    port map (
            O => \N__37752\,
            I => \N__37746\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__37749\,
            I => \N__37743\
        );

    \I__7862\ : InMux
    port map (
            O => \N__37746\,
            I => \N__37740\
        );

    \I__7861\ : Odrv4
    port map (
            O => \N__37743\,
            I => \ALU.r4_RNID26E8_0Z0Z_0\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__37740\,
            I => \ALU.r4_RNID26E8_0Z0Z_0\
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__37735\,
            I => \N__37731\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__37734\,
            I => \N__37727\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37723\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37720\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37717\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37714\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37723\,
            I => \N__37709\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__37720\,
            I => \N__37709\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37717\,
            I => \N__37704\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37714\,
            I => \N__37704\
        );

    \I__7849\ : Span4Mux_h
    port map (
            O => \N__37709\,
            I => \N__37701\
        );

    \I__7848\ : Span4Mux_s0_v
    port map (
            O => \N__37704\,
            I => \N__37698\
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__37701\,
            I => \ALU.rshift_6\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__37698\,
            I => \ALU.rshift_6\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37690\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__37690\,
            I => \N__37685\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__37689\,
            I => \N__37682\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37679\
        );

    \I__7841\ : Span4Mux_h
    port map (
            O => \N__37685\,
            I => \N__37676\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37673\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__37679\,
            I => \N__37670\
        );

    \I__7838\ : Odrv4
    port map (
            O => \N__37676\,
            I => \ALU.lshift_6\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__37673\,
            I => \ALU.lshift_6\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__37670\,
            I => \ALU.lshift_6\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__37663\,
            I => \N__37660\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37657\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37657\,
            I => \ALU.r0_12_prm_8_6_s0_c_RNOZ0\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37651\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37651\,
            I => \N__37647\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37644\
        );

    \I__7829\ : Span4Mux_v
    port map (
            O => \N__37647\,
            I => \N__37641\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37644\,
            I => \N__37638\
        );

    \I__7827\ : Span4Mux_h
    port map (
            O => \N__37641\,
            I => \N__37633\
        );

    \I__7826\ : Span4Mux_h
    port map (
            O => \N__37638\,
            I => \N__37630\
        );

    \I__7825\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37627\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37624\
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__37633\,
            I => \ALU.un2_addsub_cry_11_c_RNICP8AEZ0\
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__37630\,
            I => \ALU.un2_addsub_cry_11_c_RNICP8AEZ0\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__37627\,
            I => \ALU.un2_addsub_cry_11_c_RNICP8AEZ0\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37624\,
            I => \ALU.un2_addsub_cry_11_c_RNICP8AEZ0\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__37615\,
            I => \N__37612\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37612\,
            I => \N__37609\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37609\,
            I => \N__37606\
        );

    \I__7816\ : Odrv4
    port map (
            O => \N__37606\,
            I => \ALU.r0_12_prm_2_12_s1_c_RNOZ0\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37600\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__37600\,
            I => \N__37597\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__37597\,
            I => \ALU.r0_12_prm_1_12_s1_c_RNOZ0\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37590\
        );

    \I__7811\ : CascadeMux
    port map (
            O => \N__37593\,
            I => \N__37587\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37590\,
            I => \N__37583\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37580\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37586\,
            I => \N__37577\
        );

    \I__7807\ : Span4Mux_v
    port map (
            O => \N__37583\,
            I => \N__37573\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37580\,
            I => \N__37568\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37577\,
            I => \N__37568\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37576\,
            I => \N__37565\
        );

    \I__7803\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37558\
        );

    \I__7802\ : Span4Mux_v
    port map (
            O => \N__37568\,
            I => \N__37558\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37558\
        );

    \I__7800\ : Odrv4
    port map (
            O => \N__37558\,
            I => \ALU.un9_addsub_cry_11_c_RNIAHI1AZ0\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37555\,
            I => \ALU.r0_12_s1_12\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37549\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37549\,
            I => \N__37546\
        );

    \I__7796\ : Span12Mux_v
    port map (
            O => \N__37546\,
            I => \N__37543\
        );

    \I__7795\ : Odrv12
    port map (
            O => \N__37543\,
            I => \ALU.r0_12_s1_12_THRU_CO\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__37540\,
            I => \N__37537\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37534\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37534\,
            I => \N__37531\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__37531\,
            I => \N__37528\
        );

    \I__7790\ : Span4Mux_h
    port map (
            O => \N__37528\,
            I => \N__37525\
        );

    \I__7789\ : Span4Mux_h
    port map (
            O => \N__37525\,
            I => \N__37522\
        );

    \I__7788\ : Odrv4
    port map (
            O => \N__37522\,
            I => \ALU.r0_12_prm_5_15_s1_c_RNOZ0\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37519\,
            I => \N__37516\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37516\,
            I => \N__37513\
        );

    \I__7785\ : Span12Mux_s7_h
    port map (
            O => \N__37513\,
            I => \N__37510\
        );

    \I__7784\ : Span12Mux_v
    port map (
            O => \N__37510\,
            I => \N__37507\
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__37507\,
            I => \ALU.r0_12_prm_8_15_s1_c_RNOZ0Z_1\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37504\,
            I => \N__37501\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37501\,
            I => \ALU.r0_12_prm_8_0_s1_c_RNOZ0\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37498\,
            I => \N__37495\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37495\,
            I => \N__37492\
        );

    \I__7778\ : Span4Mux_h
    port map (
            O => \N__37492\,
            I => \N__37489\
        );

    \I__7777\ : Odrv4
    port map (
            O => \N__37489\,
            I => \ALU.r5_RNIAV175Z0Z_15\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37482\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37479\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37482\,
            I => \ALU.r4_RNIQK1V71Z0Z_5\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37479\,
            I => \ALU.r4_RNIQK1V71Z0Z_5\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37471\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37471\,
            I => \ALU.r0_12_prm_8_12_s1_c_RNOZ0\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37465\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37465\,
            I => \N__37461\
        );

    \I__7768\ : CascadeMux
    port map (
            O => \N__37464\,
            I => \N__37458\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__37461\,
            I => \N__37455\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37452\
        );

    \I__7765\ : Odrv4
    port map (
            O => \N__37455\,
            I => \ALU.lshift_12\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37452\,
            I => \ALU.lshift_12\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37447\,
            I => \N__37444\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37444\,
            I => \ALU.r0_12_prm_7_12_s1_c_RNOZ0\
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__37441\,
            I => \N__37438\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37434\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37431\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37428\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37425\
        );

    \I__7756\ : Span4Mux_v
    port map (
            O => \N__37428\,
            I => \N__37422\
        );

    \I__7755\ : Span4Mux_v
    port map (
            O => \N__37425\,
            I => \N__37417\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__37422\,
            I => \N__37417\
        );

    \I__7753\ : Odrv4
    port map (
            O => \N__37417\,
            I => \ALU.r5_RNISP2L9_0Z0Z_12\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37414\,
            I => \N__37411\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37411\,
            I => \N__37407\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37410\,
            I => \N__37404\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__37407\,
            I => \N__37401\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__37404\,
            I => \N__37398\
        );

    \I__7747\ : Sp12to4
    port map (
            O => \N__37401\,
            I => \N__37395\
        );

    \I__7746\ : Span4Mux_h
    port map (
            O => \N__37398\,
            I => \N__37392\
        );

    \I__7745\ : Span12Mux_v
    port map (
            O => \N__37395\,
            I => \N__37389\
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__37392\,
            I => \ALU.un14_log_0_i_12\
        );

    \I__7743\ : Odrv12
    port map (
            O => \N__37389\,
            I => \ALU.un14_log_0_i_12\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37381\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__37381\,
            I => \N__37378\
        );

    \I__7740\ : Span4Mux_h
    port map (
            O => \N__37378\,
            I => \N__37375\
        );

    \I__7739\ : Span4Mux_v
    port map (
            O => \N__37375\,
            I => \N__37372\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__37372\,
            I => \ALU.r0_12_prm_5_12_s1_c_RNOZ0\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37366\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37366\,
            I => \N__37363\
        );

    \I__7735\ : Span4Mux_h
    port map (
            O => \N__37363\,
            I => \N__37359\
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__37362\,
            I => \N__37356\
        );

    \I__7733\ : Span4Mux_h
    port map (
            O => \N__37359\,
            I => \N__37353\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37350\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__37353\,
            I => \ALU.r5_RNISP2L9_1Z0Z_12\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__37350\,
            I => \ALU.r5_RNISP2L9_1Z0Z_12\
        );

    \I__7729\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37342\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__37342\,
            I => \N__37339\
        );

    \I__7727\ : Span4Mux_v
    port map (
            O => \N__37339\,
            I => \N__37336\
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__37336\,
            I => \ALU.r0_12_prm_4_12_s1_c_RNOZ0\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__37333\,
            I => \N__37330\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37327\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__37327\,
            I => \N__37324\
        );

    \I__7722\ : Span4Mux_h
    port map (
            O => \N__37324\,
            I => \N__37320\
        );

    \I__7721\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37317\
        );

    \I__7720\ : Span4Mux_h
    port map (
            O => \N__37320\,
            I => \N__37314\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__37317\,
            I => \ALU.a_i_12\
        );

    \I__7718\ : Odrv4
    port map (
            O => \N__37314\,
            I => \ALU.a_i_12\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37309\,
            I => \ALU.r0_12_s0_8\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__37306\,
            I => \N__37303\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37300\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37300\,
            I => \ALU.r0_12_prm_1_8_s0_c_RNOZ0\
        );

    \I__7713\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37294\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37294\,
            I => \N__37291\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__37291\,
            I => \N__37287\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__37290\,
            I => \N__37284\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__37287\,
            I => \N__37280\
        );

    \I__7708\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37277\
        );

    \I__7707\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37274\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__37280\,
            I => \N__37270\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__37277\,
            I => \N__37267\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__37274\,
            I => \N__37264\
        );

    \I__7703\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37261\
        );

    \I__7702\ : Odrv4
    port map (
            O => \N__37270\,
            I => \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9\
        );

    \I__7701\ : Odrv12
    port map (
            O => \N__37267\,
            I => \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9\
        );

    \I__7700\ : Odrv4
    port map (
            O => \N__37264\,
            I => \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__37261\,
            I => \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__37252\,
            I => \N__37249\
        );

    \I__7697\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37246\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__37246\,
            I => \N__37243\
        );

    \I__7695\ : Span4Mux_h
    port map (
            O => \N__37243\,
            I => \N__37240\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__37240\,
            I => \N__37237\
        );

    \I__7693\ : Odrv4
    port map (
            O => \N__37237\,
            I => \ALU.r0_12_prm_1_15_s1_c_RNOZ0\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37231\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37231\,
            I => \N__37228\
        );

    \I__7690\ : Span4Mux_h
    port map (
            O => \N__37228\,
            I => \N__37225\
        );

    \I__7689\ : Span4Mux_h
    port map (
            O => \N__37225\,
            I => \N__37222\
        );

    \I__7688\ : Odrv4
    port map (
            O => \N__37222\,
            I => \ALU.mult_5\
        );

    \I__7687\ : InMux
    port map (
            O => \N__37219\,
            I => \ALU.r0_12_s0_5\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37213\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__37213\,
            I => \N__37205\
        );

    \I__7684\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37202\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37199\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37210\,
            I => \N__37196\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37193\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37208\,
            I => \N__37190\
        );

    \I__7679\ : Span4Mux_v
    port map (
            O => \N__37205\,
            I => \N__37180\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__37202\,
            I => \N__37180\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__37199\,
            I => \N__37180\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37180\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__37193\,
            I => \N__37177\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37190\,
            I => \N__37174\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37171\
        );

    \I__7672\ : Span4Mux_v
    port map (
            O => \N__37180\,
            I => \N__37168\
        );

    \I__7671\ : Span4Mux_h
    port map (
            O => \N__37177\,
            I => \N__37165\
        );

    \I__7670\ : Span4Mux_v
    port map (
            O => \N__37174\,
            I => \N__37160\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__37171\,
            I => \N__37160\
        );

    \I__7668\ : Span4Mux_h
    port map (
            O => \N__37168\,
            I => \N__37157\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__37165\,
            I => \N__37154\
        );

    \I__7666\ : Span4Mux_v
    port map (
            O => \N__37160\,
            I => \N__37151\
        );

    \I__7665\ : Span4Mux_h
    port map (
            O => \N__37157\,
            I => \N__37147\
        );

    \I__7664\ : Span4Mux_h
    port map (
            O => \N__37154\,
            I => \N__37144\
        );

    \I__7663\ : Span4Mux_h
    port map (
            O => \N__37151\,
            I => \N__37141\
        );

    \I__7662\ : InMux
    port map (
            O => \N__37150\,
            I => \N__37138\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__37147\,
            I => \ALU.r0_12_5\
        );

    \I__7660\ : Odrv4
    port map (
            O => \N__37144\,
            I => \ALU.r0_12_5\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__37141\,
            I => \ALU.r0_12_5\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__37138\,
            I => \ALU.r0_12_5\
        );

    \I__7657\ : CascadeMux
    port map (
            O => \N__37129\,
            I => \N__37126\
        );

    \I__7656\ : InMux
    port map (
            O => \N__37126\,
            I => \N__37121\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37118\
        );

    \I__7654\ : CascadeMux
    port map (
            O => \N__37124\,
            I => \N__37115\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37112\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__37118\,
            I => \N__37109\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37106\
        );

    \I__7650\ : Span4Mux_v
    port map (
            O => \N__37112\,
            I => \N__37103\
        );

    \I__7649\ : Sp12to4
    port map (
            O => \N__37109\,
            I => \N__37100\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37097\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__37103\,
            I => \N__37094\
        );

    \I__7646\ : Span12Mux_v
    port map (
            O => \N__37100\,
            I => \N__37089\
        );

    \I__7645\ : Span12Mux_s5_h
    port map (
            O => \N__37097\,
            I => \N__37089\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__37094\,
            I => r1_5
        );

    \I__7643\ : Odrv12
    port map (
            O => \N__37089\,
            I => r1_5
        );

    \I__7642\ : InMux
    port map (
            O => \N__37084\,
            I => \N__37081\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__37081\,
            I => \N__37078\
        );

    \I__7640\ : Span4Mux_v
    port map (
            O => \N__37078\,
            I => \N__37075\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__37075\,
            I => \N__37072\
        );

    \I__7638\ : Span4Mux_h
    port map (
            O => \N__37072\,
            I => \N__37069\
        );

    \I__7637\ : Odrv4
    port map (
            O => \N__37069\,
            I => \ALU.r0_12_prm_6_8_s0_c_RNOZ0\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37066\,
            I => \N__37063\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__37063\,
            I => \ALU.r0_12_prm_3_8_s0_sf\
        );

    \I__7634\ : CascadeMux
    port map (
            O => \N__37060\,
            I => \N__37057\
        );

    \I__7633\ : InMux
    port map (
            O => \N__37057\,
            I => \N__37054\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__37054\,
            I => \N__37051\
        );

    \I__7631\ : Span4Mux_v
    port map (
            O => \N__37051\,
            I => \N__37048\
        );

    \I__7630\ : Sp12to4
    port map (
            O => \N__37048\,
            I => \N__37045\
        );

    \I__7629\ : Odrv12
    port map (
            O => \N__37045\,
            I => \ALU.r0_12_prm_7_5_s0_c_RNOZ0\
        );

    \I__7628\ : CascadeMux
    port map (
            O => \N__37042\,
            I => \N__37039\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37039\,
            I => \N__37036\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__37036\,
            I => \N__37033\
        );

    \I__7625\ : Span4Mux_v
    port map (
            O => \N__37033\,
            I => \N__37030\
        );

    \I__7624\ : Span4Mux_h
    port map (
            O => \N__37030\,
            I => \N__37027\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__37027\,
            I => \ALU.r0_12_prm_6_5_s0_c_RNOZ0\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__37024\,
            I => \N__37021\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37021\,
            I => \N__37018\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__7619\ : Odrv12
    port map (
            O => \N__37015\,
            I => \ALU.r0_12_prm_5_5_s0_c_RNOZ0\
        );

    \I__7618\ : CascadeMux
    port map (
            O => \N__37012\,
            I => \N__37009\
        );

    \I__7617\ : InMux
    port map (
            O => \N__37009\,
            I => \N__37006\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37006\,
            I => \N__37003\
        );

    \I__7615\ : Span4Mux_h
    port map (
            O => \N__37003\,
            I => \N__37000\
        );

    \I__7614\ : Span4Mux_v
    port map (
            O => \N__37000\,
            I => \N__36997\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__36997\,
            I => \ALU.r4_RNIM8HG5Z0Z_5\
        );

    \I__7612\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36991\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__36991\,
            I => \ALU.r0_12_prm_3_5_s0_sf\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__36988\,
            I => \N__36985\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36982\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__7607\ : Odrv4
    port map (
            O => \N__36979\,
            I => \ALU.r0_12_prm_2_5_s0_c_RNOZ0\
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__36976\,
            I => \N__36973\
        );

    \I__7605\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36970\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__36970\,
            I => \N__36967\
        );

    \I__7603\ : Odrv4
    port map (
            O => \N__36967\,
            I => \ALU.r0_12_prm_6_7_s0_c_RNOZ0\
        );

    \I__7602\ : CascadeMux
    port map (
            O => \N__36964\,
            I => \N__36961\
        );

    \I__7601\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36958\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__36958\,
            I => \ALU.r4_RNIFR136Z0Z_7\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36952\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__36952\,
            I => \ALU.r0_12_prm_3_7_s0_sf\
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__36949\,
            I => \N__36946\
        );

    \I__7596\ : InMux
    port map (
            O => \N__36946\,
            I => \N__36943\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36943\,
            I => \ALU.r0_12_prm_1_7_s0_c_RNOZ0\
        );

    \I__7594\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36937\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__36937\,
            I => \N__36934\
        );

    \I__7592\ : Span4Mux_v
    port map (
            O => \N__36934\,
            I => \N__36931\
        );

    \I__7591\ : Span4Mux_h
    port map (
            O => \N__36931\,
            I => \N__36928\
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__36928\,
            I => \ALU.mult_7\
        );

    \I__7589\ : InMux
    port map (
            O => \N__36925\,
            I => \ALU.r0_12_s0_7\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__36922\,
            I => \N__36919\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36914\
        );

    \I__7586\ : InMux
    port map (
            O => \N__36918\,
            I => \N__36909\
        );

    \I__7585\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36909\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__36914\,
            I => \N__36906\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__36909\,
            I => \N__36903\
        );

    \I__7582\ : Span4Mux_h
    port map (
            O => \N__36906\,
            I => \N__36900\
        );

    \I__7581\ : Odrv4
    port map (
            O => \N__36903\,
            I => r1_7
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__36900\,
            I => r1_7
        );

    \I__7579\ : CascadeMux
    port map (
            O => \N__36895\,
            I => \N__36892\
        );

    \I__7578\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36889\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__36889\,
            I => \ALU.lshift_3_ns_1_5\
        );

    \I__7576\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36883\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__36883\,
            I => \N__36880\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__36880\,
            I => \ALU.lshift_15_ns_1_9\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__36877\,
            I => \ALU.r4_RNIF01FKZ0Z_2_cascade_\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36871\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36868\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__36868\,
            I => \N__36864\
        );

    \I__7569\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36861\
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__36864\,
            I => \ALU.r4_RNI2H9PKZ0Z_6\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__36861\,
            I => \ALU.r4_RNI2H9PKZ0Z_6\
        );

    \I__7566\ : CascadeMux
    port map (
            O => \N__36856\,
            I => \ALU.lshift_9_cascade_\
        );

    \I__7565\ : CascadeMux
    port map (
            O => \N__36853\,
            I => \N__36850\
        );

    \I__7564\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36847\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__36847\,
            I => \N__36844\
        );

    \I__7562\ : Span4Mux_v
    port map (
            O => \N__36844\,
            I => \N__36841\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__36841\,
            I => \N__36838\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__36838\,
            I => \ALU.r0_12_prm_8_9_s0_c_RNOZ0\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36835\,
            I => \N__36832\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36832\,
            I => \N__36829\
        );

    \I__7557\ : Odrv4
    port map (
            O => \N__36829\,
            I => \ALU.rshift_15_ns_1_6\
        );

    \I__7556\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36823\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__36823\,
            I => \ALU.rshift_3_ns_1_5\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__36820\,
            I => \ALU.r4_RNI9OH6AZ0Z_1_cascade_\
        );

    \I__7553\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36814\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36814\,
            I => \N__36811\
        );

    \I__7551\ : Span12Mux_s9_v
    port map (
            O => \N__36811\,
            I => \N__36808\
        );

    \I__7550\ : Odrv12
    port map (
            O => \N__36808\,
            I => \ALU.r5_RNIVQN52Z0Z_10\
        );

    \I__7549\ : InMux
    port map (
            O => \N__36805\,
            I => \N__36802\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__36802\,
            I => \N__36799\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__36799\,
            I => \N__36796\
        );

    \I__7546\ : Span4Mux_h
    port map (
            O => \N__36796\,
            I => \N__36792\
        );

    \I__7545\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36789\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__36792\,
            I => \ALU.r6_RNIP3372Z0Z_10\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__36789\,
            I => \ALU.r6_RNIP3372Z0Z_10\
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__36784\,
            I => \N__36779\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__36783\,
            I => \N__36775\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__36782\,
            I => \N__36772\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36779\,
            I => \N__36760\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__36778\,
            I => \N__36756\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36775\,
            I => \N__36750\
        );

    \I__7536\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36747\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__36771\,
            I => \N__36744\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__36770\,
            I => \N__36741\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__36769\,
            I => \N__36738\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__36768\,
            I => \N__36735\
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__36767\,
            I => \N__36731\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__36766\,
            I => \N__36728\
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__36765\,
            I => \N__36725\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36722\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__36763\,
            I => \N__36719\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36760\,
            I => \N__36716\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36759\,
            I => \N__36711\
        );

    \I__7524\ : InMux
    port map (
            O => \N__36756\,
            I => \N__36711\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__36755\,
            I => \N__36708\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__36754\,
            I => \N__36705\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36753\,
            I => \N__36702\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36699\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__36747\,
            I => \N__36694\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36744\,
            I => \N__36689\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36689\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36686\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36682\
        );

    \I__7514\ : InMux
    port map (
            O => \N__36734\,
            I => \N__36677\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36674\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36671\
        );

    \I__7511\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36668\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36665\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36661\
        );

    \I__7508\ : Span4Mux_h
    port map (
            O => \N__36716\,
            I => \N__36656\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__36711\,
            I => \N__36656\
        );

    \I__7506\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36651\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36651\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36648\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__36699\,
            I => \N__36645\
        );

    \I__7502\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36640\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36640\
        );

    \I__7500\ : Span4Mux_s1_v
    port map (
            O => \N__36694\,
            I => \N__36635\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36635\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36686\,
            I => \N__36632\
        );

    \I__7497\ : CascadeMux
    port map (
            O => \N__36685\,
            I => \N__36629\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__36682\,
            I => \N__36626\
        );

    \I__7495\ : CascadeMux
    port map (
            O => \N__36681\,
            I => \N__36622\
        );

    \I__7494\ : CascadeMux
    port map (
            O => \N__36680\,
            I => \N__36618\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36677\,
            I => \N__36615\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36610\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36610\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36607\
        );

    \I__7489\ : Span4Mux_s2_h
    port map (
            O => \N__36665\,
            I => \N__36604\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36601\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36661\,
            I => \N__36596\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__36656\,
            I => \N__36596\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__36651\,
            I => \N__36593\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36648\,
            I => \N__36590\
        );

    \I__7483\ : Span4Mux_s1_h
    port map (
            O => \N__36645\,
            I => \N__36585\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__36640\,
            I => \N__36585\
        );

    \I__7481\ : Span4Mux_h
    port map (
            O => \N__36635\,
            I => \N__36580\
        );

    \I__7480\ : Span4Mux_v
    port map (
            O => \N__36632\,
            I => \N__36580\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36577\
        );

    \I__7478\ : Span4Mux_h
    port map (
            O => \N__36626\,
            I => \N__36574\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36571\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36564\
        );

    \I__7475\ : InMux
    port map (
            O => \N__36621\,
            I => \N__36564\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36564\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__36615\,
            I => \N__36560\
        );

    \I__7472\ : Span4Mux_v
    port map (
            O => \N__36610\,
            I => \N__36557\
        );

    \I__7471\ : Sp12to4
    port map (
            O => \N__36607\,
            I => \N__36554\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__36604\,
            I => \N__36549\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36601\,
            I => \N__36549\
        );

    \I__7468\ : Span4Mux_s2_h
    port map (
            O => \N__36596\,
            I => \N__36546\
        );

    \I__7467\ : Span4Mux_v
    port map (
            O => \N__36593\,
            I => \N__36543\
        );

    \I__7466\ : Span4Mux_s1_v
    port map (
            O => \N__36590\,
            I => \N__36534\
        );

    \I__7465\ : Span4Mux_h
    port map (
            O => \N__36585\,
            I => \N__36534\
        );

    \I__7464\ : Span4Mux_h
    port map (
            O => \N__36580\,
            I => \N__36534\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36534\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__36574\,
            I => \N__36531\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__36571\,
            I => \N__36526\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__36564\,
            I => \N__36526\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36523\
        );

    \I__7458\ : Span4Mux_h
    port map (
            O => \N__36560\,
            I => \N__36520\
        );

    \I__7457\ : Sp12to4
    port map (
            O => \N__36557\,
            I => \N__36515\
        );

    \I__7456\ : Span12Mux_s8_v
    port map (
            O => \N__36554\,
            I => \N__36515\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__36549\,
            I => \N__36508\
        );

    \I__7454\ : Span4Mux_v
    port map (
            O => \N__36546\,
            I => \N__36508\
        );

    \I__7453\ : Span4Mux_s2_h
    port map (
            O => \N__36543\,
            I => \N__36508\
        );

    \I__7452\ : Span4Mux_v
    port map (
            O => \N__36534\,
            I => \N__36505\
        );

    \I__7451\ : Sp12to4
    port map (
            O => \N__36531\,
            I => \N__36500\
        );

    \I__7450\ : Span12Mux_s8_v
    port map (
            O => \N__36526\,
            I => \N__36500\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36523\,
            I => \a_1_repZ0Z2\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__36520\,
            I => \a_1_repZ0Z2\
        );

    \I__7447\ : Odrv12
    port map (
            O => \N__36515\,
            I => \a_1_repZ0Z2\
        );

    \I__7446\ : Odrv4
    port map (
            O => \N__36508\,
            I => \a_1_repZ0Z2\
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__36505\,
            I => \a_1_repZ0Z2\
        );

    \I__7444\ : Odrv12
    port map (
            O => \N__36500\,
            I => \a_1_repZ0Z2\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36481\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36481\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__36481\,
            I => \N__36478\
        );

    \I__7440\ : Span4Mux_s3_h
    port map (
            O => \N__36478\,
            I => \N__36475\
        );

    \I__7439\ : Span4Mux_h
    port map (
            O => \N__36475\,
            I => \N__36472\
        );

    \I__7438\ : Span4Mux_h
    port map (
            O => \N__36472\,
            I => \N__36469\
        );

    \I__7437\ : Sp12to4
    port map (
            O => \N__36469\,
            I => \N__36466\
        );

    \I__7436\ : Odrv12
    port map (
            O => \N__36466\,
            I => \ALU.a10_b_4\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36460\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36460\,
            I => \N__36457\
        );

    \I__7433\ : Span4Mux_s2_v
    port map (
            O => \N__36457\,
            I => \N__36454\
        );

    \I__7432\ : Span4Mux_h
    port map (
            O => \N__36454\,
            I => \N__36451\
        );

    \I__7431\ : Odrv4
    port map (
            O => \N__36451\,
            I => \ALU.r0_12_prm_3_0_s1_c_RNOZ0\
        );

    \I__7430\ : CascadeMux
    port map (
            O => \N__36448\,
            I => \N__36444\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__36447\,
            I => \N__36441\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36444\,
            I => \N__36434\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36434\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36429\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36429\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36426\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__36429\,
            I => \N__36421\
        );

    \I__7422\ : Span4Mux_h
    port map (
            O => \N__36426\,
            I => \N__36421\
        );

    \I__7421\ : Span4Mux_v
    port map (
            O => \N__36421\,
            I => \N__36418\
        );

    \I__7420\ : Odrv4
    port map (
            O => \N__36418\,
            I => \ALU.mult_0\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36412\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36409\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__36409\,
            I => \N__36406\
        );

    \I__7416\ : Sp12to4
    port map (
            O => \N__36406\,
            I => \N__36403\
        );

    \I__7415\ : Odrv12
    port map (
            O => \N__36403\,
            I => \ALU.r0_12_prm_1_0_s1_c_RNOZ0\
        );

    \I__7414\ : CascadeMux
    port map (
            O => \N__36400\,
            I => \N__36396\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36393\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36396\,
            I => \N__36390\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__36393\,
            I => \ALU.un9_addsub_axb_0\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36390\,
            I => \ALU.un9_addsub_axb_0\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36385\,
            I => \bfn_12_3_0_\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36379\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__36379\,
            I => \ALU.r0_12_s1_0_THRU_CO\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36373\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__36373\,
            I => \N__36370\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__36370\,
            I => \ALU.rshift_15_ns_1_0\
        );

    \I__7403\ : CascadeMux
    port map (
            O => \N__36367\,
            I => \N__36364\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36361\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__36361\,
            I => \ALU.r0_12_prm_2_0_s0_c_RNOZ0\
        );

    \I__7400\ : CascadeMux
    port map (
            O => \N__36358\,
            I => \N__36355\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36352\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__36352\,
            I => \ALU.r0_12_prm_1_6_s1_c_RNOZ0\
        );

    \I__7397\ : CascadeMux
    port map (
            O => \N__36349\,
            I => \ALU.rshift_3_ns_1_4_cascade_\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36346\,
            I => \N__36343\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__36343\,
            I => \N__36340\
        );

    \I__7394\ : Span4Mux_s2_v
    port map (
            O => \N__36340\,
            I => \N__36337\
        );

    \I__7393\ : Odrv4
    port map (
            O => \N__36337\,
            I => \ALU.r0_12_prm_7_0_s1_c_RNOZ0\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36331\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__36331\,
            I => \N__36328\
        );

    \I__7390\ : Span4Mux_s1_v
    port map (
            O => \N__36328\,
            I => \N__36325\
        );

    \I__7389\ : Span4Mux_h
    port map (
            O => \N__36325\,
            I => \N__36322\
        );

    \I__7388\ : Span4Mux_h
    port map (
            O => \N__36322\,
            I => \N__36319\
        );

    \I__7387\ : Odrv4
    port map (
            O => \N__36319\,
            I => \ALU.r0_12_prm_6_0_s1_c_RNOZ0\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__36316\,
            I => \N__36313\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36309\
        );

    \I__7384\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36306\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__36309\,
            I => \N__36303\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36298\
        );

    \I__7381\ : Span4Mux_s2_v
    port map (
            O => \N__36303\,
            I => \N__36298\
        );

    \I__7380\ : Span4Mux_h
    port map (
            O => \N__36298\,
            I => \N__36295\
        );

    \I__7379\ : Odrv4
    port map (
            O => \N__36295\,
            I => \ALU.un14_log_0_i_0\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36289\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__36289\,
            I => \ALU.r0_12_prm_5_0_s1_c_RNOZ0\
        );

    \I__7376\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36283\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36283\,
            I => \ALU.r0_12_prm_4_0_s1_c_RNOZ0\
        );

    \I__7374\ : CascadeMux
    port map (
            O => \N__36280\,
            I => \N__36276\
        );

    \I__7373\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36273\
        );

    \I__7372\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36270\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__36273\,
            I => \ALU.N_883_i\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__36270\,
            I => \ALU.N_883_i\
        );

    \I__7369\ : InMux
    port map (
            O => \N__36265\,
            I => \N__36262\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__36262\,
            I => \ALU.r0_12_prm_3_15_s0_sf\
        );

    \I__7367\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36256\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36253\
        );

    \I__7365\ : Span4Mux_h
    port map (
            O => \N__36253\,
            I => \N__36249\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36245\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__36249\,
            I => \N__36242\
        );

    \I__7362\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36239\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36245\,
            I => \N__36236\
        );

    \I__7360\ : Span4Mux_v
    port map (
            O => \N__36242\,
            I => \N__36232\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__36239\,
            I => \N__36229\
        );

    \I__7358\ : Span4Mux_v
    port map (
            O => \N__36236\,
            I => \N__36226\
        );

    \I__7357\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36223\
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__36232\,
            I => \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__36229\,
            I => \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9\
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__36226\,
            I => \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__36223\,
            I => \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9\
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__36214\,
            I => \N__36211\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36208\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36208\,
            I => \N__36205\
        );

    \I__7349\ : Odrv4
    port map (
            O => \N__36205\,
            I => \ALU.r0_12_prm_2_15_s0_c_RNOZ0\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36199\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__36196\
        );

    \I__7346\ : Odrv12
    port map (
            O => \N__36196\,
            I => \ALU.r0_12_prm_1_15_s0_c_RNOZ0\
        );

    \I__7345\ : InMux
    port map (
            O => \N__36193\,
            I => \ALU.r0_12_s0_15\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36187\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__36187\,
            I => \N__36184\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__36184\,
            I => \N__36181\
        );

    \I__7341\ : Sp12to4
    port map (
            O => \N__36181\,
            I => \N__36178\
        );

    \I__7340\ : Odrv12
    port map (
            O => \N__36178\,
            I => \ALU.r0_12_s0_15_THRU_CO\
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__36175\,
            I => \N__36172\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36172\,
            I => \N__36169\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__36169\,
            I => \N__36166\
        );

    \I__7336\ : Span4Mux_h
    port map (
            O => \N__36166\,
            I => \N__36163\
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__36163\,
            I => \ALU.r5_RNIB8HG5Z0Z_12\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36156\
        );

    \I__7333\ : CascadeMux
    port map (
            O => \N__36159\,
            I => \N__36153\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__36156\,
            I => \N__36150\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36147\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__36150\,
            I => \N__36142\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__36147\,
            I => \N__36142\
        );

    \I__7328\ : Span4Mux_h
    port map (
            O => \N__36142\,
            I => \N__36137\
        );

    \I__7327\ : InMux
    port map (
            O => \N__36141\,
            I => \N__36134\
        );

    \I__7326\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36131\
        );

    \I__7325\ : Sp12to4
    port map (
            O => \N__36137\,
            I => \N__36124\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__36134\,
            I => \N__36124\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36131\,
            I => \N__36124\
        );

    \I__7322\ : Span12Mux_v
    port map (
            O => \N__36124\,
            I => \N__36121\
        );

    \I__7321\ : Odrv12
    port map (
            O => \N__36121\,
            I => \ALU.lshift_13\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36118\,
            I => \N__36115\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36112\
        );

    \I__7318\ : Odrv4
    port map (
            O => \N__36112\,
            I => \ALU.r0_12_prm_8_13_s1_c_RNOZ0\
        );

    \I__7317\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36105\
        );

    \I__7316\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36102\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__36105\,
            I => \N__36097\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__36102\,
            I => \N__36094\
        );

    \I__7313\ : InMux
    port map (
            O => \N__36101\,
            I => \N__36091\
        );

    \I__7312\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36088\
        );

    \I__7311\ : Span4Mux_h
    port map (
            O => \N__36097\,
            I => \N__36081\
        );

    \I__7310\ : Span4Mux_v
    port map (
            O => \N__36094\,
            I => \N__36081\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__36091\,
            I => \N__36081\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__36088\,
            I => \N__36078\
        );

    \I__7307\ : Odrv4
    port map (
            O => \N__36081\,
            I => \ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8\
        );

    \I__7306\ : Odrv12
    port map (
            O => \N__36078\,
            I => \ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8\
        );

    \I__7305\ : CascadeMux
    port map (
            O => \N__36073\,
            I => \N__36070\
        );

    \I__7304\ : InMux
    port map (
            O => \N__36070\,
            I => \N__36067\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__36067\,
            I => \ALU.r0_12_prm_1_10_s1_c_RNOZ0\
        );

    \I__7302\ : CascadeMux
    port map (
            O => \N__36064\,
            I => \N__36061\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36061\,
            I => \N__36058\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__36058\,
            I => \N__36055\
        );

    \I__7299\ : Odrv12
    port map (
            O => \N__36055\,
            I => \ALU.r0_12_prm_1_12_s0_c_RNOZ0\
        );

    \I__7298\ : CascadeMux
    port map (
            O => \N__36052\,
            I => \N__36049\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36046\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36043\
        );

    \I__7295\ : Span4Mux_h
    port map (
            O => \N__36043\,
            I => \N__36040\
        );

    \I__7294\ : Odrv4
    port map (
            O => \N__36040\,
            I => \ALU.r0_12_prm_2_14_s0_c_RNOZ0\
        );

    \I__7293\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36034\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36034\,
            I => \ALU.rshift_15\
        );

    \I__7291\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36028\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__36028\,
            I => \N__36024\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36027\,
            I => \N__36021\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__36024\,
            I => \N__36018\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__36015\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__36018\,
            I => \N__36008\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__36015\,
            I => \N__36008\
        );

    \I__7284\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36005\
        );

    \I__7283\ : InMux
    port map (
            O => \N__36013\,
            I => \N__36002\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__36008\,
            I => \ALU.lshift_15\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__36005\,
            I => \ALU.lshift_15\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__36002\,
            I => \ALU.lshift_15\
        );

    \I__7279\ : CascadeMux
    port map (
            O => \N__35995\,
            I => \N__35992\
        );

    \I__7278\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35989\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__35989\,
            I => \ALU.r0_12_prm_8_15_s0_c_RNOZ0\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35983\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__35983\,
            I => \N__35979\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__35982\,
            I => \N__35976\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__35979\,
            I => \N__35973\
        );

    \I__7272\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35970\
        );

    \I__7271\ : Sp12to4
    port map (
            O => \N__35973\,
            I => \N__35965\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__35970\,
            I => \N__35965\
        );

    \I__7269\ : Odrv12
    port map (
            O => \N__35965\,
            I => \ALU.r2_RNI7AQC9_0Z0Z_15\
        );

    \I__7268\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35959\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__35959\,
            I => \N__35956\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__35956\,
            I => \ALU.r0_12_prm_6_15_s0_c_RNOZ0\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__7264\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35946\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35943\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__35946\,
            I => \N__35940\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35943\,
            I => \N__35937\
        );

    \I__7260\ : Span4Mux_v
    port map (
            O => \N__35940\,
            I => \N__35934\
        );

    \I__7259\ : Span4Mux_h
    port map (
            O => \N__35937\,
            I => \N__35931\
        );

    \I__7258\ : Sp12to4
    port map (
            O => \N__35934\,
            I => \N__35928\
        );

    \I__7257\ : Sp12to4
    port map (
            O => \N__35931\,
            I => \N__35923\
        );

    \I__7256\ : Span12Mux_h
    port map (
            O => \N__35928\,
            I => \N__35923\
        );

    \I__7255\ : Odrv12
    port map (
            O => \N__35923\,
            I => \ALU.un14_log_0_i_15\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35917\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__35917\,
            I => \N__35914\
        );

    \I__7252\ : Odrv12
    port map (
            O => \N__35914\,
            I => \ALU.r0_12_prm_5_15_s0_c_RNOZ0\
        );

    \I__7251\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35907\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__35910\,
            I => \N__35904\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__35907\,
            I => \N__35901\
        );

    \I__7248\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35898\
        );

    \I__7247\ : Span4Mux_h
    port map (
            O => \N__35901\,
            I => \N__35895\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__35898\,
            I => \N__35892\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__35895\,
            I => \ALU.r2_RNI7AQC9_1Z0Z_15\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__35892\,
            I => \ALU.r2_RNI7AQC9_1Z0Z_15\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35884\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__35884\,
            I => \ALU.r5_RNI5P1F5Z0Z_15\
        );

    \I__7241\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35878\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35875\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__35875\,
            I => \N__35871\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__35874\,
            I => \N__35868\
        );

    \I__7237\ : Span4Mux_h
    port map (
            O => \N__35871\,
            I => \N__35865\
        );

    \I__7236\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35862\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__35865\,
            I => \ALU.a_i_15\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__35862\,
            I => \ALU.a_i_15\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__35857\,
            I => \N__35854\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35851\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__35851\,
            I => \N__35848\
        );

    \I__7230\ : Odrv12
    port map (
            O => \N__35848\,
            I => \ALU.r0_12_prm_2_10_s0_c_RNOZ0\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__35845\,
            I => \N__35841\
        );

    \I__7228\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35838\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35835\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__35838\,
            I => \N__35828\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__35835\,
            I => \N__35828\
        );

    \I__7224\ : InMux
    port map (
            O => \N__35834\,
            I => \N__35825\
        );

    \I__7223\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35822\
        );

    \I__7222\ : Span12Mux_v
    port map (
            O => \N__35828\,
            I => \N__35819\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__35825\,
            I => \N__35816\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35813\
        );

    \I__7219\ : Odrv12
    port map (
            O => \N__35819\,
            I => \ALU.un2_addsub_cry_10_c_RNIS4T7DZ0\
        );

    \I__7218\ : Odrv4
    port map (
            O => \N__35816\,
            I => \ALU.un2_addsub_cry_10_c_RNIS4T7DZ0\
        );

    \I__7217\ : Odrv4
    port map (
            O => \N__35813\,
            I => \ALU.un2_addsub_cry_10_c_RNIS4T7DZ0\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__35806\,
            I => \N__35803\
        );

    \I__7215\ : InMux
    port map (
            O => \N__35803\,
            I => \N__35800\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__35800\,
            I => \N__35797\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__35797\,
            I => \N__35794\
        );

    \I__7212\ : Span4Mux_h
    port map (
            O => \N__35794\,
            I => \N__35791\
        );

    \I__7211\ : Span4Mux_h
    port map (
            O => \N__35791\,
            I => \N__35788\
        );

    \I__7210\ : Odrv4
    port map (
            O => \N__35788\,
            I => \ALU.r0_12_prm_2_11_s1_c_RNOZ0\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35782\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35782\,
            I => \ALU.r5_RNIAP7U9Z0Z_10\
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__35779\,
            I => \ALU.r5_RNIKU3HJZ0Z_10_cascade_\
        );

    \I__7206\ : CascadeMux
    port map (
            O => \N__35776\,
            I => \ALU.r4_RNIQK1V71Z0Z_5_cascade_\
        );

    \I__7205\ : InMux
    port map (
            O => \N__35773\,
            I => \N__35769\
        );

    \I__7204\ : InMux
    port map (
            O => \N__35772\,
            I => \N__35765\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35769\,
            I => \N__35762\
        );

    \I__7202\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35759\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35752\
        );

    \I__7200\ : Span4Mux_v
    port map (
            O => \N__35762\,
            I => \N__35752\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__35759\,
            I => \N__35752\
        );

    \I__7198\ : Span4Mux_v
    port map (
            O => \N__35752\,
            I => \N__35749\
        );

    \I__7197\ : Span4Mux_h
    port map (
            O => \N__35749\,
            I => \N__35745\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35742\
        );

    \I__7195\ : Span4Mux_h
    port map (
            O => \N__35745\,
            I => \N__35739\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35736\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__35739\,
            I => \ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__35736\,
            I => \ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__35731\,
            I => \N__35728\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35725\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35722\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__35722\,
            I => \N__35719\
        );

    \I__7187\ : Span4Mux_h
    port map (
            O => \N__35719\,
            I => \N__35716\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__35716\,
            I => \ALU.r0_12_prm_1_11_s0_c_RNOZ0\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__35713\,
            I => \N__35710\
        );

    \I__7184\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35707\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__35707\,
            I => \N__35704\
        );

    \I__7182\ : Span4Mux_h
    port map (
            O => \N__35704\,
            I => \N__35701\
        );

    \I__7181\ : Span4Mux_v
    port map (
            O => \N__35701\,
            I => \N__35698\
        );

    \I__7180\ : Odrv4
    port map (
            O => \N__35698\,
            I => \ALU.r0_12_prm_8_13_s0_c_RNOZ0\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__35695\,
            I => \N__35692\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35692\,
            I => \N__35689\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35686\
        );

    \I__7176\ : Span4Mux_h
    port map (
            O => \N__35686\,
            I => \N__35683\
        );

    \I__7175\ : Span4Mux_v
    port map (
            O => \N__35683\,
            I => \N__35680\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__35680\,
            I => \ALU.r0_12_prm_2_12_s0_c_RNOZ0\
        );

    \I__7173\ : CascadeMux
    port map (
            O => \N__35677\,
            I => \N__35674\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35674\,
            I => \N__35671\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__35671\,
            I => \N__35668\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__35668\,
            I => \ALU.r0_12_prm_1_9_s0_c_RNOZ0\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35662\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__35662\,
            I => \N__35659\
        );

    \I__7167\ : Odrv12
    port map (
            O => \N__35659\,
            I => \ALU.lshift_3_ns_1_13\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35653\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35653\,
            I => \N__35650\
        );

    \I__7164\ : Span4Mux_v
    port map (
            O => \N__35650\,
            I => \N__35647\
        );

    \I__7163\ : Span4Mux_h
    port map (
            O => \N__35647\,
            I => \N__35644\
        );

    \I__7162\ : Odrv4
    port map (
            O => \N__35644\,
            I => \ALU.rshift_12\
        );

    \I__7161\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35638\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__35638\,
            I => \N__35633\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35629\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35626\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35623\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35620\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35629\,
            I => \N__35615\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__35626\,
            I => \N__35615\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__35623\,
            I => \ALU.un2_addsub_cry_9_c_RNIS67KDZ0\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35620\,
            I => \ALU.un2_addsub_cry_9_c_RNIS67KDZ0\
        );

    \I__7151\ : Odrv12
    port map (
            O => \N__35615\,
            I => \ALU.un2_addsub_cry_9_c_RNIS67KDZ0\
        );

    \I__7150\ : InMux
    port map (
            O => \N__35608\,
            I => \ALU.un9_addsub_cry_9\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35601\
        );

    \I__7148\ : CascadeMux
    port map (
            O => \N__35604\,
            I => \N__35598\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__35601\,
            I => \N__35595\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35589\
        );

    \I__7145\ : Span4Mux_v
    port map (
            O => \N__35595\,
            I => \N__35585\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35582\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__35593\,
            I => \N__35574\
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__35592\,
            I => \N__35570\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__35589\,
            I => \N__35563\
        );

    \I__7140\ : CascadeMux
    port map (
            O => \N__35588\,
            I => \N__35559\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__35585\,
            I => \N__35554\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35582\,
            I => \N__35554\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35551\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35548\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35541\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35541\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35541\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35534\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35534\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35531\
        );

    \I__7129\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35528\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35521\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35521\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35521\
        );

    \I__7125\ : Span4Mux_v
    port map (
            O => \N__35563\,
            I => \N__35518\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35515\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35512\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__35554\,
            I => \N__35507\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35507\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35502\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__35541\,
            I => \N__35502\
        );

    \I__7118\ : CascadeMux
    port map (
            O => \N__35540\,
            I => \N__35497\
        );

    \I__7117\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35493\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35534\,
            I => \N__35490\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35483\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35528\,
            I => \N__35483\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35521\,
            I => \N__35483\
        );

    \I__7112\ : Span4Mux_h
    port map (
            O => \N__35518\,
            I => \N__35478\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__35515\,
            I => \N__35478\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35473\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__35507\,
            I => \N__35473\
        );

    \I__7108\ : Span12Mux_v
    port map (
            O => \N__35502\,
            I => \N__35470\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35467\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35460\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35460\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35496\,
            I => \N__35460\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__35493\,
            I => \N__35453\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__35490\,
            I => \N__35453\
        );

    \I__7101\ : Span4Mux_v
    port map (
            O => \N__35483\,
            I => \N__35453\
        );

    \I__7100\ : Span4Mux_h
    port map (
            O => \N__35478\,
            I => \N__35450\
        );

    \I__7099\ : Span4Mux_v
    port map (
            O => \N__35473\,
            I => \N__35447\
        );

    \I__7098\ : Odrv12
    port map (
            O => \N__35470\,
            I => \ALU.b_11\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__35467\,
            I => \ALU.b_11\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__35460\,
            I => \ALU.b_11\
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__35453\,
            I => \ALU.b_11\
        );

    \I__7094\ : Odrv4
    port map (
            O => \N__35450\,
            I => \ALU.b_11\
        );

    \I__7093\ : Odrv4
    port map (
            O => \N__35447\,
            I => \ALU.b_11\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35434\,
            I => \ALU.un9_addsub_cry_10\
        );

    \I__7091\ : InMux
    port map (
            O => \N__35431\,
            I => \ALU.un9_addsub_cry_11\
        );

    \I__7090\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35421\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__35427\,
            I => \N__35418\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__35426\,
            I => \N__35415\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \N__35412\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__35424\,
            I => \N__35407\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35421\,
            I => \N__35404\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35393\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35393\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35412\,
            I => \N__35393\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35393\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35393\
        );

    \I__7079\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35389\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__35404\,
            I => \N__35384\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35381\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35378\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__35389\,
            I => \N__35375\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35388\,
            I => \N__35368\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35387\,
            I => \N__35368\
        );

    \I__7072\ : Span4Mux_h
    port map (
            O => \N__35384\,
            I => \N__35361\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__35381\,
            I => \N__35361\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35378\,
            I => \N__35361\
        );

    \I__7069\ : Span4Mux_v
    port map (
            O => \N__35375\,
            I => \N__35358\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35374\,
            I => \N__35355\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35373\,
            I => \N__35352\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35368\,
            I => \N__35349\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__35361\,
            I => \N__35344\
        );

    \I__7064\ : Span4Mux_h
    port map (
            O => \N__35358\,
            I => \N__35341\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35355\,
            I => \N__35338\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__35352\,
            I => \N__35335\
        );

    \I__7061\ : Span4Mux_v
    port map (
            O => \N__35349\,
            I => \N__35332\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35327\
        );

    \I__7059\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35327\
        );

    \I__7058\ : Sp12to4
    port map (
            O => \N__35344\,
            I => \N__35324\
        );

    \I__7057\ : Span4Mux_h
    port map (
            O => \N__35341\,
            I => \N__35321\
        );

    \I__7056\ : Span4Mux_v
    port map (
            O => \N__35338\,
            I => \N__35318\
        );

    \I__7055\ : Span4Mux_s1_h
    port map (
            O => \N__35335\,
            I => \N__35313\
        );

    \I__7054\ : Span4Mux_v
    port map (
            O => \N__35332\,
            I => \N__35313\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__35327\,
            I => \ALU.b_13\
        );

    \I__7052\ : Odrv12
    port map (
            O => \N__35324\,
            I => \ALU.b_13\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__35321\,
            I => \ALU.b_13\
        );

    \I__7050\ : Odrv4
    port map (
            O => \N__35318\,
            I => \ALU.b_13\
        );

    \I__7049\ : Odrv4
    port map (
            O => \N__35313\,
            I => \ALU.b_13\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35297\
        );

    \I__7047\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35291\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35291\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35288\
        );

    \I__7044\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35285\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__35291\,
            I => \N__35282\
        );

    \I__7042\ : Span4Mux_v
    port map (
            O => \N__35288\,
            I => \N__35279\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35285\,
            I => \N__35274\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__35282\,
            I => \N__35274\
        );

    \I__7039\ : Span4Mux_h
    port map (
            O => \N__35279\,
            I => \N__35269\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__35274\,
            I => \N__35269\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__35269\,
            I => \ALU.un9_addsub_cry_12_c_RNISR30AZ0\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35266\,
            I => \ALU.un9_addsub_cry_12\
        );

    \I__7035\ : InMux
    port map (
            O => \N__35263\,
            I => \ALU.un9_addsub_cry_13\
        );

    \I__7034\ : InMux
    port map (
            O => \N__35260\,
            I => \ALU.un9_addsub_cry_14\
        );

    \I__7033\ : CascadeMux
    port map (
            O => \N__35257\,
            I => \N__35254\
        );

    \I__7032\ : InMux
    port map (
            O => \N__35254\,
            I => \N__35251\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35248\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__35248\,
            I => \N__35245\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__35245\,
            I => \N__35242\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__35242\,
            I => \ALU.r0_12_prm_6_10_s0_c_RNOZ0\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__35239\,
            I => \N__35236\
        );

    \I__7026\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35233\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35233\,
            I => \N__35230\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__35230\,
            I => \N__35227\
        );

    \I__7023\ : Span4Mux_v
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__7022\ : Odrv4
    port map (
            O => \N__35224\,
            I => \ALU.r4_RNI90J9EZ0Z_1\
        );

    \I__7021\ : InMux
    port map (
            O => \N__35221\,
            I => \ALU.un9_addsub_cry_0\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35215\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__35215\,
            I => \ALU.r4_RNI468UDZ0Z_2\
        );

    \I__7018\ : InMux
    port map (
            O => \N__35212\,
            I => \ALU.un9_addsub_cry_1\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__35209\,
            I => \N__35206\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35203\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35200\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__35200\,
            I => \N__35197\
        );

    \I__7013\ : Odrv4
    port map (
            O => \N__35197\,
            I => \ALU.r4_RNIUU8UDZ0Z_3\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35194\,
            I => \ALU.un9_addsub_cry_2\
        );

    \I__7011\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35188\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__35188\,
            I => \N__35185\
        );

    \I__7009\ : Odrv4
    port map (
            O => \N__35185\,
            I => \ALU.r4_RNIQK1EDZ0Z_4\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35182\,
            I => \ALU.un9_addsub_cry_3\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35179\,
            I => \ALU.un9_addsub_cry_4\
        );

    \I__7006\ : InMux
    port map (
            O => \N__35176\,
            I => \ALU.un9_addsub_cry_5\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35173\,
            I => \ALU.un9_addsub_cry_6\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35170\,
            I => \bfn_11_9_0_\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35167\,
            I => \ALU.un9_addsub_cry_8\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__35164\,
            I => \ALU.r5_RNI9S2TIZ0Z_11_cascade_\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__35161\,
            I => \ALU.lshift_15_ns_1_13_cascade_\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35158\,
            I => \N__35155\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__35155\,
            I => \N__35152\
        );

    \I__6998\ : Odrv4
    port map (
            O => \N__35152\,
            I => \ALU.un9_addsub_axb_2\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__35149\,
            I => \N__35146\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35142\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35139\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35142\,
            I => \N__35136\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35133\
        );

    \I__6992\ : Span4Mux_h
    port map (
            O => \N__35136\,
            I => \N__35130\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__35133\,
            I => \N__35125\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__35130\,
            I => \N__35125\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__35125\,
            I => \N__35122\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__35122\,
            I => \N__35119\
        );

    \I__6987\ : Odrv4
    port map (
            O => \N__35119\,
            I => \ALU.un14_log_0_i_11\
        );

    \I__6986\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35110\
        );

    \I__6985\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35110\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__35110\,
            I => \N__35107\
        );

    \I__6983\ : Span4Mux_h
    port map (
            O => \N__35107\,
            I => \N__35104\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__35104\,
            I => \ALU.a6_b_0\
        );

    \I__6981\ : CascadeMux
    port map (
            O => \N__35101\,
            I => \ALU.lshift_3_ns_1_8_cascade_\
        );

    \I__6980\ : CascadeMux
    port map (
            O => \N__35098\,
            I => \ALU.r4_RNILIPV9Z0Z_6_cascade_\
        );

    \I__6979\ : CascadeMux
    port map (
            O => \N__35095\,
            I => \ALU.r4_RNI1G9PKZ0Z_6_cascade_\
        );

    \I__6978\ : CascadeMux
    port map (
            O => \N__35092\,
            I => \N__35089\
        );

    \I__6977\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35086\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__35086\,
            I => \N__35083\
        );

    \I__6975\ : Span4Mux_h
    port map (
            O => \N__35083\,
            I => \N__35079\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35076\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__35079\,
            I => \N__35073\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35070\
        );

    \I__6971\ : Span4Mux_v
    port map (
            O => \N__35073\,
            I => \N__35066\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__35070\,
            I => \N__35063\
        );

    \I__6969\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35060\
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__35066\,
            I => r0_1
        );

    \I__6967\ : Odrv4
    port map (
            O => \N__35063\,
            I => r0_1
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__35060\,
            I => r0_1
        );

    \I__6965\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35050\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35046\
        );

    \I__6963\ : InMux
    port map (
            O => \N__35049\,
            I => \N__35043\
        );

    \I__6962\ : Span4Mux_h
    port map (
            O => \N__35046\,
            I => \N__35037\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__35043\,
            I => \N__35037\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35034\
        );

    \I__6959\ : Span4Mux_h
    port map (
            O => \N__35037\,
            I => \N__35031\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__35034\,
            I => r0_3
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__35031\,
            I => r0_3
        );

    \I__6956\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35022\
        );

    \I__6955\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35019\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__35022\,
            I => \N__35013\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__35019\,
            I => \N__35013\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35010\
        );

    \I__6951\ : Span4Mux_v
    port map (
            O => \N__35013\,
            I => \N__35004\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35010\,
            I => \N__35004\
        );

    \I__6949\ : InMux
    port map (
            O => \N__35009\,
            I => \N__35001\
        );

    \I__6948\ : Span4Mux_v
    port map (
            O => \N__35004\,
            I => \N__34997\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34994\
        );

    \I__6946\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34991\
        );

    \I__6945\ : Span4Mux_v
    port map (
            O => \N__34997\,
            I => \N__34988\
        );

    \I__6944\ : Sp12to4
    port map (
            O => \N__34994\,
            I => \N__34983\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__34991\,
            I => \N__34980\
        );

    \I__6942\ : Span4Mux_h
    port map (
            O => \N__34988\,
            I => \N__34977\
        );

    \I__6941\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34974\
        );

    \I__6940\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34971\
        );

    \I__6939\ : Span12Mux_v
    port map (
            O => \N__34983\,
            I => \N__34967\
        );

    \I__6938\ : Span12Mux_s10_h
    port map (
            O => \N__34980\,
            I => \N__34964\
        );

    \I__6937\ : Span4Mux_h
    port map (
            O => \N__34977\,
            I => \N__34959\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34974\,
            I => \N__34959\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__34971\,
            I => \N__34956\
        );

    \I__6934\ : InMux
    port map (
            O => \N__34970\,
            I => \N__34953\
        );

    \I__6933\ : Odrv12
    port map (
            O => \N__34967\,
            I => \ALU.r0_12_0\
        );

    \I__6932\ : Odrv12
    port map (
            O => \N__34964\,
            I => \ALU.r0_12_0\
        );

    \I__6931\ : Odrv4
    port map (
            O => \N__34959\,
            I => \ALU.r0_12_0\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__34956\,
            I => \ALU.r0_12_0\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__34953\,
            I => \ALU.r0_12_0\
        );

    \I__6928\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34936\
        );

    \I__6927\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34936\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__34936\,
            I => \N__34933\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__34933\,
            I => \N__34929\
        );

    \I__6924\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34926\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__34929\,
            I => r0_0
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__34926\,
            I => r0_0
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__34921\,
            I => \N__34918\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34918\,
            I => \N__34915\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__34915\,
            I => \ALU.r0_12_prm_5_0_s0_c_RNOZ0\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__34912\,
            I => \N__34909\
        );

    \I__6917\ : InMux
    port map (
            O => \N__34909\,
            I => \N__34906\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__34906\,
            I => \N__34903\
        );

    \I__6915\ : Span4Mux_s2_v
    port map (
            O => \N__34903\,
            I => \N__34900\
        );

    \I__6914\ : Span4Mux_h
    port map (
            O => \N__34900\,
            I => \N__34897\
        );

    \I__6913\ : Odrv4
    port map (
            O => \N__34897\,
            I => \ALU.r2_RNIKG5N5Z0Z_0\
        );

    \I__6912\ : CascadeMux
    port map (
            O => \N__34894\,
            I => \N__34891\
        );

    \I__6911\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34888\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__34888\,
            I => \N__34885\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__34885\,
            I => \ALU.r0_12_prm_3_0_s0_c_RNOZ0\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__34882\,
            I => \N__34879\
        );

    \I__6907\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34876\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__34876\,
            I => \N__34873\
        );

    \I__6905\ : Span4Mux_h
    port map (
            O => \N__34873\,
            I => \N__34870\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__34870\,
            I => \ALU.r0_12_prm_1_0_s0_c_RNOZ0\
        );

    \I__6903\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34864\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__34864\,
            I => \N__34861\
        );

    \I__6901\ : Odrv4
    port map (
            O => \N__34861\,
            I => \ALU.rshift_0\
        );

    \I__6900\ : InMux
    port map (
            O => \N__34858\,
            I => \bfn_11_4_0_\
        );

    \I__6899\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34848\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34848\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__34853\,
            I => \N__34845\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34848\,
            I => \N__34842\
        );

    \I__6895\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34839\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__34842\,
            I => \N__34836\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34833\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__34836\,
            I => \N__34828\
        );

    \I__6891\ : Span4Mux_v
    port map (
            O => \N__34833\,
            I => \N__34828\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__34828\,
            I => r1_0
        );

    \I__6889\ : InMux
    port map (
            O => \N__34825\,
            I => \ALU.r0_12_s1_6\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__34822\,
            I => \ALU.lshift_6_cascade_\
        );

    \I__6887\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34816\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__34816\,
            I => \ALU.r0_12_prm_8_6_s1_c_RNOZ0\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__34813\,
            I => \N__34810\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34807\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34807\,
            I => \N__34804\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__34804\,
            I => \ALU.r0_12_prm_7_0_s0_c_RNOZ0\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__34801\,
            I => \N__34798\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34795\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34795\,
            I => \N__34792\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__34792\,
            I => \ALU.r0_12_prm_6_0_s0_c_RNOZ0\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__34789\,
            I => \N__34786\
        );

    \I__6876\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34783\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__34783\,
            I => \ALU.r0_12_prm_7_6_s1_c_RNOZ0\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34777\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__34777\,
            I => \ALU.r0_12_prm_6_6_s1_c_RNOZ0\
        );

    \I__6872\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34771\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34768\
        );

    \I__6870\ : Odrv4
    port map (
            O => \N__34768\,
            I => \ALU.r0_12_prm_5_6_s1_c_RNOZ0\
        );

    \I__6869\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34762\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34759\
        );

    \I__6867\ : Span4Mux_h
    port map (
            O => \N__34759\,
            I => \N__34756\
        );

    \I__6866\ : Odrv4
    port map (
            O => \N__34756\,
            I => \ALU.r0_12_prm_4_6_s1_c_RNOZ0\
        );

    \I__6865\ : CascadeMux
    port map (
            O => \N__34753\,
            I => \N__34750\
        );

    \I__6864\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34747\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__34747\,
            I => \ALU.r0_12_prm_2_6_s1_c_RNOZ0\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34744\,
            I => \N__34741\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34741\,
            I => \ALU.r0_12_prm_6_10_s1_c_RNOZ0\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__34738\,
            I => \N__34734\
        );

    \I__6859\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34731\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34728\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__34731\,
            I => \N__34725\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34728\,
            I => \N__34722\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__34725\,
            I => \N__34719\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__34722\,
            I => \N__34716\
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__34719\,
            I => \ALU.un14_log_0_i_10\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__34716\,
            I => \ALU.un14_log_0_i_10\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34708\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__34708\,
            I => \ALU.r0_12_prm_5_10_s1_c_RNOZ0\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__34705\,
            I => \N__34702\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34699\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34699\,
            I => \N__34695\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34692\
        );

    \I__6845\ : Span4Mux_h
    port map (
            O => \N__34695\,
            I => \N__34689\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34684\
        );

    \I__6843\ : Span4Mux_v
    port map (
            O => \N__34689\,
            I => \N__34684\
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__34684\,
            I => \ALU.r5_RNIUF9K8_1Z0Z_10\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34678\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34678\,
            I => \ALU.r0_12_prm_4_10_s1_c_RNOZ0\
        );

    \I__6839\ : CascadeMux
    port map (
            O => \N__34675\,
            I => \N__34672\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34669\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__34669\,
            I => \N__34666\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__34666\,
            I => \N__34662\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34665\,
            I => \N__34659\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__34662\,
            I => \N__34656\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__34659\,
            I => \ALU.a_i_10\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__34656\,
            I => \ALU.a_i_10\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__34651\,
            I => \N__34648\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34648\,
            I => \N__34645\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34645\,
            I => \ALU.r0_12_prm_2_10_s1_c_RNOZ0\
        );

    \I__6828\ : InMux
    port map (
            O => \N__34642\,
            I => \ALU.r0_12_s1_10\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34636\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34633\
        );

    \I__6825\ : Span4Mux_h
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__6824\ : Span4Mux_v
    port map (
            O => \N__34630\,
            I => \N__34627\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__34627\,
            I => \ALU.r0_12_s1_10_THRU_CO\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34618\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34615\
        );

    \I__6819\ : Odrv12
    port map (
            O => \N__34615\,
            I => \ALU.r0_12_prm_1_13_s0_c_RNOZ0\
        );

    \I__6818\ : CascadeMux
    port map (
            O => \N__34612\,
            I => \N__34609\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34606\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34603\
        );

    \I__6815\ : Span4Mux_h
    port map (
            O => \N__34603\,
            I => \N__34600\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__34600\,
            I => \ALU.r5_RNI27VE5Z0Z_10\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34593\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__34596\,
            I => \N__34590\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__34593\,
            I => \N__34586\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34583\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34580\
        );

    \I__6808\ : Span4Mux_v
    port map (
            O => \N__34586\,
            I => \N__34576\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34583\,
            I => \N__34571\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34580\,
            I => \N__34571\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34579\,
            I => \N__34568\
        );

    \I__6804\ : Span4Mux_h
    port map (
            O => \N__34576\,
            I => \N__34563\
        );

    \I__6803\ : Span4Mux_v
    port map (
            O => \N__34571\,
            I => \N__34563\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__34568\,
            I => \N__34560\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__34563\,
            I => \ALU.un2_addsub_cry_12_c_RNI74A7EZ0\
        );

    \I__6800\ : Odrv12
    port map (
            O => \N__34560\,
            I => \ALU.un2_addsub_cry_12_c_RNI74A7EZ0\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34552\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34552\,
            I => \ALU.r0_12_prm_2_13_s1_c_RNOZ0\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34546\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__34546\,
            I => \N__34543\
        );

    \I__6795\ : Span4Mux_h
    port map (
            O => \N__34543\,
            I => \N__34540\
        );

    \I__6794\ : Span4Mux_h
    port map (
            O => \N__34540\,
            I => \N__34537\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__34537\,
            I => \ALU.rshift_11\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34531\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34531\,
            I => \N__34528\
        );

    \I__6790\ : Span12Mux_v
    port map (
            O => \N__34528\,
            I => \N__34525\
        );

    \I__6789\ : Odrv12
    port map (
            O => \N__34525\,
            I => \ALU.r0_12_prm_8_10_s1_c_RNOZ0Z_1\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34519\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34519\,
            I => \N__34516\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__34516\,
            I => \ALU.r0_12_prm_7_10_s1_c_RNOZ0\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34509\
        );

    \I__6784\ : CascadeMux
    port map (
            O => \N__34512\,
            I => \N__34506\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__34509\,
            I => \N__34503\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34500\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__34503\,
            I => \N__34497\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34500\,
            I => \N__34494\
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__34497\,
            I => \ALU.r5_RNIUF9K8_0Z0Z_10\
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__34494\,
            I => \ALU.r5_RNIUF9K8_0Z0Z_10\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34489\,
            I => \N__34486\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__34486\,
            I => \N__34483\
        );

    \I__6775\ : Odrv12
    port map (
            O => \N__34483\,
            I => \ALU.N_884_i\
        );

    \I__6774\ : CascadeMux
    port map (
            O => \N__34480\,
            I => \N__34477\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34474\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__34474\,
            I => \N__34471\
        );

    \I__6771\ : Span4Mux_v
    port map (
            O => \N__34471\,
            I => \N__34468\
        );

    \I__6770\ : Odrv4
    port map (
            O => \N__34468\,
            I => \ALU.r0_12_prm_8_12_s0_c_RNOZ0\
        );

    \I__6769\ : CascadeMux
    port map (
            O => \N__34465\,
            I => \ALU.lshift_3_ns_1_3_cascade_\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34458\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34455\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__34458\,
            I => \N__34450\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__34455\,
            I => \N__34450\
        );

    \I__6764\ : Odrv12
    port map (
            O => \N__34450\,
            I => \ALU.r4_RNI1RK3KZ0Z_9\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__34447\,
            I => \ALU.r4_RNIOK1781Z0Z_9_cascade_\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34440\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34443\,
            I => \N__34437\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34440\,
            I => \N__34434\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__34437\,
            I => \N__34431\
        );

    \I__6758\ : Span4Mux_h
    port map (
            O => \N__34434\,
            I => \N__34428\
        );

    \I__6757\ : Span4Mux_h
    port map (
            O => \N__34431\,
            I => \N__34425\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__34428\,
            I => \N__34418\
        );

    \I__6755\ : Span4Mux_h
    port map (
            O => \N__34425\,
            I => \N__34418\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34415\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34412\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__34418\,
            I => \ALU.lshift_11\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34415\,
            I => \ALU.lshift_11\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__34412\,
            I => \ALU.lshift_11\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34402\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34402\,
            I => \N__34398\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34395\
        );

    \I__6746\ : Span4Mux_h
    port map (
            O => \N__34398\,
            I => \N__34392\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34395\,
            I => \N__34388\
        );

    \I__6744\ : Span4Mux_v
    port map (
            O => \N__34392\,
            I => \N__34385\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34391\,
            I => \N__34382\
        );

    \I__6742\ : Span12Mux_s10_v
    port map (
            O => \N__34388\,
            I => \N__34379\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__34385\,
            I => \N__34374\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34374\
        );

    \I__6739\ : Odrv12
    port map (
            O => \N__34379\,
            I => r4_9
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__34374\,
            I => r4_9
        );

    \I__6737\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34365\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34362\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__34365\,
            I => \N__34358\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__34362\,
            I => \N__34355\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34361\,
            I => \N__34352\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__34358\,
            I => \N__34349\
        );

    \I__6731\ : Span4Mux_h
    port map (
            O => \N__34355\,
            I => \N__34346\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34343\
        );

    \I__6729\ : Span4Mux_h
    port map (
            O => \N__34349\,
            I => \N__34338\
        );

    \I__6728\ : Span4Mux_v
    port map (
            O => \N__34346\,
            I => \N__34338\
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__34343\,
            I => r4_1
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__34338\,
            I => r4_1
        );

    \I__6725\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34330\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34326\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34322\
        );

    \I__6722\ : Span4Mux_v
    port map (
            O => \N__34326\,
            I => \N__34319\
        );

    \I__6721\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34316\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34313\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__34319\,
            I => \N__34310\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34305\
        );

    \I__6717\ : Span4Mux_h
    port map (
            O => \N__34313\,
            I => \N__34305\
        );

    \I__6716\ : Odrv4
    port map (
            O => \N__34310\,
            I => r4_2
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__34305\,
            I => r4_2
        );

    \I__6714\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34297\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34297\,
            I => \N__34294\
        );

    \I__6712\ : Span4Mux_v
    port map (
            O => \N__34294\,
            I => \N__34291\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__34291\,
            I => \N__34286\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34283\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34280\
        );

    \I__6708\ : Span4Mux_h
    port map (
            O => \N__34286\,
            I => \N__34277\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__34283\,
            I => \N__34274\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34271\
        );

    \I__6705\ : Span4Mux_h
    port map (
            O => \N__34277\,
            I => \N__34268\
        );

    \I__6704\ : Span4Mux_h
    port map (
            O => \N__34274\,
            I => \N__34263\
        );

    \I__6703\ : Span4Mux_v
    port map (
            O => \N__34271\,
            I => \N__34263\
        );

    \I__6702\ : Odrv4
    port map (
            O => \N__34268\,
            I => r4_4
        );

    \I__6701\ : Odrv4
    port map (
            O => \N__34263\,
            I => r4_4
        );

    \I__6700\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34255\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34252\
        );

    \I__6698\ : Span4Mux_h
    port map (
            O => \N__34252\,
            I => \N__34249\
        );

    \I__6697\ : Span4Mux_v
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__6696\ : Span4Mux_h
    port map (
            O => \N__34246\,
            I => \N__34243\
        );

    \I__6695\ : Span4Mux_h
    port map (
            O => \N__34243\,
            I => \N__34240\
        );

    \I__6694\ : Odrv4
    port map (
            O => \N__34240\,
            I => \ALU.r5_RNIVF7TIZ0Z_13\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__34237\,
            I => \ALU.lshift_15_ns_1_15_cascade_\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34231\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__34231\,
            I => \N__34228\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__34228\,
            I => \N__34225\
        );

    \I__6689\ : Span4Mux_h
    port map (
            O => \N__34225\,
            I => \N__34222\
        );

    \I__6688\ : Span4Mux_h
    port map (
            O => \N__34222\,
            I => \N__34219\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__34219\,
            I => \ALU.r0_12_prm_8_11_s1_c_RNOZ0Z_1\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34213\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34213\,
            I => \N__34210\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__34210\,
            I => \N__34207\
        );

    \I__6683\ : Span4Mux_h
    port map (
            O => \N__34207\,
            I => \N__34204\
        );

    \I__6682\ : Odrv4
    port map (
            O => \N__34204\,
            I => \ALU.r0_12_prm_2_11_s0_c_RNOZ0\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__34201\,
            I => \N__34198\
        );

    \I__6680\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34195\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34192\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__34192\,
            I => \ALU.r0_12_prm_1_10_s0_c_RNOZ0\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__34189\,
            I => \N__34186\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__6674\ : Span4Mux_h
    port map (
            O => \N__34180\,
            I => \N__34177\
        );

    \I__6673\ : Span4Mux_h
    port map (
            O => \N__34177\,
            I => \N__34174\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__34174\,
            I => \ALU.r5_RNIUF9K8_2Z0Z_10\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34171\,
            I => \ALU.un2_addsub_cry_9\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34162\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__34162\,
            I => \N__34159\
        );

    \I__6667\ : Span4Mux_v
    port map (
            O => \N__34159\,
            I => \N__34156\
        );

    \I__6666\ : Span4Mux_h
    port map (
            O => \N__34156\,
            I => \N__34153\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__34153\,
            I => \N__34150\
        );

    \I__6664\ : Odrv4
    port map (
            O => \N__34150\,
            I => \ALU.r5_RNIE0AK8_2Z0Z_11\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34147\,
            I => \ALU.un2_addsub_cry_10\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__34144\,
            I => \N__34141\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34138\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34135\
        );

    \I__6659\ : Odrv12
    port map (
            O => \N__34135\,
            I => \ALU.r5_RNISP2L9_2Z0Z_12\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34132\,
            I => \ALU.un2_addsub_cry_11\
        );

    \I__6657\ : CascadeMux
    port map (
            O => \N__34129\,
            I => \N__34126\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34126\,
            I => \N__34123\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34123\,
            I => \N__34120\
        );

    \I__6654\ : Span4Mux_h
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__34117\,
            I => \N__34114\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__34114\,
            I => \ALU.r5_RNID2JJ9_2Z0Z_13\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34111\,
            I => \ALU.un2_addsub_cry_12\
        );

    \I__6650\ : CascadeMux
    port map (
            O => \N__34108\,
            I => \N__34105\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34102\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__34099\
        );

    \I__6647\ : Odrv12
    port map (
            O => \N__34099\,
            I => \ALU.r2_RNINPPC9_2Z0Z_14\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34096\,
            I => \ALU.un2_addsub_cry_13\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34093\,
            I => \ALU.un2_addsub_cry_14\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34084\
        );

    \I__6643\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34084\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__34084\,
            I => \N__34080\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34077\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__34080\,
            I => \N__34072\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34077\,
            I => \N__34072\
        );

    \I__6638\ : Odrv4
    port map (
            O => \N__34072\,
            I => r4_7
        );

    \I__6637\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34066\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__34066\,
            I => \N__34062\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34059\
        );

    \I__6634\ : Span4Mux_s2_v
    port map (
            O => \N__34062\,
            I => \N__34056\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__34059\,
            I => \N__34052\
        );

    \I__6632\ : Span4Mux_h
    port map (
            O => \N__34056\,
            I => \N__34049\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34055\,
            I => \N__34046\
        );

    \I__6630\ : Span4Mux_h
    port map (
            O => \N__34052\,
            I => \N__34043\
        );

    \I__6629\ : Span4Mux_v
    port map (
            O => \N__34049\,
            I => \N__34038\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__34038\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__34043\,
            I => r4_8
        );

    \I__6626\ : Odrv4
    port map (
            O => \N__34038\,
            I => r4_8
        );

    \I__6625\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34028\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34023\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34019\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__34028\,
            I => \N__34016\
        );

    \I__6621\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34011\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34008\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__34005\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34022\,
            I => \N__34002\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34019\,
            I => \N__33997\
        );

    \I__6616\ : Span4Mux_v
    port map (
            O => \N__34016\,
            I => \N__33997\
        );

    \I__6615\ : InMux
    port map (
            O => \N__34015\,
            I => \N__33994\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34014\,
            I => \N__33991\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__34011\,
            I => \N__33988\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__33983\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__34005\,
            I => \N__33983\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__34002\,
            I => \N__33978\
        );

    \I__6609\ : Span4Mux_h
    port map (
            O => \N__33997\,
            I => \N__33978\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__33994\,
            I => \N__33969\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__33991\,
            I => \N__33969\
        );

    \I__6606\ : Span4Mux_v
    port map (
            O => \N__33988\,
            I => \N__33969\
        );

    \I__6605\ : Span4Mux_h
    port map (
            O => \N__33983\,
            I => \N__33969\
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__33978\,
            I => \ALU.r0_12_9\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__33969\,
            I => \ALU.r0_12_9\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33964\,
            I => \ALU.un2_addsub_cry_0\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33961\,
            I => \N__33958\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33958\,
            I => \N__33955\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__33955\,
            I => \N__33952\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__33952\,
            I => \ALU.r4_RNIUM9JCZ0Z_2\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__33949\,
            I => \N__33946\
        );

    \I__6596\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33943\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__33943\,
            I => \N__33940\
        );

    \I__6594\ : Span4Mux_v
    port map (
            O => \N__33940\,
            I => \N__33937\
        );

    \I__6593\ : Span4Mux_v
    port map (
            O => \N__33937\,
            I => \N__33933\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33930\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__33933\,
            I => \ALU.b_i_2\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__33930\,
            I => \ALU.b_i_2\
        );

    \I__6589\ : InMux
    port map (
            O => \N__33925\,
            I => \ALU.un2_addsub_cry_1\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33919\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__33919\,
            I => \N__33916\
        );

    \I__6586\ : Sp12to4
    port map (
            O => \N__33916\,
            I => \N__33913\
        );

    \I__6585\ : Odrv12
    port map (
            O => \N__33913\,
            I => \ALU.r4_RNINFAJCZ0Z_3\
        );

    \I__6584\ : CascadeMux
    port map (
            O => \N__33910\,
            I => \N__33907\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33904\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33901\
        );

    \I__6581\ : Span12Mux_h
    port map (
            O => \N__33901\,
            I => \N__33898\
        );

    \I__6580\ : Odrv12
    port map (
            O => \N__33898\,
            I => \ALU.b_i_3\
        );

    \I__6579\ : InMux
    port map (
            O => \N__33895\,
            I => \ALU.un2_addsub_cry_2\
        );

    \I__6578\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33889\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33886\
        );

    \I__6576\ : Odrv12
    port map (
            O => \N__33886\,
            I => \ALU.r4_RNI20C8CZ0Z_4\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__33883\,
            I => \N__33879\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33876\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33873\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__33876\,
            I => \N__33870\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__33873\,
            I => \N__33867\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__33870\,
            I => \N__33864\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__33867\,
            I => \N__33859\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__33864\,
            I => \N__33859\
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__33859\,
            I => \ALU.b_i_4\
        );

    \I__6566\ : InMux
    port map (
            O => \N__33856\,
            I => \ALU.un2_addsub_cry_3\
        );

    \I__6565\ : CascadeMux
    port map (
            O => \N__33853\,
            I => \N__33850\
        );

    \I__6564\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33847\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33844\
        );

    \I__6562\ : Span4Mux_v
    port map (
            O => \N__33844\,
            I => \N__33841\
        );

    \I__6561\ : Sp12to4
    port map (
            O => \N__33841\,
            I => \N__33838\
        );

    \I__6560\ : Odrv12
    port map (
            O => \N__33838\,
            I => \ALU.r4_RNI8B628_1Z0Z_5\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33835\,
            I => \ALU.un2_addsub_cry_4\
        );

    \I__6558\ : CascadeMux
    port map (
            O => \N__33832\,
            I => \N__33829\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33826\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__33826\,
            I => \N__33823\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__33823\,
            I => \N__33820\
        );

    \I__6554\ : Span4Mux_h
    port map (
            O => \N__33820\,
            I => \N__33817\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__33817\,
            I => \N__33814\
        );

    \I__6552\ : Span4Mux_s3_v
    port map (
            O => \N__33814\,
            I => \N__33811\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__33811\,
            I => \ALU.r4_RNI2BKQ8_1Z0Z_6\
        );

    \I__6550\ : InMux
    port map (
            O => \N__33808\,
            I => \ALU.un2_addsub_cry_5\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33805\,
            I => \ALU.un2_addsub_cry_6\
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__33802\,
            I => \N__33799\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33796\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__33796\,
            I => \N__33793\
        );

    \I__6545\ : Odrv12
    port map (
            O => \N__33793\,
            I => \ALU.r4_RNIKUMQ8_1Z0Z_8\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33790\,
            I => \bfn_10_10_0_\
        );

    \I__6543\ : InMux
    port map (
            O => \N__33787\,
            I => \ALU.un2_addsub_cry_8\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33780\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33777\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33774\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33771\
        );

    \I__6538\ : Span4Mux_v
    port map (
            O => \N__33774\,
            I => \N__33767\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__33771\,
            I => \N__33764\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33761\
        );

    \I__6535\ : Span4Mux_h
    port map (
            O => \N__33767\,
            I => \N__33758\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__33764\,
            I => \N__33753\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__33761\,
            I => \N__33753\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__33758\,
            I => \N__33748\
        );

    \I__6531\ : Span4Mux_h
    port map (
            O => \N__33753\,
            I => \N__33748\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__33748\,
            I => r5_6
        );

    \I__6529\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33739\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33739\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__33739\,
            I => \N__33735\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33732\
        );

    \I__6525\ : Odrv4
    port map (
            O => \N__33735\,
            I => r5_7
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__33732\,
            I => r5_7
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__33727\,
            I => \N__33724\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33721\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__6520\ : Span4Mux_s2_v
    port map (
            O => \N__33718\,
            I => \N__33713\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33710\
        );

    \I__6518\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33707\
        );

    \I__6517\ : Span4Mux_h
    port map (
            O => \N__33713\,
            I => \N__33704\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33710\,
            I => \N__33699\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__33707\,
            I => \N__33699\
        );

    \I__6514\ : Span4Mux_v
    port map (
            O => \N__33704\,
            I => \N__33696\
        );

    \I__6513\ : Odrv12
    port map (
            O => \N__33699\,
            I => r5_8
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__33696\,
            I => r5_8
        );

    \I__6511\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33688\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33688\,
            I => \N__33684\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33681\
        );

    \I__6508\ : Span4Mux_h
    port map (
            O => \N__33684\,
            I => \N__33677\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33681\,
            I => \N__33674\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33671\
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__33677\,
            I => r5_9
        );

    \I__6504\ : Odrv12
    port map (
            O => \N__33674\,
            I => r5_9
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__33671\,
            I => r5_9
        );

    \I__6502\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33660\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33657\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__33660\,
            I => \N__33654\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__33657\,
            I => \N__33650\
        );

    \I__6498\ : Span4Mux_v
    port map (
            O => \N__33654\,
            I => \N__33647\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33644\
        );

    \I__6496\ : Span4Mux_h
    port map (
            O => \N__33650\,
            I => \N__33641\
        );

    \I__6495\ : Odrv4
    port map (
            O => \N__33647\,
            I => r5_1
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33644\,
            I => r5_1
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__33641\,
            I => r5_1
        );

    \I__6492\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33631\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33628\
        );

    \I__6490\ : Span4Mux_v
    port map (
            O => \N__33628\,
            I => \N__33623\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33620\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33617\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33623\,
            I => r5_2
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33620\,
            I => r5_2
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33617\,
            I => r5_2
        );

    \I__6484\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33604\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__33604\,
            I => \N__33600\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__33603\,
            I => \N__33597\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__33600\,
            I => \N__33594\
        );

    \I__6479\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33591\
        );

    \I__6478\ : Span4Mux_v
    port map (
            O => \N__33594\,
            I => \N__33586\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33591\,
            I => \N__33586\
        );

    \I__6476\ : Span4Mux_h
    port map (
            O => \N__33586\,
            I => \N__33582\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33579\
        );

    \I__6474\ : Odrv4
    port map (
            O => \N__33582\,
            I => r5_3
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__33579\,
            I => r5_3
        );

    \I__6472\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33571\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33571\,
            I => \N__33568\
        );

    \I__6470\ : Span4Mux_v
    port map (
            O => \N__33568\,
            I => \N__33565\
        );

    \I__6469\ : Span4Mux_h
    port map (
            O => \N__33565\,
            I => \N__33562\
        );

    \I__6468\ : Span4Mux_h
    port map (
            O => \N__33562\,
            I => \N__33557\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33554\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33551\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__33557\,
            I => r5_4
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__33554\,
            I => r5_4
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__33551\,
            I => r5_4
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__33544\,
            I => \N__33541\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33538\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__33538\,
            I => \N__33535\
        );

    \I__6459\ : Span4Mux_v
    port map (
            O => \N__33535\,
            I => \N__33532\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__33532\,
            I => \N__33529\
        );

    \I__6457\ : Span4Mux_h
    port map (
            O => \N__33529\,
            I => \N__33526\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__33526\,
            I => \ALU.r4_RNIUES39Z0Z_1\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33520\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__33520\,
            I => \N__33517\
        );

    \I__6453\ : Span4Mux_h
    port map (
            O => \N__33517\,
            I => \N__33514\
        );

    \I__6452\ : Odrv4
    port map (
            O => \N__33514\,
            I => \ALU.b_3_ns_1_0\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__33508\,
            I => \N__33504\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33501\
        );

    \I__6448\ : Span4Mux_h
    port map (
            O => \N__33504\,
            I => \N__33498\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__33501\,
            I => \N__33494\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__33498\,
            I => \N__33491\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33488\
        );

    \I__6444\ : Span4Mux_h
    port map (
            O => \N__33494\,
            I => \N__33485\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__33491\,
            I => r0_4
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__33488\,
            I => r0_4
        );

    \I__6441\ : Odrv4
    port map (
            O => \N__33485\,
            I => r0_4
        );

    \I__6440\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33475\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__33475\,
            I => \N__33472\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__33472\,
            I => \N__33469\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__33469\,
            I => \N__33464\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__33468\,
            I => \N__33461\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33458\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__33464\,
            I => \N__33455\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33452\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__33458\,
            I => \N__33449\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__33455\,
            I => r1_4
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33452\,
            I => r1_4
        );

    \I__6429\ : Odrv12
    port map (
            O => \N__33449\,
            I => r1_4
        );

    \I__6428\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \ALU.b_3_ns_1_4_cascade_\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33435\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33432\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__33435\,
            I => \N__33429\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33432\,
            I => \N__33426\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__33429\,
            I => \N__33421\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__33426\,
            I => \N__33421\
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__33421\,
            I => \ALU.r4_RNISLNE1Z0Z_4\
        );

    \I__6420\ : InMux
    port map (
            O => \N__33418\,
            I => \N__33415\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__33415\,
            I => \N__33412\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__33412\,
            I => \N__33408\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33404\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__33408\,
            I => \N__33401\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33398\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__33404\,
            I => \N__33395\
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__33401\,
            I => r0_2
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33398\,
            I => r0_2
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__33395\,
            I => r0_2
        );

    \I__6410\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33385\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33381\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__33384\,
            I => \N__33377\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__33381\,
            I => \N__33374\
        );

    \I__6406\ : CascadeMux
    port map (
            O => \N__33380\,
            I => \N__33371\
        );

    \I__6405\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33368\
        );

    \I__6404\ : Span4Mux_h
    port map (
            O => \N__33374\,
            I => \N__33365\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33362\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__33368\,
            I => \N__33359\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__33365\,
            I => r1_2
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__33362\,
            I => r1_2
        );

    \I__6399\ : Odrv12
    port map (
            O => \N__33359\,
            I => r1_2
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__33352\,
            I => \ALU.b_3_ns_1_2_cascade_\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33344\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33348\,
            I => \N__33341\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33337\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__33344\,
            I => \N__33334\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__33341\,
            I => \N__33331\
        );

    \I__6392\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33328\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__33337\,
            I => \N__33325\
        );

    \I__6390\ : Span4Mux_h
    port map (
            O => \N__33334\,
            I => \N__33322\
        );

    \I__6389\ : Span12Mux_s8_h
    port map (
            O => \N__33331\,
            I => \N__33319\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33328\,
            I => \N__33316\
        );

    \I__6387\ : Span4Mux_h
    port map (
            O => \N__33325\,
            I => \N__33313\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__33322\,
            I => \ALU.r4_RNIKDNE1Z0Z_2\
        );

    \I__6385\ : Odrv12
    port map (
            O => \N__33319\,
            I => \ALU.r4_RNIKDNE1Z0Z_2\
        );

    \I__6384\ : Odrv4
    port map (
            O => \N__33316\,
            I => \ALU.r4_RNIKDNE1Z0Z_2\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__33313\,
            I => \ALU.r4_RNIKDNE1Z0Z_2\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__33304\,
            I => \N__33300\
        );

    \I__6381\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33292\
        );

    \I__6380\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33285\
        );

    \I__6379\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33276\
        );

    \I__6378\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33276\
        );

    \I__6377\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33276\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33276\
        );

    \I__6375\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33273\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__33292\,
            I => \N__33270\
        );

    \I__6373\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33261\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33261\
        );

    \I__6371\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33261\
        );

    \I__6370\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33261\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__33285\,
            I => \N__33258\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__33276\,
            I => \N__33255\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__33273\,
            I => \b_fastZ0Z_2\
        );

    \I__6366\ : Odrv4
    port map (
            O => \N__33270\,
            I => \b_fastZ0Z_2\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33261\,
            I => \b_fastZ0Z_2\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__33258\,
            I => \b_fastZ0Z_2\
        );

    \I__6363\ : Odrv12
    port map (
            O => \N__33255\,
            I => \b_fastZ0Z_2\
        );

    \I__6362\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33241\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33238\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__33238\,
            I => \N__33234\
        );

    \I__6359\ : CascadeMux
    port map (
            O => \N__33237\,
            I => \N__33230\
        );

    \I__6358\ : Sp12to4
    port map (
            O => \N__33234\,
            I => \N__33227\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__33233\,
            I => \N__33224\
        );

    \I__6356\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33221\
        );

    \I__6355\ : Span12Mux_s8_h
    port map (
            O => \N__33227\,
            I => \N__33218\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33215\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33212\
        );

    \I__6352\ : Odrv12
    port map (
            O => \N__33218\,
            I => r1_3
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__33215\,
            I => r1_3
        );

    \I__6350\ : Odrv4
    port map (
            O => \N__33212\,
            I => r1_3
        );

    \I__6349\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33197\
        );

    \I__6348\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33197\
        );

    \I__6347\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33194\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33191\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__33197\,
            I => \N__33188\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33185\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33178\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__33188\,
            I => \N__33175\
        );

    \I__6341\ : Span4Mux_h
    port map (
            O => \N__33185\,
            I => \N__33171\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33168\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33161\
        );

    \I__6338\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33161\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33161\
        );

    \I__6336\ : Span4Mux_h
    port map (
            O => \N__33178\,
            I => \N__33156\
        );

    \I__6335\ : Span4Mux_h
    port map (
            O => \N__33175\,
            I => \N__33156\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33153\
        );

    \I__6333\ : Odrv4
    port map (
            O => \N__33171\,
            I => \b_fastZ0Z_0\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__33168\,
            I => \b_fastZ0Z_0\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33161\,
            I => \b_fastZ0Z_0\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__33156\,
            I => \b_fastZ0Z_0\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__33153\,
            I => \b_fastZ0Z_0\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33132\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33127\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33127\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33139\,
            I => \N__33124\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33121\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33114\
        );

    \I__6322\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33114\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33114\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33108\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33105\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33102\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33097\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33114\,
            I => \N__33097\
        );

    \I__6315\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33094\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33091\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33088\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__33108\,
            I => \N__33083\
        );

    \I__6311\ : Span4Mux_h
    port map (
            O => \N__33105\,
            I => \N__33083\
        );

    \I__6310\ : Span4Mux_h
    port map (
            O => \N__33102\,
            I => \N__33080\
        );

    \I__6309\ : Span4Mux_h
    port map (
            O => \N__33097\,
            I => \N__33077\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__33094\,
            I => \b_2_repZ0Z1\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__33091\,
            I => \b_2_repZ0Z1\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__33088\,
            I => \b_2_repZ0Z1\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__33083\,
            I => \b_2_repZ0Z1\
        );

    \I__6304\ : Odrv4
    port map (
            O => \N__33080\,
            I => \b_2_repZ0Z1\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__33077\,
            I => \b_2_repZ0Z1\
        );

    \I__6302\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33061\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__33061\,
            I => \N__33058\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__33058\,
            I => \N__33053\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33048\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33048\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__33053\,
            I => \N__33045\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__33048\,
            I => r4_3
        );

    \I__6295\ : Odrv4
    port map (
            O => \N__33045\,
            I => r4_3
        );

    \I__6294\ : CascadeMux
    port map (
            O => \N__33040\,
            I => \ALU.b_3_ns_1_3_cascade_\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33037\,
            I => \N__33031\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33031\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__33031\,
            I => \N__33027\
        );

    \I__6290\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33024\
        );

    \I__6289\ : Span4Mux_v
    port map (
            O => \N__33027\,
            I => \N__33021\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__33018\
        );

    \I__6287\ : Span4Mux_h
    port map (
            O => \N__33021\,
            I => \N__33013\
        );

    \I__6286\ : Span4Mux_v
    port map (
            O => \N__33018\,
            I => \N__33013\
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__33013\,
            I => \ALU.r4_RNIOHNE1Z0Z_3\
        );

    \I__6284\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__33007\,
            I => \N__33004\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__33004\,
            I => \N__33001\
        );

    \I__6281\ : Span4Mux_v
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__32998\,
            I => \ALU.rshift_10\
        );

    \I__6279\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32992\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32992\,
            I => \N__32989\
        );

    \I__6277\ : Span4Mux_h
    port map (
            O => \N__32989\,
            I => \N__32986\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__32986\,
            I => \ALU.madd_76_0\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__32983\,
            I => \ALU.lshift_3_ns_1_11_cascade_\
        );

    \I__6274\ : CascadeMux
    port map (
            O => \N__32980\,
            I => \N__32977\
        );

    \I__6273\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__32974\,
            I => \ALU.un9_addsub_axb_4\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__32968\,
            I => \N__32965\
        );

    \I__6269\ : Span4Mux_h
    port map (
            O => \N__32965\,
            I => \N__32962\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__32962\,
            I => \ALU.lshift_3_ns_1_9\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32956\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32951\
        );

    \I__6265\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32948\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32945\
        );

    \I__6263\ : Span4Mux_h
    port map (
            O => \N__32951\,
            I => \N__32940\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__32948\,
            I => \N__32940\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__32945\,
            I => r1_1
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__32940\,
            I => r1_1
        );

    \I__6259\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32932\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32929\
        );

    \I__6257\ : Span4Mux_h
    port map (
            O => \N__32929\,
            I => \N__32926\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__32926\,
            I => \ALU.r0_RNIE5LHZ0Z_1\
        );

    \I__6255\ : CascadeMux
    port map (
            O => \N__32923\,
            I => \ALU.rshift_3_ns_1_3_cascade_\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__32920\,
            I => \ALU.r0_12_prm_8_3_c_RNOZ0Z_3_cascade_\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32914\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32911\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__32911\,
            I => \N__32907\
        );

    \I__6250\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32904\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__32907\,
            I => \N__32901\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__32904\,
            I => \ALU.r5_RNI67NNKZ0Z_10\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__32901\,
            I => \ALU.r5_RNI67NNKZ0Z_10\
        );

    \I__6246\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32888\
        );

    \I__6245\ : CascadeMux
    port map (
            O => \N__32895\,
            I => \N__32884\
        );

    \I__6244\ : CascadeMux
    port map (
            O => \N__32894\,
            I => \N__32880\
        );

    \I__6243\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32877\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32874\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32871\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32868\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32887\,
            I => \N__32865\
        );

    \I__6238\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32856\
        );

    \I__6237\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32856\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32853\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__32877\,
            I => \N__32842\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32874\,
            I => \N__32842\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32842\
        );

    \I__6232\ : Span4Mux_v
    port map (
            O => \N__32868\,
            I => \N__32842\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32842\
        );

    \I__6230\ : CascadeMux
    port map (
            O => \N__32864\,
            I => \N__32838\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__32863\,
            I => \N__32835\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32831\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32827\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__32856\,
            I => \N__32824\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32821\
        );

    \I__6224\ : Span4Mux_v
    port map (
            O => \N__32842\,
            I => \N__32818\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__32841\,
            I => \N__32812\
        );

    \I__6222\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32807\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32807\
        );

    \I__6220\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32804\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__32831\,
            I => \N__32801\
        );

    \I__6218\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32798\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32827\,
            I => \N__32795\
        );

    \I__6216\ : Span4Mux_s2_h
    port map (
            O => \N__32824\,
            I => \N__32788\
        );

    \I__6215\ : Span4Mux_v
    port map (
            O => \N__32821\,
            I => \N__32788\
        );

    \I__6214\ : Span4Mux_s2_h
    port map (
            O => \N__32818\,
            I => \N__32788\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32781\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32781\
        );

    \I__6211\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32781\
        );

    \I__6210\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32778\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32775\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32768\
        );

    \I__6207\ : Span12Mux_h
    port map (
            O => \N__32801\,
            I => \N__32768\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__32798\,
            I => \N__32768\
        );

    \I__6205\ : Span4Mux_h
    port map (
            O => \N__32795\,
            I => \N__32763\
        );

    \I__6204\ : Span4Mux_h
    port map (
            O => \N__32788\,
            I => \N__32763\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32781\,
            I => \bZ0Z_1\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__32778\,
            I => \bZ0Z_1\
        );

    \I__6201\ : Odrv12
    port map (
            O => \N__32775\,
            I => \bZ0Z_1\
        );

    \I__6200\ : Odrv12
    port map (
            O => \N__32768\,
            I => \bZ0Z_1\
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__32763\,
            I => \bZ0Z_1\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32752\,
            I => \N__32749\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__32749\,
            I => \N__32745\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32741\
        );

    \I__6195\ : Span4Mux_v
    port map (
            O => \N__32745\,
            I => \N__32738\
        );

    \I__6194\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32735\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32732\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__32738\,
            I => \N__32729\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__32735\,
            I => \N__32726\
        );

    \I__6190\ : Odrv12
    port map (
            O => \N__32732\,
            I => \ALU.r6_RNI6TET1Z0Z_0\
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__32729\,
            I => \ALU.r6_RNI6TET1Z0Z_0\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__32726\,
            I => \ALU.r6_RNI6TET1Z0Z_0\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32715\
        );

    \I__6186\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32712\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32709\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32705\
        );

    \I__6183\ : Span4Mux_h
    port map (
            O => \N__32709\,
            I => \N__32702\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32699\
        );

    \I__6181\ : Odrv12
    port map (
            O => \N__32705\,
            I => \ALU.r4_RNIC5NE1Z0Z_0\
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__32702\,
            I => \ALU.r4_RNIC5NE1Z0Z_0\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32699\,
            I => \ALU.r4_RNIC5NE1Z0Z_0\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32692\,
            I => \N__32686\
        );

    \I__6177\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32686\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__32686\,
            I => \N__32681\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32685\,
            I => \N__32678\
        );

    \I__6174\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32672\
        );

    \I__6173\ : Span4Mux_s1_v
    port map (
            O => \N__32681\,
            I => \N__32667\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__32678\,
            I => \N__32667\
        );

    \I__6171\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32660\
        );

    \I__6170\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32660\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32657\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32652\
        );

    \I__6167\ : Span4Mux_h
    port map (
            O => \N__32667\,
            I => \N__32649\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32646\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32643\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32638\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32657\,
            I => \N__32638\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32635\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32632\
        );

    \I__6160\ : Span4Mux_v
    port map (
            O => \N__32652\,
            I => \N__32629\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__32649\,
            I => \N__32624\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32646\,
            I => \N__32624\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__32643\,
            I => \N__32621\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__32638\,
            I => \N__32616\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32616\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32613\
        );

    \I__6153\ : Sp12to4
    port map (
            O => \N__32629\,
            I => \N__32610\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__32624\,
            I => \N__32605\
        );

    \I__6151\ : Span4Mux_v
    port map (
            O => \N__32621\,
            I => \N__32605\
        );

    \I__6150\ : Span4Mux_h
    port map (
            O => \N__32616\,
            I => \N__32602\
        );

    \I__6149\ : Odrv12
    port map (
            O => \N__32613\,
            I => \ALU.r6_RNIBF8D2Z0Z_2\
        );

    \I__6148\ : Odrv12
    port map (
            O => \N__32610\,
            I => \ALU.r6_RNIBF8D2Z0Z_2\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__32605\,
            I => \ALU.r6_RNIBF8D2Z0Z_2\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__32602\,
            I => \ALU.r6_RNIBF8D2Z0Z_2\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32586\
        );

    \I__6144\ : CascadeMux
    port map (
            O => \N__32592\,
            I => \N__32583\
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__32591\,
            I => \N__32580\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32575\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32571\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__32586\,
            I => \N__32567\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32583\,
            I => \N__32564\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32559\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32559\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32556\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__32575\,
            I => \N__32553\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32574\,
            I => \N__32550\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__32571\,
            I => \N__32545\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32542\
        );

    \I__6131\ : Span4Mux_v
    port map (
            O => \N__32567\,
            I => \N__32537\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__32564\,
            I => \N__32537\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__32559\,
            I => \N__32534\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32556\,
            I => \N__32531\
        );

    \I__6127\ : Span4Mux_h
    port map (
            O => \N__32553\,
            I => \N__32526\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__32550\,
            I => \N__32526\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32521\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32521\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__32545\,
            I => \N__32518\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32542\,
            I => \N__32515\
        );

    \I__6121\ : Span4Mux_h
    port map (
            O => \N__32537\,
            I => \N__32510\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__32534\,
            I => \N__32510\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__32531\,
            I => \N__32507\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__32526\,
            I => \N__32504\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32521\,
            I => \N__32501\
        );

    \I__6116\ : Span4Mux_h
    port map (
            O => \N__32518\,
            I => \N__32498\
        );

    \I__6115\ : Span12Mux_s8_h
    port map (
            O => \N__32515\,
            I => \N__32495\
        );

    \I__6114\ : Span4Mux_v
    port map (
            O => \N__32510\,
            I => \N__32492\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__32507\,
            I => \N__32487\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__32504\,
            I => \N__32487\
        );

    \I__6111\ : Odrv12
    port map (
            O => \N__32501\,
            I => \ALU.r4_RNIHM992Z0Z_2\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__32498\,
            I => \ALU.r4_RNIHM992Z0Z_2\
        );

    \I__6109\ : Odrv12
    port map (
            O => \N__32495\,
            I => \ALU.r4_RNIHM992Z0Z_2\
        );

    \I__6108\ : Odrv4
    port map (
            O => \N__32492\,
            I => \ALU.r4_RNIHM992Z0Z_2\
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__32487\,
            I => \ALU.r4_RNIHM992Z0Z_2\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32473\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32465\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32461\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32457\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32454\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32448\
        );

    \I__6100\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32448\
        );

    \I__6099\ : Span4Mux_s1_v
    port map (
            O => \N__32465\,
            I => \N__32444\
        );

    \I__6098\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32441\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32438\
        );

    \I__6096\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32435\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__32457\,
            I => \N__32432\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32429\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32426\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32423\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32420\
        );

    \I__6090\ : Span4Mux_v
    port map (
            O => \N__32444\,
            I => \N__32417\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__32441\,
            I => \N__32414\
        );

    \I__6088\ : Span4Mux_s2_v
    port map (
            O => \N__32438\,
            I => \N__32407\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32435\,
            I => \N__32407\
        );

    \I__6086\ : Span4Mux_h
    port map (
            O => \N__32432\,
            I => \N__32407\
        );

    \I__6085\ : Span4Mux_h
    port map (
            O => \N__32429\,
            I => \N__32402\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32426\,
            I => \N__32402\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__32423\,
            I => \N__32397\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__32420\,
            I => \N__32397\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__32417\,
            I => \N__32394\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__32414\,
            I => \N__32389\
        );

    \I__6079\ : Span4Mux_v
    port map (
            O => \N__32407\,
            I => \N__32389\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__32402\,
            I => \N__32384\
        );

    \I__6077\ : Span4Mux_h
    port map (
            O => \N__32397\,
            I => \N__32384\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__32394\,
            I => \ALU.r6_RNI403D2Z0Z_4\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__32389\,
            I => \ALU.r6_RNI403D2Z0Z_4\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__32384\,
            I => \ALU.r6_RNI403D2Z0Z_4\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32369\
        );

    \I__6072\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32366\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32363\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__32374\,
            I => \N__32357\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32354\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32351\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32345\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32366\,
            I => \N__32345\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32342\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32339\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32336\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32331\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32331\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32328\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32325\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32322\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__32345\,
            I => \N__32319\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__32342\,
            I => \N__32312\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32312\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__32336\,
            I => \N__32312\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32331\,
            I => \N__32309\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__32328\,
            I => \N__32306\
        );

    \I__6051\ : Span4Mux_v
    port map (
            O => \N__32325\,
            I => \N__32303\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32322\,
            I => \N__32300\
        );

    \I__6049\ : Span4Mux_h
    port map (
            O => \N__32319\,
            I => \N__32295\
        );

    \I__6048\ : Span4Mux_v
    port map (
            O => \N__32312\,
            I => \N__32295\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__32309\,
            I => \N__32290\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__32306\,
            I => \N__32290\
        );

    \I__6045\ : Span4Mux_h
    port map (
            O => \N__32303\,
            I => \N__32283\
        );

    \I__6044\ : Span4Mux_v
    port map (
            O => \N__32300\,
            I => \N__32283\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__32295\,
            I => \N__32283\
        );

    \I__6042\ : Odrv4
    port map (
            O => \N__32290\,
            I => \ALU.r4_RNIQU992Z0Z_4\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__32283\,
            I => \ALU.r4_RNIQU992Z0Z_4\
        );

    \I__6040\ : CascadeMux
    port map (
            O => \N__32278\,
            I => \N__32273\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__32277\,
            I => \N__32269\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__32276\,
            I => \N__32266\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32258\
        );

    \I__6036\ : CascadeMux
    port map (
            O => \N__32272\,
            I => \N__32254\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32269\,
            I => \N__32249\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32249\
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__32265\,
            I => \N__32246\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__32264\,
            I => \N__32242\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__32263\,
            I => \N__32239\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__32262\,
            I => \N__32233\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__32261\,
            I => \N__32230\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__32258\,
            I => \N__32225\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__32257\,
            I => \N__32220\
        );

    \I__6026\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32217\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32249\,
            I => \N__32214\
        );

    \I__6024\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32211\
        );

    \I__6023\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32206\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32206\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32203\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__32238\,
            I => \N__32196\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__32237\,
            I => \N__32193\
        );

    \I__6018\ : CascadeMux
    port map (
            O => \N__32236\,
            I => \N__32190\
        );

    \I__6017\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32187\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32182\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__32229\,
            I => \N__32179\
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__32228\,
            I => \N__32175\
        );

    \I__6013\ : Span4Mux_s2_h
    port map (
            O => \N__32225\,
            I => \N__32170\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32224\,
            I => \N__32163\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32163\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32163\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32156\
        );

    \I__6008\ : Span4Mux_s2_v
    port map (
            O => \N__32214\,
            I => \N__32156\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__32211\,
            I => \N__32149\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__32206\,
            I => \N__32149\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__32203\,
            I => \N__32149\
        );

    \I__6004\ : CascadeMux
    port map (
            O => \N__32202\,
            I => \N__32146\
        );

    \I__6003\ : CascadeMux
    port map (
            O => \N__32201\,
            I => \N__32143\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__32200\,
            I => \N__32140\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32199\,
            I => \N__32133\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32133\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32133\
        );

    \I__5998\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32130\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32187\,
            I => \N__32126\
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__32186\,
            I => \N__32123\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__32185\,
            I => \N__32120\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32182\,
            I => \N__32117\
        );

    \I__5993\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32110\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32110\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32110\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__32174\,
            I => \N__32107\
        );

    \I__5989\ : CascadeMux
    port map (
            O => \N__32173\,
            I => \N__32103\
        );

    \I__5988\ : Span4Mux_h
    port map (
            O => \N__32170\,
            I => \N__32099\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32096\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32091\
        );

    \I__5985\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32091\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__32156\,
            I => \N__32086\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__32149\,
            I => \N__32086\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32083\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32078\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32078\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__32133\,
            I => \N__32075\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32072\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32069\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__32126\,
            I => \N__32066\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32063\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32060\
        );

    \I__5973\ : Span4Mux_s1_v
    port map (
            O => \N__32117\,
            I => \N__32055\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32055\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32050\
        );

    \I__5970\ : InMux
    port map (
            O => \N__32106\,
            I => \N__32050\
        );

    \I__5969\ : InMux
    port map (
            O => \N__32103\,
            I => \N__32045\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32045\
        );

    \I__5967\ : Span4Mux_v
    port map (
            O => \N__32099\,
            I => \N__32037\
        );

    \I__5966\ : Span4Mux_v
    port map (
            O => \N__32096\,
            I => \N__32037\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32034\
        );

    \I__5964\ : Sp12to4
    port map (
            O => \N__32086\,
            I => \N__32031\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__32083\,
            I => \N__32026\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__32078\,
            I => \N__32026\
        );

    \I__5961\ : Span4Mux_v
    port map (
            O => \N__32075\,
            I => \N__32023\
        );

    \I__5960\ : Span4Mux_h
    port map (
            O => \N__32072\,
            I => \N__32014\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32014\
        );

    \I__5958\ : Span4Mux_h
    port map (
            O => \N__32066\,
            I => \N__32014\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__32063\,
            I => \N__32014\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__32060\,
            I => \N__32011\
        );

    \I__5955\ : Span4Mux_h
    port map (
            O => \N__32055\,
            I => \N__32004\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__32004\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__32045\,
            I => \N__32004\
        );

    \I__5952\ : InMux
    port map (
            O => \N__32044\,
            I => \N__31997\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32043\,
            I => \N__31997\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32042\,
            I => \N__31997\
        );

    \I__5949\ : Span4Mux_h
    port map (
            O => \N__32037\,
            I => \N__31994\
        );

    \I__5948\ : Sp12to4
    port map (
            O => \N__32034\,
            I => \N__31987\
        );

    \I__5947\ : Span12Mux_h
    port map (
            O => \N__32031\,
            I => \N__31987\
        );

    \I__5946\ : Span12Mux_s5_h
    port map (
            O => \N__32026\,
            I => \N__31987\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__32023\,
            I => \N__31982\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__32014\,
            I => \N__31982\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__32011\,
            I => \N__31977\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__32004\,
            I => \N__31977\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__31997\,
            I => \aZ0Z_1\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__31994\,
            I => \aZ0Z_1\
        );

    \I__5939\ : Odrv12
    port map (
            O => \N__31987\,
            I => \aZ0Z_1\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__31982\,
            I => \aZ0Z_1\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__31977\,
            I => \aZ0Z_1\
        );

    \I__5936\ : CascadeMux
    port map (
            O => \N__31966\,
            I => \ALU.un2_addsub_axb_4_cascade_\
        );

    \I__5935\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31960\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31957\
        );

    \I__5933\ : Odrv12
    port map (
            O => \N__31957\,
            I => \ALU.un9_addsub_axb_3\
        );

    \I__5932\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31951\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31948\
        );

    \I__5930\ : Span4Mux_v
    port map (
            O => \N__31948\,
            I => \N__31945\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__31945\,
            I => \N__31942\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__31942\,
            I => \N__31939\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__31939\,
            I => \ALU.madd_490_5\
        );

    \I__5926\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31931\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31928\
        );

    \I__5924\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31925\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31918\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31915\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31912\
        );

    \I__5920\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31908\
        );

    \I__5919\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31903\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31903\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31898\
        );

    \I__5916\ : Span4Mux_h
    port map (
            O => \N__31918\,
            I => \N__31893\
        );

    \I__5915\ : Span4Mux_s1_v
    port map (
            O => \N__31915\,
            I => \N__31893\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__31912\,
            I => \N__31890\
        );

    \I__5913\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31887\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31882\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__31903\,
            I => \N__31882\
        );

    \I__5910\ : InMux
    port map (
            O => \N__31902\,
            I => \N__31879\
        );

    \I__5909\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31876\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31873\
        );

    \I__5907\ : Span4Mux_v
    port map (
            O => \N__31893\,
            I => \N__31870\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__31890\,
            I => \N__31863\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31863\
        );

    \I__5904\ : Span4Mux_h
    port map (
            O => \N__31882\,
            I => \N__31863\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31879\,
            I => \N__31858\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__31876\,
            I => \N__31858\
        );

    \I__5901\ : Span4Mux_v
    port map (
            O => \N__31873\,
            I => \N__31853\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__31870\,
            I => \N__31853\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__31863\,
            I => \N__31850\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__31858\,
            I => \N__31847\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__31853\,
            I => \ALU.r6_RNIFJ8D2Z0Z_3\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__31850\,
            I => \ALU.r6_RNIFJ8D2Z0Z_3\
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__31847\,
            I => \ALU.r6_RNIFJ8D2Z0Z_3\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__31840\,
            I => \N__31836\
        );

    \I__5893\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31830\
        );

    \I__5892\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31825\
        );

    \I__5891\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31819\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31834\,
            I => \N__31819\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__31833\,
            I => \N__31816\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31813\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31810\
        );

    \I__5886\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31807\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__31825\,
            I => \N__31804\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31824\,
            I => \N__31801\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31819\,
            I => \N__31798\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31793\
        );

    \I__5881\ : Span4Mux_v
    port map (
            O => \N__31813\,
            I => \N__31788\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31788\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__31807\,
            I => \N__31785\
        );

    \I__5878\ : Span4Mux_s3_v
    port map (
            O => \N__31804\,
            I => \N__31782\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31779\
        );

    \I__5876\ : Span4Mux_v
    port map (
            O => \N__31798\,
            I => \N__31776\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31771\
        );

    \I__5874\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31771\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__31793\,
            I => \N__31768\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__31788\,
            I => \N__31765\
        );

    \I__5871\ : Span4Mux_s3_v
    port map (
            O => \N__31785\,
            I => \N__31760\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__31782\,
            I => \N__31760\
        );

    \I__5869\ : Span4Mux_v
    port map (
            O => \N__31779\,
            I => \N__31755\
        );

    \I__5868\ : Span4Mux_h
    port map (
            O => \N__31776\,
            I => \N__31755\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31771\,
            I => \N__31752\
        );

    \I__5866\ : Odrv12
    port map (
            O => \N__31768\,
            I => \ALU.r4_RNIMQ992Z0Z_3\
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__31765\,
            I => \ALU.r4_RNIMQ992Z0Z_3\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__31760\,
            I => \ALU.r4_RNIMQ992Z0Z_3\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__31755\,
            I => \ALU.r4_RNIMQ992Z0Z_3\
        );

    \I__5862\ : Odrv12
    port map (
            O => \N__31752\,
            I => \ALU.r4_RNIMQ992Z0Z_3\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31735\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__31740\,
            I => \N__31732\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31726\
        );

    \I__5858\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31726\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__31735\,
            I => \N__31723\
        );

    \I__5856\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31714\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31714\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31726\,
            I => \N__31711\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__31723\,
            I => \N__31708\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31701\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31701\
        );

    \I__5850\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31701\
        );

    \I__5849\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31698\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__31714\,
            I => \N__31695\
        );

    \I__5847\ : Span4Mux_s3_v
    port map (
            O => \N__31711\,
            I => \N__31692\
        );

    \I__5846\ : Span4Mux_h
    port map (
            O => \N__31708\,
            I => \N__31687\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31687\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31698\,
            I => \N__31684\
        );

    \I__5843\ : Span4Mux_s3_v
    port map (
            O => \N__31695\,
            I => \N__31681\
        );

    \I__5842\ : Span4Mux_v
    port map (
            O => \N__31692\,
            I => \N__31678\
        );

    \I__5841\ : Span4Mux_h
    port map (
            O => \N__31687\,
            I => \N__31675\
        );

    \I__5840\ : Odrv12
    port map (
            O => \N__31684\,
            I => \ALU.r4_RNIDI992Z0Z_1\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__31681\,
            I => \ALU.r4_RNIDI992Z0Z_1\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__31678\,
            I => \ALU.r4_RNIDI992Z0Z_1\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__31675\,
            I => \ALU.r4_RNIDI992Z0Z_1\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31661\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31665\,
            I => \N__31656\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31656\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31652\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N__31649\
        );

    \I__5831\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31644\
        );

    \I__5830\ : Span4Mux_s1_v
    port map (
            O => \N__31652\,
            I => \N__31641\
        );

    \I__5829\ : Span4Mux_s1_v
    port map (
            O => \N__31649\,
            I => \N__31638\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31633\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31633\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__31644\,
            I => \N__31627\
        );

    \I__5825\ : Span4Mux_v
    port map (
            O => \N__31641\,
            I => \N__31622\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__31638\,
            I => \N__31622\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31633\,
            I => \N__31619\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31612\
        );

    \I__5821\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31612\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31612\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__31627\,
            I => \N__31609\
        );

    \I__5818\ : Span4Mux_h
    port map (
            O => \N__31622\,
            I => \N__31606\
        );

    \I__5817\ : Span12Mux_s8_v
    port map (
            O => \N__31619\,
            I => \N__31603\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__31612\,
            I => \N__31600\
        );

    \I__5815\ : Odrv4
    port map (
            O => \N__31609\,
            I => \ALU.r6_RNI7B8D2Z0Z_1\
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__31606\,
            I => \ALU.r6_RNI7B8D2Z0Z_1\
        );

    \I__5813\ : Odrv12
    port map (
            O => \N__31603\,
            I => \ALU.r6_RNI7B8D2Z0Z_1\
        );

    \I__5812\ : Odrv12
    port map (
            O => \N__31600\,
            I => \ALU.r6_RNI7B8D2Z0Z_1\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31582\
        );

    \I__5810\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31582\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31582\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__5807\ : Odrv4
    port map (
            O => \N__31579\,
            I => \ALU.a1_b_3\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__31576\,
            I => \N__31572\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__31575\,
            I => \N__31569\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31564\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31564\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31560\
        );

    \I__5801\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31557\
        );

    \I__5800\ : Span4Mux_s1_v
    port map (
            O => \N__31560\,
            I => \N__31554\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__31557\,
            I => \N__31551\
        );

    \I__5798\ : Span4Mux_s2_h
    port map (
            O => \N__31554\,
            I => \N__31548\
        );

    \I__5797\ : Span4Mux_h
    port map (
            O => \N__31551\,
            I => \N__31543\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__31548\,
            I => \N__31543\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__31543\,
            I => \ALU.madd_135_0\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31537\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31537\,
            I => \N__31534\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__31534\,
            I => \ALU.lshift_3_ns_1_6\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31531\,
            I => \N__31528\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__31528\,
            I => \N__31525\
        );

    \I__5789\ : Span4Mux_s3_v
    port map (
            O => \N__31525\,
            I => \N__31522\
        );

    \I__5788\ : Span4Mux_h
    port map (
            O => \N__31522\,
            I => \N__31519\
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__31519\,
            I => \ALU.lshift_3_ns_1_7\
        );

    \I__5786\ : InMux
    port map (
            O => \N__31516\,
            I => \ALU.r0_12_s1_13\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31510\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31507\
        );

    \I__5783\ : Odrv12
    port map (
            O => \N__31507\,
            I => \ALU.r0_12_s1_13_THRU_CO\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__31504\,
            I => \N__31501\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31498\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31498\,
            I => \ALU.r0_12_prm_1_13_s1_c_RNOZ0\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__31495\,
            I => \ALU.rshift_3_ns_1_2_cascade_\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31489\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__31486\,
            I => \N__31483\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__31483\,
            I => \N__31480\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__31480\,
            I => \ALU.r0_12_prm_7_13_s1_c_RNOZ0\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__31477\,
            I => \N__31473\
        );

    \I__5772\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31470\
        );

    \I__5771\ : InMux
    port map (
            O => \N__31473\,
            I => \N__31467\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31470\,
            I => \N__31464\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31461\
        );

    \I__5768\ : Span4Mux_v
    port map (
            O => \N__31464\,
            I => \N__31458\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__31461\,
            I => \N__31455\
        );

    \I__5766\ : Span4Mux_h
    port map (
            O => \N__31458\,
            I => \N__31452\
        );

    \I__5765\ : Sp12to4
    port map (
            O => \N__31455\,
            I => \N__31449\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__31452\,
            I => \ALU.r5_RNID2JJ9_0Z0Z_13\
        );

    \I__5763\ : Odrv12
    port map (
            O => \N__31449\,
            I => \ALU.r5_RNID2JJ9_0Z0Z_13\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31441\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__31441\,
            I => \N__31438\
        );

    \I__5760\ : Span4Mux_h
    port map (
            O => \N__31438\,
            I => \N__31435\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__31435\,
            I => \ALU.r0_12_prm_6_13_s1_c_RNOZ0\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31429\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31425\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__31425\,
            I => \N__31419\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31416\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__31419\,
            I => \ALU.un14_log_0_i_13\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__31416\,
            I => \ALU.un14_log_0_i_13\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31408\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__31408\,
            I => \N__31405\
        );

    \I__5749\ : Span4Mux_h
    port map (
            O => \N__31405\,
            I => \N__31402\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__31402\,
            I => \ALU.r0_12_prm_5_13_s1_c_RNOZ0\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__31399\,
            I => \N__31395\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__31398\,
            I => \N__31392\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31389\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31386\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31389\,
            I => \N__31383\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31378\
        );

    \I__5741\ : Span4Mux_h
    port map (
            O => \N__31383\,
            I => \N__31378\
        );

    \I__5740\ : Span4Mux_h
    port map (
            O => \N__31378\,
            I => \N__31375\
        );

    \I__5739\ : Odrv4
    port map (
            O => \N__31375\,
            I => \ALU.r5_RNID2JJ9_1Z0Z_13\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31369\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__31369\,
            I => \N__31366\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__31366\,
            I => \N__31363\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__31363\,
            I => \ALU.r0_12_prm_4_13_s1_c_RNOZ0\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__31360\,
            I => \N__31356\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31353\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31350\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31353\,
            I => \N__31345\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31350\,
            I => \N__31345\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__31345\,
            I => \ALU.a_i_13\
        );

    \I__5728\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31339\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31339\,
            I => \ALU.rshift_10_ns_1_3\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__31336\,
            I => \ALU.r5_RNI465TIZ0Z_13_cascade_\
        );

    \I__5725\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31330\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__31330\,
            I => \N__31327\
        );

    \I__5723\ : Span4Mux_v
    port map (
            O => \N__31327\,
            I => \N__31324\
        );

    \I__5722\ : Span4Mux_v
    port map (
            O => \N__31324\,
            I => \N__31321\
        );

    \I__5721\ : Odrv4
    port map (
            O => \N__31321\,
            I => \ALU.r5_RNIOL1S71Z0Z_10\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__31318\,
            I => \N__31315\
        );

    \I__5719\ : InMux
    port map (
            O => \N__31315\,
            I => \N__31312\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__31312\,
            I => \N__31309\
        );

    \I__5717\ : Span4Mux_h
    port map (
            O => \N__31309\,
            I => \N__31306\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__31306\,
            I => \ALU.r0_12_prm_5_12_s0_c_RNOZ0\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__31303\,
            I => \N__31300\
        );

    \I__5714\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31297\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31294\
        );

    \I__5712\ : Span4Mux_v
    port map (
            O => \N__31294\,
            I => \N__31291\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__31291\,
            I => \N__31288\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__31288\,
            I => \ALU.r0_12_prm_8_11_s0_c_RNOZ0\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__31285\,
            I => \N__31282\
        );

    \I__5708\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31279\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__31279\,
            I => \N__31276\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__31276\,
            I => \N__31273\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__31273\,
            I => \ALU.r0_12_prm_7_12_s0_c_RNOZ0\
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__31270\,
            I => \N__31267\
        );

    \I__5703\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31261\
        );

    \I__5701\ : Span4Mux_v
    port map (
            O => \N__31261\,
            I => \N__31258\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__5699\ : Sp12to4
    port map (
            O => \N__31255\,
            I => \N__31252\
        );

    \I__5698\ : Odrv12
    port map (
            O => \N__31252\,
            I => \ALU.r0_12_prm_6_12_s0_c_RNOZ0\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__31249\,
            I => \N__31246\
        );

    \I__5696\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31243\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__31243\,
            I => \N__31240\
        );

    \I__5694\ : Span4Mux_h
    port map (
            O => \N__31240\,
            I => \N__31237\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__31237\,
            I => \ALU.r0_12_prm_2_15_s1_c_RNOZ0\
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__31234\,
            I => \N__31231\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31228\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__31228\,
            I => \N__31225\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__31225\,
            I => \N__31222\
        );

    \I__5688\ : Span4Mux_h
    port map (
            O => \N__31222\,
            I => \N__31219\
        );

    \I__5687\ : Odrv4
    port map (
            O => \N__31219\,
            I => \ALU.r0_12_prm_2_13_s0_c_RNOZ0\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__31216\,
            I => \N__31213\
        );

    \I__5685\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31210\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31210\,
            I => \N__31207\
        );

    \I__5683\ : Span4Mux_h
    port map (
            O => \N__31207\,
            I => \N__31204\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__31204\,
            I => \ALU.r0_12_prm_1_14_s0_c_RNOZ0\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__31201\,
            I => \N__31198\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31195\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__31195\,
            I => \N__31192\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__31192\,
            I => \N__31189\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__31189\,
            I => \ALU.r0_12_prm_8_15_s1_c_RNOZ0\
        );

    \I__5676\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31183\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__31183\,
            I => \ALU.r0_12_prm_3_9_s0_sf\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__31180\,
            I => \N__31177\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31177\,
            I => \N__31174\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__31174\,
            I => \N__31171\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__31171\,
            I => \N__31168\
        );

    \I__5670\ : Span4Mux_h
    port map (
            O => \N__31168\,
            I => \N__31165\
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__31165\,
            I => \ALU.r0_12_prm_2_9_s0_c_RNOZ0\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31159\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31159\,
            I => \N__31156\
        );

    \I__5666\ : Span4Mux_v
    port map (
            O => \N__31156\,
            I => \N__31153\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__31153\,
            I => \ALU.mult_9\
        );

    \I__5664\ : InMux
    port map (
            O => \N__31150\,
            I => \ALU.r0_12_s0_9\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31143\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31140\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__31143\,
            I => \N__31135\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__31140\,
            I => \N__31135\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__31135\,
            I => \N__31131\
        );

    \I__5658\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31128\
        );

    \I__5657\ : Span4Mux_h
    port map (
            O => \N__31131\,
            I => \N__31123\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31123\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__31123\,
            I => r0_9
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31114\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__31114\,
            I => \N__31111\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__31111\,
            I => \N__31108\
        );

    \I__5650\ : Span4Mux_h
    port map (
            O => \N__31108\,
            I => \N__31105\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__31105\,
            I => \N__31102\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__31102\,
            I => \ALU.r0_12_prm_8_11_s1_c_RNOZ0\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__31099\,
            I => \ALU.a_3_ns_1_4_cascade_\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31092\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__31092\,
            I => \N__31081\
        );

    \I__5643\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31072\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31072\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31072\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31072\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__31085\,
            I => \N__31069\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__31084\,
            I => \N__31063\
        );

    \I__5637\ : Span4Mux_s1_h
    port map (
            O => \N__31081\,
            I => \N__31057\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31072\,
            I => \N__31054\
        );

    \I__5635\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31047\
        );

    \I__5634\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31047\
        );

    \I__5633\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31047\
        );

    \I__5632\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31044\
        );

    \I__5631\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31041\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31062\,
            I => \N__31038\
        );

    \I__5629\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31033\
        );

    \I__5628\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31033\
        );

    \I__5627\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31028\
        );

    \I__5626\ : Span4Mux_h
    port map (
            O => \N__31054\,
            I => \N__31028\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__31047\,
            I => \N__31025\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__31044\,
            I => \a_fastZ0Z_2\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__31041\,
            I => \a_fastZ0Z_2\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__31038\,
            I => \a_fastZ0Z_2\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__31033\,
            I => \a_fastZ0Z_2\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__31028\,
            I => \a_fastZ0Z_2\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__31025\,
            I => \a_fastZ0Z_2\
        );

    \I__5618\ : CascadeMux
    port map (
            O => \N__31012\,
            I => \N__31007\
        );

    \I__5617\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31004\
        );

    \I__5616\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31001\
        );

    \I__5615\ : InMux
    port map (
            O => \N__31007\,
            I => \N__30998\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__31004\,
            I => \N__30995\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__31001\,
            I => \N__30990\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30990\
        );

    \I__5611\ : Span4Mux_h
    port map (
            O => \N__30995\,
            I => \N__30987\
        );

    \I__5610\ : Span4Mux_h
    port map (
            O => \N__30990\,
            I => \N__30984\
        );

    \I__5609\ : Odrv4
    port map (
            O => \N__30987\,
            I => r1_9
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__30984\,
            I => r1_9
        );

    \I__5607\ : InMux
    port map (
            O => \N__30979\,
            I => \N__30965\
        );

    \I__5606\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30965\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30958\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30976\,
            I => \N__30958\
        );

    \I__5603\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30958\
        );

    \I__5602\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30947\
        );

    \I__5601\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30947\
        );

    \I__5600\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30947\
        );

    \I__5599\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30947\
        );

    \I__5598\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30947\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__30965\,
            I => \N__30944\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__30958\,
            I => \a_fastZ0Z_0\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__30947\,
            I => \a_fastZ0Z_0\
        );

    \I__5594\ : Odrv4
    port map (
            O => \N__30944\,
            I => \a_fastZ0Z_0\
        );

    \I__5593\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30931\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30931\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__30931\,
            I => \N__30921\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30916\
        );

    \I__5589\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30916\
        );

    \I__5588\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30909\
        );

    \I__5587\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30906\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30903\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30925\,
            I => \N__30900\
        );

    \I__5584\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30897\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__30921\,
            I => \N__30894\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30891\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30880\
        );

    \I__5580\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30880\
        );

    \I__5579\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30875\
        );

    \I__5578\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30875\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__30909\,
            I => \N__30872\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__30906\,
            I => \N__30867\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__30903\,
            I => \N__30867\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30900\,
            I => \N__30862\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__30897\,
            I => \N__30862\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__30894\,
            I => \N__30857\
        );

    \I__5571\ : Span4Mux_v
    port map (
            O => \N__30891\,
            I => \N__30857\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30852\
        );

    \I__5569\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30852\
        );

    \I__5568\ : InMux
    port map (
            O => \N__30888\,
            I => \N__30845\
        );

    \I__5567\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30845\
        );

    \I__5566\ : InMux
    port map (
            O => \N__30886\,
            I => \N__30845\
        );

    \I__5565\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30842\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30833\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30833\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__30872\,
            I => \N__30833\
        );

    \I__5561\ : Span4Mux_h
    port map (
            O => \N__30867\,
            I => \N__30833\
        );

    \I__5560\ : Span4Mux_v
    port map (
            O => \N__30862\,
            I => \N__30828\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__30857\,
            I => \N__30828\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__30852\,
            I => \a_2_repZ0Z2\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__30845\,
            I => \a_2_repZ0Z2\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__30842\,
            I => \a_2_repZ0Z2\
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__30833\,
            I => \a_2_repZ0Z2\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__30828\,
            I => \a_2_repZ0Z2\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__30817\,
            I => \ALU.a_3_ns_1_9_cascade_\
        );

    \I__5552\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30808\
        );

    \I__5551\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30805\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30812\,
            I => \N__30802\
        );

    \I__5549\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30799\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__30808\,
            I => \N__30796\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__30805\,
            I => \N__30791\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30802\,
            I => \N__30791\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__30799\,
            I => \N__30788\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__30796\,
            I => \N__30785\
        );

    \I__5543\ : Span4Mux_h
    port map (
            O => \N__30791\,
            I => \N__30782\
        );

    \I__5542\ : Span4Mux_h
    port map (
            O => \N__30788\,
            I => \N__30779\
        );

    \I__5541\ : Span4Mux_h
    port map (
            O => \N__30785\,
            I => \N__30774\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__30782\,
            I => \N__30774\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__30779\,
            I => \ALU.r4_RNIEJA92Z0Z_9\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__30774\,
            I => \ALU.r4_RNIEJA92Z0Z_9\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__30769\,
            I => \N__30766\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30763\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30760\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__30760\,
            I => \N__30757\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__30757\,
            I => \N__30754\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__30754\,
            I => \ALU.r0_12_prm_6_9_s0_c_RNOZ0\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30751\,
            I => \N__30748\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__30748\,
            I => \N__30745\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__30745\,
            I => \N__30742\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__30742\,
            I => \N__30737\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30732\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30732\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__30737\,
            I => r0_7
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30732\,
            I => r0_7
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__30727\,
            I => \ALU.a_3_ns_1_7_cascade_\
        );

    \I__5522\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30719\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30716\
        );

    \I__5520\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30712\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__30719\,
            I => \N__30708\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30705\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30702\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__30712\,
            I => \N__30699\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30696\
        );

    \I__5514\ : Span4Mux_h
    port map (
            O => \N__30708\,
            I => \N__30693\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__30705\,
            I => \N__30688\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30702\,
            I => \N__30688\
        );

    \I__5511\ : Span4Mux_v
    port map (
            O => \N__30699\,
            I => \N__30685\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30696\,
            I => \N__30682\
        );

    \I__5509\ : Span4Mux_h
    port map (
            O => \N__30693\,
            I => \N__30679\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__30688\,
            I => \N__30676\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__30685\,
            I => \N__30671\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__30682\,
            I => \N__30671\
        );

    \I__5505\ : Odrv4
    port map (
            O => \N__30679\,
            I => \ALU.r4_RNI6BA92Z0Z_7\
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__30676\,
            I => \ALU.r4_RNI6BA92Z0Z_7\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__30671\,
            I => \ALU.r4_RNI6BA92Z0Z_7\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__30664\,
            I => \N__30660\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__30663\,
            I => \N__30657\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30653\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30650\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30647\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30653\,
            I => \N__30644\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30650\,
            I => \N__30641\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__30647\,
            I => \N__30638\
        );

    \I__5494\ : Span12Mux_s10_v
    port map (
            O => \N__30644\,
            I => \N__30635\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__30641\,
            I => \N__30632\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__30638\,
            I => r1_8
        );

    \I__5491\ : Odrv12
    port map (
            O => \N__30635\,
            I => r1_8
        );

    \I__5490\ : Odrv4
    port map (
            O => \N__30632\,
            I => r1_8
        );

    \I__5489\ : CascadeMux
    port map (
            O => \N__30625\,
            I => \ALU.a_3_ns_1_8_cascade_\
        );

    \I__5488\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30618\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__30621\,
            I => \N__30615\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__30618\,
            I => \N__30610\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30605\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30605\
        );

    \I__5483\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30602\
        );

    \I__5482\ : Span4Mux_v
    port map (
            O => \N__30610\,
            I => \N__30599\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30605\,
            I => \N__30594\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30602\,
            I => \N__30594\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__30599\,
            I => \N__30591\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__30594\,
            I => \N__30588\
        );

    \I__5477\ : Odrv4
    port map (
            O => \N__30591\,
            I => \ALU.r4_RNIAFA92Z0Z_8\
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__30588\,
            I => \ALU.r4_RNIAFA92Z0Z_8\
        );

    \I__5475\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30580\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30580\,
            I => \N__30577\
        );

    \I__5473\ : Odrv4
    port map (
            O => \N__30577\,
            I => \ALU.a_3_ns_1_3\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__30574\,
            I => \ALU.a_3_ns_1_2_cascade_\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30564\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30560\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30554\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30550\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30547\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30564\,
            I => \N__30544\
        );

    \I__5465\ : CascadeMux
    port map (
            O => \N__30563\,
            I => \N__30538\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__30560\,
            I => \N__30535\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30528\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30528\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30528\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30554\,
            I => \N__30525\
        );

    \I__5459\ : InMux
    port map (
            O => \N__30553\,
            I => \N__30522\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__30550\,
            I => \N__30515\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30547\,
            I => \N__30515\
        );

    \I__5456\ : Span4Mux_v
    port map (
            O => \N__30544\,
            I => \N__30515\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30506\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30542\,
            I => \N__30506\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30506\
        );

    \I__5452\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30506\
        );

    \I__5451\ : Span4Mux_h
    port map (
            O => \N__30535\,
            I => \N__30503\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30528\,
            I => \N__30498\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__30525\,
            I => \N__30498\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30522\,
            I => \a_2_repZ0Z1\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__30515\,
            I => \a_2_repZ0Z1\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__30506\,
            I => \a_2_repZ0Z1\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__30503\,
            I => \a_2_repZ0Z1\
        );

    \I__5444\ : Odrv4
    port map (
            O => \N__30498\,
            I => \a_2_repZ0Z1\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30484\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__30484\,
            I => \N__30481\
        );

    \I__5441\ : Span4Mux_h
    port map (
            O => \N__30481\,
            I => \N__30476\
        );

    \I__5440\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30473\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__30479\,
            I => \N__30470\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__30476\,
            I => \N__30465\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30473\,
            I => \N__30465\
        );

    \I__5436\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30462\
        );

    \I__5435\ : Span4Mux_v
    port map (
            O => \N__30465\,
            I => \N__30459\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30456\
        );

    \I__5433\ : Odrv4
    port map (
            O => \N__30459\,
            I => r1_15
        );

    \I__5432\ : Odrv4
    port map (
            O => \N__30456\,
            I => r1_15
        );

    \I__5431\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30448\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30448\,
            I => \N__30444\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30441\
        );

    \I__5428\ : Span4Mux_h
    port map (
            O => \N__30444\,
            I => \N__30438\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30435\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__30438\,
            I => \N__30429\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__30435\,
            I => \N__30429\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30426\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__30429\,
            I => r5_15
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30426\,
            I => r5_15
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__30421\,
            I => \TXbuffer_18_10_ns_1_7_cascade_\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__30418\,
            I => \N__30411\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__30417\,
            I => \N__30408\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__30416\,
            I => \N__30405\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__30415\,
            I => \N__30402\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__30414\,
            I => \N__30399\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30389\
        );

    \I__5414\ : InMux
    port map (
            O => \N__30408\,
            I => \N__30389\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30381\
        );

    \I__5412\ : InMux
    port map (
            O => \N__30402\,
            I => \N__30381\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30378\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__30398\,
            I => \N__30375\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__30397\,
            I => \N__30372\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__30396\,
            I => \N__30368\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__30395\,
            I => \N__30365\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__30394\,
            I => \N__30361\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30356\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__30388\,
            I => \N__30351\
        );

    \I__5403\ : CascadeMux
    port map (
            O => \N__30387\,
            I => \N__30348\
        );

    \I__5402\ : InMux
    port map (
            O => \N__30386\,
            I => \N__30345\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__30381\,
            I => \N__30340\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__30378\,
            I => \N__30340\
        );

    \I__5399\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30337\
        );

    \I__5398\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30331\
        );

    \I__5397\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30331\
        );

    \I__5396\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30328\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30325\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__30364\,
            I => \N__30321\
        );

    \I__5393\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30318\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__30360\,
            I => \N__30314\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__30359\,
            I => \N__30311\
        );

    \I__5390\ : Span4Mux_v
    port map (
            O => \N__30356\,
            I => \N__30306\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__30355\,
            I => \N__30300\
        );

    \I__5388\ : CascadeMux
    port map (
            O => \N__30354\,
            I => \N__30297\
        );

    \I__5387\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30292\
        );

    \I__5386\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30292\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__30345\,
            I => \N__30285\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__30340\,
            I => \N__30285\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30337\,
            I => \N__30285\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__30336\,
            I => \N__30282\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__30331\,
            I => \N__30276\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__30328\,
            I => \N__30276\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__30325\,
            I => \N__30273\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__30324\,
            I => \N__30270\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30265\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30262\
        );

    \I__5375\ : InMux
    port map (
            O => \N__30317\,
            I => \N__30259\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30256\
        );

    \I__5373\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30253\
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__30310\,
            I => \N__30250\
        );

    \I__5371\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30247\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__30306\,
            I => \N__30244\
        );

    \I__5369\ : InMux
    port map (
            O => \N__30305\,
            I => \N__30241\
        );

    \I__5368\ : CascadeMux
    port map (
            O => \N__30304\,
            I => \N__30237\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30230\
        );

    \I__5366\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30230\
        );

    \I__5365\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30230\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30225\
        );

    \I__5363\ : Span4Mux_h
    port map (
            O => \N__30285\,
            I => \N__30225\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30220\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30220\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__30276\,
            I => \N__30215\
        );

    \I__5359\ : Span4Mux_v
    port map (
            O => \N__30273\,
            I => \N__30215\
        );

    \I__5358\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30210\
        );

    \I__5357\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30210\
        );

    \I__5356\ : CascadeMux
    port map (
            O => \N__30268\,
            I => \N__30205\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__30265\,
            I => \N__30202\
        );

    \I__5354\ : Span4Mux_v
    port map (
            O => \N__30262\,
            I => \N__30193\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__30259\,
            I => \N__30193\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__30256\,
            I => \N__30193\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__30253\,
            I => \N__30193\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30190\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__30247\,
            I => \N__30183\
        );

    \I__5348\ : Sp12to4
    port map (
            O => \N__30244\,
            I => \N__30183\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__30241\,
            I => \N__30183\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30178\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30178\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__30230\,
            I => \N__30175\
        );

    \I__5343\ : Span4Mux_s1_h
    port map (
            O => \N__30225\,
            I => \N__30172\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__30220\,
            I => \N__30167\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__30215\,
            I => \N__30167\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__30210\,
            I => \N__30164\
        );

    \I__5339\ : InMux
    port map (
            O => \N__30209\,
            I => \N__30161\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30208\,
            I => \N__30156\
        );

    \I__5337\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30156\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__30202\,
            I => \N__30153\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__30193\,
            I => \N__30150\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__30190\,
            I => \N__30145\
        );

    \I__5333\ : Span12Mux_h
    port map (
            O => \N__30183\,
            I => \N__30145\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30138\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__30175\,
            I => \N__30138\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__30172\,
            I => \N__30138\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__30167\,
            I => \N__30135\
        );

    \I__5328\ : Odrv12
    port map (
            O => \N__30164\,
            I => \clkdivZ0Z_7\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30161\,
            I => \clkdivZ0Z_7\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30156\,
            I => \clkdivZ0Z_7\
        );

    \I__5325\ : Odrv4
    port map (
            O => \N__30153\,
            I => \clkdivZ0Z_7\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__30150\,
            I => \clkdivZ0Z_7\
        );

    \I__5323\ : Odrv12
    port map (
            O => \N__30145\,
            I => \clkdivZ0Z_7\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__30138\,
            I => \clkdivZ0Z_7\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__30135\,
            I => \clkdivZ0Z_7\
        );

    \I__5320\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30114\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30111\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30108\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__30111\,
            I => \N__30104\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__30108\,
            I => \N__30101\
        );

    \I__5315\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30098\
        );

    \I__5314\ : Span4Mux_h
    port map (
            O => \N__30104\,
            I => \N__30095\
        );

    \I__5313\ : Span4Mux_v
    port map (
            O => \N__30101\,
            I => \N__30090\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30090\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__30095\,
            I => r0_15
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__30090\,
            I => r0_15
        );

    \I__5309\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30074\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30074\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30069\
        );

    \I__5306\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30069\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__30081\,
            I => \N__30055\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__30080\,
            I => \N__30051\
        );

    \I__5303\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30033\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__30074\,
            I => \N__30028\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__30028\
        );

    \I__5300\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30021\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30021\
        );

    \I__5298\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30021\
        );

    \I__5297\ : InMux
    port map (
            O => \N__30065\,
            I => \N__30012\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30064\,
            I => \N__30012\
        );

    \I__5295\ : InMux
    port map (
            O => \N__30063\,
            I => \N__30012\
        );

    \I__5294\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30012\
        );

    \I__5293\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30005\
        );

    \I__5292\ : InMux
    port map (
            O => \N__30060\,
            I => \N__30005\
        );

    \I__5291\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30005\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30058\,
            I => \N__29998\
        );

    \I__5289\ : InMux
    port map (
            O => \N__30055\,
            I => \N__29998\
        );

    \I__5288\ : InMux
    port map (
            O => \N__30054\,
            I => \N__29998\
        );

    \I__5287\ : InMux
    port map (
            O => \N__30051\,
            I => \N__29991\
        );

    \I__5286\ : InMux
    port map (
            O => \N__30050\,
            I => \N__29991\
        );

    \I__5285\ : InMux
    port map (
            O => \N__30049\,
            I => \N__29991\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__30048\,
            I => \N__29982\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30047\,
            I => \N__29977\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30046\,
            I => \N__29977\
        );

    \I__5281\ : InMux
    port map (
            O => \N__30045\,
            I => \N__29962\
        );

    \I__5280\ : InMux
    port map (
            O => \N__30044\,
            I => \N__29962\
        );

    \I__5279\ : InMux
    port map (
            O => \N__30043\,
            I => \N__29953\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30042\,
            I => \N__29953\
        );

    \I__5277\ : InMux
    port map (
            O => \N__30041\,
            I => \N__29953\
        );

    \I__5276\ : InMux
    port map (
            O => \N__30040\,
            I => \N__29953\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30039\,
            I => \N__29944\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30038\,
            I => \N__29944\
        );

    \I__5273\ : InMux
    port map (
            O => \N__30037\,
            I => \N__29944\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30036\,
            I => \N__29944\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30033\,
            I => \N__29935\
        );

    \I__5270\ : Span4Mux_v
    port map (
            O => \N__30028\,
            I => \N__29935\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__30021\,
            I => \N__29935\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__30012\,
            I => \N__29935\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__30005\,
            I => \N__29924\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__29998\,
            I => \N__29924\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__29991\,
            I => \N__29921\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29914\
        );

    \I__5263\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29914\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29914\
        );

    \I__5261\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29911\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29904\
        );

    \I__5259\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29904\
        );

    \I__5258\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29904\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__29977\,
            I => \N__29900\
        );

    \I__5256\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29895\
        );

    \I__5255\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29895\
        );

    \I__5254\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29888\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29888\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29888\
        );

    \I__5251\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29881\
        );

    \I__5250\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29876\
        );

    \I__5249\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29876\
        );

    \I__5248\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29871\
        );

    \I__5247\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29871\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__29962\,
            I => \N__29868\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__29953\,
            I => \N__29865\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29944\,
            I => \N__29860\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__29935\,
            I => \N__29860\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29856\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29845\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29845\
        );

    \I__5239\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29845\
        );

    \I__5238\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29845\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29845\
        );

    \I__5236\ : Sp12to4
    port map (
            O => \N__29924\,
            I => \N__29839\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__29921\,
            I => \N__29834\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__29914\,
            I => \N__29834\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29831\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__29904\,
            I => \N__29828\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29825\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__29900\,
            I => \N__29822\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29895\,
            I => \N__29819\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29816\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29811\
        );

    \I__5226\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29811\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29806\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29806\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29797\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29797\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29797\
        );

    \I__5220\ : Span4Mux_v
    port map (
            O => \N__29868\,
            I => \N__29797\
        );

    \I__5219\ : Span4Mux_v
    port map (
            O => \N__29865\,
            I => \N__29792\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__29860\,
            I => \N__29792\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29789\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__29856\,
            I => \N__29784\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__29845\,
            I => \N__29784\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29844\,
            I => \N__29779\
        );

    \I__5213\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29779\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29776\
        );

    \I__5211\ : Span12Mux_h
    port map (
            O => \N__29839\,
            I => \N__29773\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__29834\,
            I => \N__29770\
        );

    \I__5209\ : Span4Mux_h
    port map (
            O => \N__29831\,
            I => \N__29763\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__29828\,
            I => \N__29763\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29763\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__29822\,
            I => \N__29756\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__29819\,
            I => \N__29756\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__29816\,
            I => \N__29756\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__29811\,
            I => \N__29747\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29747\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__29797\,
            I => \N__29747\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__29792\,
            I => \N__29747\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__29789\,
            I => \clkdivZ0Z_6\
        );

    \I__5198\ : Odrv12
    port map (
            O => \N__29784\,
            I => \clkdivZ0Z_6\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29779\,
            I => \clkdivZ0Z_6\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__29776\,
            I => \clkdivZ0Z_6\
        );

    \I__5195\ : Odrv12
    port map (
            O => \N__29773\,
            I => \clkdivZ0Z_6\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__29770\,
            I => \clkdivZ0Z_6\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__29763\,
            I => \clkdivZ0Z_6\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__29756\,
            I => \clkdivZ0Z_6\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__29747\,
            I => \clkdivZ0Z_6\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__29728\,
            I => \TXbuffer_18_3_ns_1_7_cascade_\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29722\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29718\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29715\
        );

    \I__5186\ : Span4Mux_v
    port map (
            O => \N__29718\,
            I => \N__29712\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29709\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__29712\,
            I => \N__29705\
        );

    \I__5183\ : Span4Mux_s2_h
    port map (
            O => \N__29709\,
            I => \N__29702\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29699\
        );

    \I__5181\ : Sp12to4
    port map (
            O => \N__29705\,
            I => \N__29696\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__29702\,
            I => \N__29693\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__29699\,
            I => \N__29690\
        );

    \I__5178\ : Odrv12
    port map (
            O => \N__29696\,
            I => r4_15
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__29693\,
            I => r4_15
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__29690\,
            I => r4_15
        );

    \I__5175\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29680\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__29677\,
            I => \N__29671\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29665\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29662\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__29674\,
            I => \N__29658\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__29671\,
            I => \N__29655\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29670\,
            I => \N__29652\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29669\,
            I => \N__29649\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29668\,
            I => \N__29646\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29643\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__29662\,
            I => \N__29640\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29637\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29634\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__29655\,
            I => \N__29629\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__29652\,
            I => \N__29629\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29649\,
            I => \N__29626\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__29646\,
            I => \N__29623\
        );

    \I__5157\ : Span12Mux_h
    port map (
            O => \N__29643\,
            I => \N__29619\
        );

    \I__5156\ : Span12Mux_v
    port map (
            O => \N__29640\,
            I => \N__29616\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29609\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29609\
        );

    \I__5153\ : Span4Mux_v
    port map (
            O => \N__29629\,
            I => \N__29609\
        );

    \I__5152\ : Span4Mux_h
    port map (
            O => \N__29626\,
            I => \N__29606\
        );

    \I__5151\ : Span4Mux_h
    port map (
            O => \N__29623\,
            I => \N__29603\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29600\
        );

    \I__5149\ : Odrv12
    port map (
            O => \N__29619\,
            I => \clkdivZ0Z_5\
        );

    \I__5148\ : Odrv12
    port map (
            O => \N__29616\,
            I => \clkdivZ0Z_5\
        );

    \I__5147\ : Odrv4
    port map (
            O => \N__29609\,
            I => \clkdivZ0Z_5\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__29606\,
            I => \clkdivZ0Z_5\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__29603\,
            I => \clkdivZ0Z_5\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29600\,
            I => \clkdivZ0Z_5\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__29587\,
            I => \TXbuffer_RNO_5Z0Z_7_cascade_\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29581\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29578\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__29578\,
            I => \N__29575\
        );

    \I__5139\ : Span4Mux_v
    port map (
            O => \N__29575\,
            I => \N__29572\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__29572\,
            I => \N__29569\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__29569\,
            I => \TXbuffer_RNO_6Z0Z_7\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__29566\,
            I => \ALU.a_3_ns_1_1_cascade_\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__29563\,
            I => \N__29559\
        );

    \I__5134\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29556\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29553\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29550\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29547\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__29550\,
            I => \N__29544\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__29547\,
            I => \ALU.a3_b_2\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__29544\,
            I => \ALU.a3_b_2\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__29539\,
            I => \ALU.rshift_3_ns_1_7_cascade_\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__29536\,
            I => \ALU.b_3_ns_1_7_cascade_\
        );

    \I__5125\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29530\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__29530\,
            I => \N__29527\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__29527\,
            I => \N__29524\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__29524\,
            I => \N__29521\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__29521\,
            I => \ALU.r4_RNI82OE1Z0Z_7\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29509\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29509\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__29516\,
            I => \N__29504\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29499\
        );

    \I__5116\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29499\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29509\,
            I => \N__29496\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29493\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29490\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29483\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__29499\,
            I => \N__29476\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__29496\,
            I => \N__29476\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__29493\,
            I => \N__29471\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__29490\,
            I => \N__29471\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29462\
        );

    \I__5106\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29462\
        );

    \I__5105\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29462\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29462\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29483\,
            I => \N__29459\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29454\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29454\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__29476\,
            I => \N__29451\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__29471\,
            I => \b_0_repZ0Z2\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__29462\,
            I => \b_0_repZ0Z2\
        );

    \I__5097\ : Odrv12
    port map (
            O => \N__29459\,
            I => \b_0_repZ0Z2\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__29454\,
            I => \b_0_repZ0Z2\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__29451\,
            I => \b_0_repZ0Z2\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29436\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29439\,
            I => \N__29433\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29436\,
            I => \N__29430\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__29433\,
            I => \N__29426\
        );

    \I__5090\ : Span4Mux_h
    port map (
            O => \N__29430\,
            I => \N__29423\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29429\,
            I => \N__29420\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__29426\,
            I => \N__29417\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__29423\,
            I => \N__29414\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29420\,
            I => r7_1
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__29417\,
            I => r7_1
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__29414\,
            I => r7_1
        );

    \I__5083\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29403\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29400\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__29403\,
            I => \N__29397\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29400\,
            I => \N__29393\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__29397\,
            I => \N__29390\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29396\,
            I => \N__29387\
        );

    \I__5077\ : Span12Mux_v
    port map (
            O => \N__29393\,
            I => \N__29384\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__29390\,
            I => \N__29381\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__29387\,
            I => r6_1
        );

    \I__5074\ : Odrv12
    port map (
            O => \N__29384\,
            I => r6_1
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__29381\,
            I => r6_1
        );

    \I__5072\ : InMux
    port map (
            O => \N__29374\,
            I => \N__29371\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__5070\ : Odrv12
    port map (
            O => \N__29368\,
            I => \ALU.r6_RNIC9P41Z0Z_1\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29361\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29356\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29361\,
            I => \N__29353\
        );

    \I__5066\ : InMux
    port map (
            O => \N__29360\,
            I => \N__29350\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29359\,
            I => \N__29347\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__29356\,
            I => \N__29344\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__29353\,
            I => \N__29339\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29350\,
            I => \N__29339\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__29347\,
            I => \ALU.r6_RNIE5FT1Z0Z_2\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__29344\,
            I => \ALU.r6_RNIE5FT1Z0Z_2\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__29339\,
            I => \ALU.r6_RNIE5FT1Z0Z_2\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29332\,
            I => \N__29326\
        );

    \I__5057\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29326\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29326\,
            I => \N__29323\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__29323\,
            I => \ALU.madd_13\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__29320\,
            I => \N__29316\
        );

    \I__5053\ : CascadeMux
    port map (
            O => \N__29319\,
            I => \N__29313\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29310\
        );

    \I__5051\ : InMux
    port map (
            O => \N__29313\,
            I => \N__29307\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__29310\,
            I => \N__29304\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__29307\,
            I => \ALU.a2_b_0\
        );

    \I__5048\ : Odrv12
    port map (
            O => \N__29304\,
            I => \ALU.a2_b_0\
        );

    \I__5047\ : CascadeMux
    port map (
            O => \N__29299\,
            I => \N__29296\
        );

    \I__5046\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29293\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__29293\,
            I => \ALU.madd_3\
        );

    \I__5044\ : InMux
    port map (
            O => \N__29290\,
            I => \N__29284\
        );

    \I__5043\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29284\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__29284\,
            I => \N__29281\
        );

    \I__5041\ : Odrv12
    port map (
            O => \N__29281\,
            I => \ALU.madd_4\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__29278\,
            I => \ALU.madd_3_cascade_\
        );

    \I__5039\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29269\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29269\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__29269\,
            I => \ALU.a0_b_3\
        );

    \I__5036\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29259\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29256\
        );

    \I__5033\ : Span4Mux_s2_v
    port map (
            O => \N__29259\,
            I => \N__29251\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29251\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__29251\,
            I => \N__29248\
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__29248\,
            I => \ALU.madd_66\
        );

    \I__5029\ : CascadeMux
    port map (
            O => \N__29245\,
            I => \N__29241\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__29244\,
            I => \N__29238\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29234\
        );

    \I__5026\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29231\
        );

    \I__5025\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29228\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__29234\,
            I => \N__29221\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29221\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__29228\,
            I => \N__29216\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__29227\,
            I => \N__29212\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__29226\,
            I => \N__29209\
        );

    \I__5019\ : Span4Mux_v
    port map (
            O => \N__29221\,
            I => \N__29203\
        );

    \I__5018\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29199\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29196\
        );

    \I__5016\ : Span4Mux_s3_v
    port map (
            O => \N__29216\,
            I => \N__29193\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29190\
        );

    \I__5014\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29187\
        );

    \I__5013\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29184\
        );

    \I__5012\ : CascadeMux
    port map (
            O => \N__29208\,
            I => \N__29180\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29177\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29174\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__29203\,
            I => \N__29171\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29168\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__29199\,
            I => \N__29161\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__29196\,
            I => \N__29161\
        );

    \I__5005\ : Span4Mux_h
    port map (
            O => \N__29193\,
            I => \N__29161\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__29190\,
            I => \N__29157\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__29187\,
            I => \N__29151\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__29184\,
            I => \N__29151\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29183\,
            I => \N__29146\
        );

    \I__5000\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29146\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29141\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29141\
        );

    \I__4997\ : Sp12to4
    port map (
            O => \N__29171\,
            I => \N__29136\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29168\,
            I => \N__29136\
        );

    \I__4995\ : Sp12to4
    port map (
            O => \N__29161\,
            I => \N__29133\
        );

    \I__4994\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29130\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__29157\,
            I => \N__29127\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29124\
        );

    \I__4991\ : Span12Mux_s5_h
    port map (
            O => \N__29151\,
            I => \N__29119\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29119\
        );

    \I__4989\ : Span12Mux_v
    port map (
            O => \N__29141\,
            I => \N__29112\
        );

    \I__4988\ : Span12Mux_s4_h
    port map (
            O => \N__29136\,
            I => \N__29112\
        );

    \I__4987\ : Span12Mux_s8_v
    port map (
            O => \N__29133\,
            I => \N__29112\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__29130\,
            I => \a_1_repZ0Z1\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__29127\,
            I => \a_1_repZ0Z1\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__29124\,
            I => \a_1_repZ0Z1\
        );

    \I__4983\ : Odrv12
    port map (
            O => \N__29119\,
            I => \a_1_repZ0Z1\
        );

    \I__4982\ : Odrv12
    port map (
            O => \N__29112\,
            I => \a_1_repZ0Z1\
        );

    \I__4981\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29097\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29091\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29097\,
            I => \N__29088\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29081\
        );

    \I__4977\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29081\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29081\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__29091\,
            I => \N__29073\
        );

    \I__4974\ : Span4Mux_s2_v
    port map (
            O => \N__29088\,
            I => \N__29068\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__29081\,
            I => \N__29068\
        );

    \I__4972\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29065\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29062\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29078\,
            I => \N__29059\
        );

    \I__4969\ : InMux
    port map (
            O => \N__29077\,
            I => \N__29056\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29076\,
            I => \N__29053\
        );

    \I__4967\ : Span4Mux_s2_v
    port map (
            O => \N__29073\,
            I => \N__29048\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__29068\,
            I => \N__29048\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29045\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__29062\,
            I => \N__29040\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29059\,
            I => \N__29040\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__29056\,
            I => \N__29037\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__29053\,
            I => \N__29034\
        );

    \I__4960\ : Span4Mux_v
    port map (
            O => \N__29048\,
            I => \N__29031\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__29045\,
            I => \N__29026\
        );

    \I__4958\ : Span4Mux_s3_v
    port map (
            O => \N__29040\,
            I => \N__29026\
        );

    \I__4957\ : Sp12to4
    port map (
            O => \N__29037\,
            I => \N__29021\
        );

    \I__4956\ : Span12Mux_s7_v
    port map (
            O => \N__29034\,
            I => \N__29021\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__29031\,
            I => \ALU.r6_RNIASIB2Z0Z_5\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__29026\,
            I => \ALU.r6_RNIASIB2Z0Z_5\
        );

    \I__4953\ : Odrv12
    port map (
            O => \N__29021\,
            I => \ALU.r6_RNIASIB2Z0Z_5\
        );

    \I__4952\ : CascadeMux
    port map (
            O => \N__29014\,
            I => \N__29010\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29013\,
            I => \N__29006\
        );

    \I__4950\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29000\
        );

    \I__4949\ : InMux
    port map (
            O => \N__29009\,
            I => \N__28994\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__29006\,
            I => \N__28991\
        );

    \I__4947\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28988\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28985\
        );

    \I__4945\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28982\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29000\,
            I => \N__28979\
        );

    \I__4943\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28971\
        );

    \I__4942\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28971\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28971\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__28994\,
            I => \N__28968\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__28991\,
            I => \N__28963\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28963\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28960\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28957\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__28979\,
            I => \N__28954\
        );

    \I__4934\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28951\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28946\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__28968\,
            I => \N__28946\
        );

    \I__4931\ : Span4Mux_s1_v
    port map (
            O => \N__28963\,
            I => \N__28943\
        );

    \I__4930\ : Span4Mux_v
    port map (
            O => \N__28960\,
            I => \N__28940\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__28957\,
            I => \N__28935\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__28954\,
            I => \N__28935\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28930\
        );

    \I__4926\ : Sp12to4
    port map (
            O => \N__28946\,
            I => \N__28930\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__28943\,
            I => \N__28925\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__28940\,
            I => \N__28925\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__28935\,
            I => \ALU.r4_RNI24Q22Z0Z_5\
        );

    \I__4922\ : Odrv12
    port map (
            O => \N__28930\,
            I => \ALU.r4_RNI24Q22Z0Z_5\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__28925\,
            I => \ALU.r4_RNI24Q22Z0Z_5\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28909\
        );

    \I__4919\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28909\
        );

    \I__4918\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28909\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__28909\,
            I => \ALU.a0_b_4\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28903\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__28903\,
            I => \N__28900\
        );

    \I__4914\ : Span4Mux_s3_v
    port map (
            O => \N__28900\,
            I => \N__28897\
        );

    \I__4913\ : Odrv4
    port map (
            O => \N__28897\,
            I => \ALU.un2_addsub_axb_2\
        );

    \I__4912\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28887\
        );

    \I__4911\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28887\
        );

    \I__4910\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28884\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28881\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__28884\,
            I => \ALU.madd_56\
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__28881\,
            I => \ALU.madd_56\
        );

    \I__4906\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28870\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__28870\,
            I => \N__28865\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28869\,
            I => \N__28860\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28860\
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__28865\,
            I => \ALU.madd_45\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__28860\,
            I => \ALU.madd_45\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__28855\,
            I => \N__28852\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28849\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__4896\ : Span4Mux_h
    port map (
            O => \N__28846\,
            I => \N__28843\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__28843\,
            I => \ALU.madd_cry_6_ma\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28835\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__28839\,
            I => \N__28832\
        );

    \I__4892\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28829\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28826\
        );

    \I__4890\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28823\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__28829\,
            I => \N__28820\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__28826\,
            I => \N__28817\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28814\
        );

    \I__4886\ : Span4Mux_s3_h
    port map (
            O => \N__28820\,
            I => \N__28811\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__28817\,
            I => \N__28808\
        );

    \I__4884\ : Span4Mux_h
    port map (
            O => \N__28814\,
            I => \N__28805\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__28811\,
            I => r3_0
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__28808\,
            I => r3_0
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__28805\,
            I => r3_0
        );

    \I__4880\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28795\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28792\
        );

    \I__4878\ : Span4Mux_v
    port map (
            O => \N__28792\,
            I => \N__28785\
        );

    \I__4877\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28772\
        );

    \I__4876\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28772\
        );

    \I__4875\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28772\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28788\,
            I => \N__28772\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__28785\,
            I => \N__28769\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28760\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28760\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28760\
        );

    \I__4869\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28760\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28772\,
            I => \a_0_repZ0Z2\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__28769\,
            I => \a_0_repZ0Z2\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__28760\,
            I => \a_0_repZ0Z2\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__4863\ : Span4Mux_s3_v
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__28744\,
            I => \ALU.r2_RNI18BOZ0Z_0\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28737\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28734\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__28737\,
            I => \N__28731\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28734\,
            I => \N__28728\
        );

    \I__4857\ : Sp12to4
    port map (
            O => \N__28731\,
            I => \N__28725\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__28728\,
            I => \N__28721\
        );

    \I__4855\ : Span12Mux_v
    port map (
            O => \N__28725\,
            I => \N__28718\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28715\
        );

    \I__4853\ : Span4Mux_h
    port map (
            O => \N__28721\,
            I => \N__28712\
        );

    \I__4852\ : Odrv12
    port map (
            O => \N__28718\,
            I => r2_0
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__28715\,
            I => r2_0
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__28712\,
            I => r2_0
        );

    \I__4849\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28702\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__28702\,
            I => \N__28697\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28694\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__28700\,
            I => \N__28691\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__28697\,
            I => \N__28688\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__28694\,
            I => \N__28685\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28682\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__28688\,
            I => \N__28679\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__28685\,
            I => \N__28676\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28673\
        );

    \I__4839\ : Span4Mux_v
    port map (
            O => \N__28679\,
            I => \N__28670\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__28676\,
            I => r3_1
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__28673\,
            I => r3_1
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__28670\,
            I => r3_1
        );

    \I__4835\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28659\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28656\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28659\,
            I => \N__28653\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__28656\,
            I => \N__28649\
        );

    \I__4831\ : Span12Mux_h
    port map (
            O => \N__28653\,
            I => \N__28646\
        );

    \I__4830\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28643\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__28649\,
            I => r2_1
        );

    \I__4828\ : Odrv12
    port map (
            O => \N__28646\,
            I => r2_1
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__28643\,
            I => r2_1
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__28636\,
            I => \N__28633\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__28630\,
            I => \N__28627\
        );

    \I__4823\ : Sp12to4
    port map (
            O => \N__28627\,
            I => \N__28624\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__28624\,
            I => \ALU.r2_RNI4H0SZ0Z_1\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28614\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28611\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__28614\,
            I => \ALU.madd_29_0\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28611\,
            I => \ALU.madd_29_0\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28603\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__28600\,
            I => \ALU.madd_18\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28594\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__28594\,
            I => \N__28590\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28587\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__28590\,
            I => \ALU.madd_34\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28587\,
            I => \ALU.madd_34\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__28582\,
            I => \ALU.madd_39_cascade_\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28576\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__28576\,
            I => \ALU.madd_39\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__28573\,
            I => \ALU.madd_23_cascade_\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28567\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__28567\,
            I => \N__28564\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__28564\,
            I => \N__28560\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28557\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__28560\,
            I => \ALU.madd_28\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28557\,
            I => \ALU.madd_28\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__28552\,
            I => \N__28549\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28543\
        );

    \I__4795\ : Span4Mux_v
    port map (
            O => \N__28543\,
            I => \N__28540\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__28540\,
            I => \ALU.madd_axb_4_l_fx\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28528\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28528\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28535\,
            I => \N__28528\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28528\,
            I => \ALU.madd_8\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28519\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28519\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28516\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__28516\,
            I => \N__28513\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28513\,
            I => \ALU.madd_19\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28507\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28507\,
            I => \N__28504\
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__28504\,
            I => \TXbuffer_RNO_1Z0Z_5\
        );

    \I__4781\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28498\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__28498\,
            I => \N__28495\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__28495\,
            I => \TXbuffer_RNO_0Z0Z_5\
        );

    \I__4778\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__28486\,
            I => \TXbuffer_18_15_ns_1_5\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__28483\,
            I => \ALU.a2_b_1_cascade_\
        );

    \I__4774\ : InMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__28477\,
            I => \ALU.a1_b_2\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28471\,
            I => \ALU.a2_b_1\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__28468\,
            I => \ALU.a1_b_2_cascade_\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28462\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__28462\,
            I => \ALU.r0_12_prm_3_12_s0_sf\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28456\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28456\,
            I => \N__28453\
        );

    \I__4765\ : Odrv12
    port map (
            O => \N__28453\,
            I => \ALU.mult_12\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28450\,
            I => \ALU.r0_12_s0_12\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__28447\,
            I => \N__28443\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28437\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28434\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28442\,
            I => \N__28431\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28428\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28424\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28420\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28415\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28431\,
            I => \N__28415\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__28428\,
            I => \N__28412\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28409\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28406\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28403\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__28420\,
            I => \N__28397\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__28415\,
            I => \N__28397\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__28412\,
            I => \N__28392\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__28409\,
            I => \N__28392\
        );

    \I__4746\ : Span4Mux_v
    port map (
            O => \N__28406\,
            I => \N__28387\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28403\,
            I => \N__28387\
        );

    \I__4744\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28384\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__28397\,
            I => \ALU.r0_12_12\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__28392\,
            I => \ALU.r0_12_12\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__28387\,
            I => \ALU.r0_12_12\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28384\,
            I => \ALU.r0_12_12\
        );

    \I__4739\ : InMux
    port map (
            O => \N__28375\,
            I => \N__28370\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28367\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28364\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__28370\,
            I => \N__28361\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__28367\,
            I => \N__28358\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__28364\,
            I => \N__28355\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__28361\,
            I => \N__28352\
        );

    \I__4732\ : Span4Mux_h
    port map (
            O => \N__28358\,
            I => \N__28349\
        );

    \I__4731\ : Span4Mux_h
    port map (
            O => \N__28355\,
            I => \N__28346\
        );

    \I__4730\ : Span4Mux_v
    port map (
            O => \N__28352\,
            I => \N__28343\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__28349\,
            I => r0_12
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__28346\,
            I => r0_12
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__28343\,
            I => r0_12
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__4725\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28330\,
            I => \ALU.r0_12_prm_3_14_s0_sf\
        );

    \I__4723\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28324\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__28324\,
            I => \N__28321\
        );

    \I__4721\ : Span4Mux_v
    port map (
            O => \N__28321\,
            I => \N__28318\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__28318\,
            I => \ALU.mult_14\
        );

    \I__4719\ : InMux
    port map (
            O => \N__28315\,
            I => \ALU.r0_12_s0_14\
        );

    \I__4718\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28305\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28302\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28299\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28296\
        );

    \I__4714\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28290\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__28305\,
            I => \N__28287\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__28302\,
            I => \N__28284\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__28299\,
            I => \N__28279\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28279\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28276\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28273\
        );

    \I__4707\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28270\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28267\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__28287\,
            I => \N__28264\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__28284\,
            I => \N__28259\
        );

    \I__4703\ : Span4Mux_v
    port map (
            O => \N__28279\,
            I => \N__28259\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__28276\,
            I => \ALU.r0_12_14\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28273\,
            I => \ALU.r0_12_14\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__28270\,
            I => \ALU.r0_12_14\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__28267\,
            I => \ALU.r0_12_14\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__28264\,
            I => \ALU.r0_12_14\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__28259\,
            I => \ALU.r0_12_14\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28242\
        );

    \I__4695\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28239\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__28242\,
            I => \N__28235\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28239\,
            I => \N__28232\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__28238\,
            I => \N__28229\
        );

    \I__4691\ : Span4Mux_h
    port map (
            O => \N__28235\,
            I => \N__28226\
        );

    \I__4690\ : Span4Mux_h
    port map (
            O => \N__28232\,
            I => \N__28223\
        );

    \I__4689\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28220\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__28226\,
            I => r1_14
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__28223\,
            I => r1_14
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__28220\,
            I => r1_14
        );

    \I__4685\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__28210\,
            I => \ALU.r0_12_prm_3_10_s0_sf\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28201\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__28201\,
            I => \N__28198\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__28198\,
            I => \ALU.mult_10\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28195\,
            I => \ALU.r0_12_s0_10\
        );

    \I__4678\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28186\
        );

    \I__4677\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28183\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28180\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28177\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__28186\,
            I => \N__28173\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28170\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28167\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__28177\,
            I => \N__28164\
        );

    \I__4670\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28161\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__28173\,
            I => \N__28153\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__28170\,
            I => \N__28153\
        );

    \I__4667\ : Span4Mux_v
    port map (
            O => \N__28167\,
            I => \N__28148\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__28164\,
            I => \N__28148\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28145\
        );

    \I__4664\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28142\
        );

    \I__4663\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28139\
        );

    \I__4662\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28136\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__28153\,
            I => \ALU.r0_12_10\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__28148\,
            I => \ALU.r0_12_10\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__28145\,
            I => \ALU.r0_12_10\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28142\,
            I => \ALU.r0_12_10\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__28139\,
            I => \ALU.r0_12_10\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__28136\,
            I => \ALU.r0_12_10\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28118\
        );

    \I__4654\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28115\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28112\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__28118\,
            I => \N__28109\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__28115\,
            I => \N__28106\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__28112\,
            I => \N__28103\
        );

    \I__4649\ : Span4Mux_h
    port map (
            O => \N__28109\,
            I => \N__28100\
        );

    \I__4648\ : Span12Mux_s6_h
    port map (
            O => \N__28106\,
            I => \N__28097\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__28103\,
            I => r0_10
        );

    \I__4646\ : Odrv4
    port map (
            O => \N__28100\,
            I => r0_10
        );

    \I__4645\ : Odrv12
    port map (
            O => \N__28097\,
            I => r0_10
        );

    \I__4644\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28083\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28083\
        );

    \I__4642\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28080\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28077\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__28080\,
            I => \N__28074\
        );

    \I__4639\ : Span4Mux_s3_h
    port map (
            O => \N__28077\,
            I => \N__28071\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__28074\,
            I => \N__28068\
        );

    \I__4637\ : Span4Mux_h
    port map (
            O => \N__28071\,
            I => \N__28065\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__28068\,
            I => r7_2
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__28065\,
            I => r7_2
        );

    \I__4634\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28056\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28053\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__28056\,
            I => \N__28050\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28047\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__28050\,
            I => \N__28041\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__28047\,
            I => \N__28041\
        );

    \I__4628\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28038\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__28041\,
            I => \N__28035\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28038\,
            I => \N__28032\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__28035\,
            I => r7_3
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__28032\,
            I => r7_3
        );

    \I__4623\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28024\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__28024\,
            I => \N__28021\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__28021\,
            I => \N__28018\
        );

    \I__4620\ : Span4Mux_h
    port map (
            O => \N__28018\,
            I => \N__28013\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28017\,
            I => \N__28008\
        );

    \I__4618\ : InMux
    port map (
            O => \N__28016\,
            I => \N__28008\
        );

    \I__4617\ : Span4Mux_v
    port map (
            O => \N__28013\,
            I => \N__28003\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__28003\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__28003\,
            I => r7_4
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__28000\,
            I => \TXbuffer_18_10_ns_1_1_cascade_\
        );

    \I__4613\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27994\,
            I => \N__27991\
        );

    \I__4611\ : Sp12to4
    port map (
            O => \N__27991\,
            I => \N__27988\
        );

    \I__4610\ : Span12Mux_v
    port map (
            O => \N__27988\,
            I => \N__27985\
        );

    \I__4609\ : Odrv12
    port map (
            O => \N__27985\,
            I => \TXbuffer_18_15_ns_1_1\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__27982\,
            I => \TXbuffer_RNO_0Z0Z_1_cascade_\
        );

    \I__4607\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27976\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__27976\,
            I => \TXbuffer_RNO_1Z0Z_1\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__27973\,
            I => \N__27969\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27966\
        );

    \I__4603\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27963\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N__27959\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__27963\,
            I => \N__27956\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__27962\,
            I => \N__27953\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__27959\,
            I => \N__27950\
        );

    \I__4598\ : Span4Mux_h
    port map (
            O => \N__27956\,
            I => \N__27947\
        );

    \I__4597\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27944\
        );

    \I__4596\ : Odrv4
    port map (
            O => \N__27950\,
            I => r1_10
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__27947\,
            I => r1_10
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__27944\,
            I => r1_10
        );

    \I__4593\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27933\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27929\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__27933\,
            I => \N__27926\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27923\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27920\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__27926\,
            I => \N__27917\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27914\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__27920\,
            I => \N__27911\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__27917\,
            I => \N__27908\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__27914\,
            I => \N__27905\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__27911\,
            I => r5_10
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__27908\,
            I => r5_10
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__27905\,
            I => r5_10
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__27898\,
            I => \TXbuffer_18_10_ns_1_2_cascade_\
        );

    \I__4579\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27892\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__27892\,
            I => \N__27889\
        );

    \I__4577\ : Span4Mux_v
    port map (
            O => \N__27889\,
            I => \N__27886\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__27886\,
            I => \TXbuffer_RNO_0Z0Z_2\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27879\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27875\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__27879\,
            I => \N__27872\
        );

    \I__4572\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27869\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__27875\,
            I => \N__27866\
        );

    \I__4570\ : Span4Mux_h
    port map (
            O => \N__27872\,
            I => \N__27863\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__27869\,
            I => \N__27860\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__27866\,
            I => \N__27853\
        );

    \I__4567\ : Span4Mux_v
    port map (
            O => \N__27863\,
            I => \N__27853\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__27860\,
            I => \N__27853\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__27853\,
            I => r7_6
        );

    \I__4564\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27847\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__27847\,
            I => \N__27844\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__27844\,
            I => \N__27839\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27834\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27834\
        );

    \I__4559\ : Sp12to4
    port map (
            O => \N__27839\,
            I => \N__27829\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27829\
        );

    \I__4557\ : Odrv12
    port map (
            O => \N__27829\,
            I => r7_7
        );

    \I__4556\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27821\
        );

    \I__4555\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27816\
        );

    \I__4554\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27816\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__27821\,
            I => \N__27813\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__27816\,
            I => \N__27810\
        );

    \I__4551\ : Span12Mux_s6_h
    port map (
            O => \N__27813\,
            I => \N__27807\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__27810\,
            I => \N__27804\
        );

    \I__4549\ : Odrv12
    port map (
            O => \N__27807\,
            I => r7_8
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__27804\,
            I => r7_8
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__4546\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27792\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27789\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__27792\,
            I => \N__27786\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27782\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__27786\,
            I => \N__27779\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27776\
        );

    \I__4540\ : Span4Mux_h
    port map (
            O => \N__27782\,
            I => \N__27773\
        );

    \I__4539\ : Span4Mux_s3_h
    port map (
            O => \N__27779\,
            I => \N__27770\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__27776\,
            I => r7_9
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__27773\,
            I => r7_9
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__27770\,
            I => r7_9
        );

    \I__4535\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27760\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__27760\,
            I => \ALU.r4_RNIJJH11Z0Z_0\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__27757\,
            I => \ALU.r0_RNIBROOZ0Z_0_cascade_\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27745\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27745\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27742\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27735\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27735\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27745\,
            I => \N__27729\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27729\
        );

    \I__4525\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27724\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27724\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27721\
        );

    \I__4522\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27717\
        );

    \I__4521\ : Span4Mux_v
    port map (
            O => \N__27729\,
            I => \N__27710\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27710\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__27721\,
            I => \N__27710\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27707\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27717\,
            I => \a_fastZ0Z_1\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__27710\,
            I => \a_fastZ0Z_1\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__27707\,
            I => \a_fastZ0Z_1\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27697\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__4512\ : Span4Mux_s2_v
    port map (
            O => \N__27694\,
            I => \N__27691\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__27691\,
            I => \N__27688\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__27688\,
            I => \ALU.a_7_ns_1_0\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27682\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__27682\,
            I => \N__27677\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27672\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27672\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__27677\,
            I => \N__27669\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__27672\,
            I => \N__27666\
        );

    \I__4503\ : Span4Mux_v
    port map (
            O => \N__27669\,
            I => \N__27661\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__27666\,
            I => \N__27661\
        );

    \I__4501\ : Odrv4
    port map (
            O => \N__27661\,
            I => r4_0
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \TXbuffer_18_3_ns_1_0_cascade_\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27649\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__27649\,
            I => \N__27646\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__27646\,
            I => \N__27643\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__27643\,
            I => \TXbuffer_RNO_5Z0Z_0\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__27640\,
            I => \TXbuffer_18_10_ns_1_0_cascade_\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__27637\,
            I => \N__27634\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27631\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__27631\,
            I => \N__27626\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27621\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27621\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__27626\,
            I => \N__27618\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27615\
        );

    \I__4486\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27610\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__27615\,
            I => \N__27610\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__27610\,
            I => r5_0
        );

    \I__4483\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27604\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27601\
        );

    \I__4481\ : Span4Mux_s2_h
    port map (
            O => \N__27601\,
            I => \N__27598\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__27598\,
            I => \N__27595\
        );

    \I__4479\ : Sp12to4
    port map (
            O => \N__27595\,
            I => \N__27592\
        );

    \I__4478\ : Odrv12
    port map (
            O => \N__27592\,
            I => \TXbuffer_RNO_0Z0Z_0\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27585\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__27588\,
            I => \N__27582\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27585\,
            I => \N__27578\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27582\,
            I => \N__27575\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27581\,
            I => \N__27572\
        );

    \I__4472\ : Span4Mux_v
    port map (
            O => \N__27578\,
            I => \N__27567\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__27575\,
            I => \N__27567\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27562\
        );

    \I__4469\ : Span4Mux_h
    port map (
            O => \N__27567\,
            I => \N__27562\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__27562\,
            I => r3_9
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__27559\,
            I => \N__27556\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27553\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__27553\,
            I => \TXbuffer_18_13_ns_1_1\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__27550\,
            I => \N__27547\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27544\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27541\
        );

    \I__4461\ : Odrv12
    port map (
            O => \N__27541\,
            I => \ALU.madd_cry_9_ma\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27538\,
            I => \ALU.madd_cry_8\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__27535\,
            I => \N__27531\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27528\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27525\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27522\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27525\,
            I => \N__27519\
        );

    \I__4454\ : Span12Mux_h
    port map (
            O => \N__27522\,
            I => \N__27516\
        );

    \I__4453\ : Span12Mux_v
    port map (
            O => \N__27519\,
            I => \N__27513\
        );

    \I__4452\ : Odrv12
    port map (
            O => \N__27516\,
            I => \ALU.madd_axb_10\
        );

    \I__4451\ : Odrv12
    port map (
            O => \N__27513\,
            I => \ALU.madd_axb_10\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__27508\,
            I => \N__27505\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27502\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27502\,
            I => \N__27499\
        );

    \I__4447\ : Span4Mux_v
    port map (
            O => \N__27499\,
            I => \N__27496\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__27496\,
            I => \N__27493\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__27493\,
            I => \ALU.madd_cry_9_THRU_CO\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27490\,
            I => \ALU.madd_cry_9\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27484\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__27484\,
            I => \N__27481\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__27481\,
            I => \N__27477\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27474\
        );

    \I__4439\ : Span4Mux_h
    port map (
            O => \N__27477\,
            I => \N__27471\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27468\
        );

    \I__4437\ : Span4Mux_v
    port map (
            O => \N__27471\,
            I => \N__27465\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__27468\,
            I => \ALU.g0_13\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__27465\,
            I => \ALU.g0_13\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__27460\,
            I => \N__27457\
        );

    \I__4433\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27454\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27451\
        );

    \I__4431\ : Span4Mux_v
    port map (
            O => \N__27451\,
            I => \N__27448\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__27448\,
            I => \ALU.madd_axb_11_l_fx\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27445\,
            I => \ALU.madd_cry_10\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27439\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__27439\,
            I => \N__27436\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__27436\,
            I => \N__27433\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__27433\,
            I => \ALU.madd_cry_12_ma\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__27430\,
            I => \N__27427\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27424\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27424\,
            I => \N__27421\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__27418\,
            I => \N__27415\
        );

    \I__4419\ : Odrv4
    port map (
            O => \N__27415\,
            I => \ALU.madd_axb_12_l_ofx\
        );

    \I__4418\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27409\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__27409\,
            I => \N__27406\
        );

    \I__4416\ : Span4Mux_v
    port map (
            O => \N__27406\,
            I => \N__27403\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__27403\,
            I => \N__27400\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__27400\,
            I => \ALU.mult_13\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27397\,
            I => \ALU.madd_cry_11\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27391\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__27388\,
            I => \N__27385\
        );

    \I__4409\ : Span4Mux_s3_h
    port map (
            O => \N__27385\,
            I => \N__27382\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__27382\,
            I => \ALU.madd_axb_13_l_ofx\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__27379\,
            I => \N__27376\
        );

    \I__4406\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27373\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27373\,
            I => \N__27370\
        );

    \I__4404\ : Span4Mux_h
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__27367\,
            I => \ALU.madd_cry_13_ma\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27364\,
            I => \ALU.madd_cry_12\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27361\,
            I => \ALU.madd_cry_13\
        );

    \I__4400\ : CascadeMux
    port map (
            O => \N__27358\,
            I => \N__27355\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27352\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27352\,
            I => \N__27349\
        );

    \I__4397\ : Span12Mux_v
    port map (
            O => \N__27349\,
            I => \N__27346\
        );

    \I__4396\ : Odrv12
    port map (
            O => \N__27346\,
            I => \ALU.madd_cry_13_THRU_CO\
        );

    \I__4395\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27338\
        );

    \I__4394\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27333\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27333\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__27338\,
            I => \ALU.a13_b_1\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__27333\,
            I => \ALU.a13_b_1\
        );

    \I__4390\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27325\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27322\
        );

    \I__4388\ : Span4Mux_v
    port map (
            O => \N__27322\,
            I => \N__27319\
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__27319\,
            I => \ALU.madd_373_0\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__27316\,
            I => \N__27313\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27310\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__27310\,
            I => \ALU.madd_368_0\
        );

    \I__4383\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27303\
        );

    \I__4382\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27300\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__27303\,
            I => \N__27297\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__27300\,
            I => \N__27294\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__27297\,
            I => \N__27291\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__27294\,
            I => \N__27288\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__27291\,
            I => \N__27285\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__27288\,
            I => \ALU.a9_b_5\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__27285\,
            I => \ALU.a9_b_5\
        );

    \I__4374\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27274\
        );

    \I__4373\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27274\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__27274\,
            I => \N__27271\
        );

    \I__4371\ : Odrv12
    port map (
            O => \N__27271\,
            I => \ALU.madd_398_0\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27268\,
            I => \ALU.madd_cry_0\
        );

    \I__4369\ : InMux
    port map (
            O => \N__27265\,
            I => \ALU.madd_cry_1\
        );

    \I__4368\ : InMux
    port map (
            O => \N__27262\,
            I => \ALU.madd_cry_2\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27259\,
            I => \ALU.madd_cry_3\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__4365\ : InMux
    port map (
            O => \N__27253\,
            I => \N__27250\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27250\,
            I => \N__27247\
        );

    \I__4363\ : Odrv12
    port map (
            O => \N__27247\,
            I => \ALU.madd_axb_5_l_fx\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27244\,
            I => \ALU.madd_cry_4\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27238\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__27238\,
            I => \N__27235\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__27235\,
            I => \N__27232\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__27232\,
            I => \ALU.madd_axb_6_l_ofx\
        );

    \I__4357\ : InMux
    port map (
            O => \N__27229\,
            I => \ALU.madd_cry_5\
        );

    \I__4356\ : InMux
    port map (
            O => \N__27226\,
            I => \ALU.madd_cry_6\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__27223\,
            I => \N__27220\
        );

    \I__4354\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27216\
        );

    \I__4353\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27213\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__27216\,
            I => \N__27210\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27207\
        );

    \I__4350\ : Span4Mux_v
    port map (
            O => \N__27210\,
            I => \N__27204\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__27207\,
            I => \N__27201\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__27204\,
            I => \ALU.madd_165\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__27201\,
            I => \ALU.madd_165\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__4345\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__4343\ : Span4Mux_v
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__27184\,
            I => \ALU.madd_axb_8_l_fx\
        );

    \I__4341\ : InMux
    port map (
            O => \N__27181\,
            I => \bfn_7_7_0_\
        );

    \I__4340\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27175\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27175\,
            I => \N__27172\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__4337\ : Odrv4
    port map (
            O => \N__27169\,
            I => \ALU.madd_axb_9_l_ofx\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__27166\,
            I => \ALU.a5_b_1_cascade_\
        );

    \I__4335\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27160\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27157\
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__27157\,
            I => \ALU.madd_50\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27150\
        );

    \I__4331\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27147\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__27150\,
            I => \ALU.madd_55\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__27147\,
            I => \ALU.madd_55\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__27142\,
            I => \ALU.madd_50_cascade_\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27135\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27132\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__27135\,
            I => \ALU.madd_73\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__27132\,
            I => \ALU.madd_73\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__27127\,
            I => \N__27124\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27118\
        );

    \I__4321\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27118\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__27118\,
            I => \ALU.madd_83\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27112\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__27112\,
            I => \N__27109\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__27109\,
            I => \N__27106\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__27106\,
            I => \N__27103\
        );

    \I__4315\ : Sp12to4
    port map (
            O => \N__27103\,
            I => \N__27100\
        );

    \I__4314\ : Odrv12
    port map (
            O => \N__27100\,
            I => \TXbuffer_RNO_1Z0Z_2\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27094\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__27094\,
            I => \N__27091\
        );

    \I__4311\ : Span4Mux_v
    port map (
            O => \N__27091\,
            I => \N__27088\
        );

    \I__4310\ : Span4Mux_h
    port map (
            O => \N__27088\,
            I => \N__27085\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__27085\,
            I => \TXbuffer_18_15_ns_1_2\
        );

    \I__4308\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27079\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__27079\,
            I => \N__27076\
        );

    \I__4306\ : Sp12to4
    port map (
            O => \N__27076\,
            I => \N__27071\
        );

    \I__4305\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27068\
        );

    \I__4304\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27065\
        );

    \I__4303\ : Span12Mux_v
    port map (
            O => \N__27071\,
            I => \N__27062\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__27068\,
            I => \clkdivZ0Z_1\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__27065\,
            I => \clkdivZ0Z_1\
        );

    \I__4300\ : Odrv12
    port map (
            O => \N__27062\,
            I => \clkdivZ0Z_1\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27052\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__27052\,
            I => \N__27047\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27044\
        );

    \I__4296\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27041\
        );

    \I__4295\ : Span12Mux_v
    port map (
            O => \N__27047\,
            I => \N__27038\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__27044\,
            I => \clkdivZ0Z_2\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__27041\,
            I => \clkdivZ0Z_2\
        );

    \I__4292\ : Odrv12
    port map (
            O => \N__27038\,
            I => \clkdivZ0Z_2\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__27031\,
            I => \N__27028\
        );

    \I__4290\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27025\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__27025\,
            I => \N__27022\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__27022\,
            I => \N__27019\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__27019\,
            I => \N__27016\
        );

    \I__4286\ : IoSpan4Mux
    port map (
            O => \N__27016\,
            I => \N__27012\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__27015\,
            I => \N__27009\
        );

    \I__4284\ : IoSpan4Mux
    port map (
            O => \N__27012\,
            I => \N__27005\
        );

    \I__4283\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27002\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26999\
        );

    \I__4281\ : Span4Mux_s1_h
    port map (
            O => \N__27005\,
            I => \N__26996\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27002\,
            I => \clkdivZ0Z_3\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__26999\,
            I => \clkdivZ0Z_3\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__26996\,
            I => \clkdivZ0Z_3\
        );

    \I__4277\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26986\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26986\,
            I => \N__26983\
        );

    \I__4275\ : Span4Mux_h
    port map (
            O => \N__26983\,
            I => \N__26980\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__26977\,
            I => \N__26972\
        );

    \I__4272\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26969\
        );

    \I__4271\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26966\
        );

    \I__4270\ : Span4Mux_v
    port map (
            O => \N__26972\,
            I => \N__26963\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__26969\,
            I => \clkdivZ0Z_0\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__26966\,
            I => \clkdivZ0Z_0\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__26963\,
            I => \clkdivZ0Z_0\
        );

    \I__4266\ : IoInMux
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__4264\ : Span12Mux_s11_h
    port map (
            O => \N__26950\,
            I => \N__26947\
        );

    \I__4263\ : Span12Mux_v
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__4262\ : Odrv12
    port map (
            O => \N__26944\,
            I => params5
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \ALU.madd_axb_3_cascade_\
        );

    \I__4260\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26932\
        );

    \I__4259\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26932\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26932\,
            I => \N__26929\
        );

    \I__4257\ : Odrv12
    port map (
            O => \N__26929\,
            I => \ALU.madd_14\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26923\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__26923\,
            I => \N__26920\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__26920\,
            I => \ALU.madd_cry_0_ma\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__26917\,
            I => \N__26914\
        );

    \I__4252\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__26908\,
            I => \ALU.madd_axb_0_l_ofx\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__26905\,
            I => \ALU.madd_73_0_cascade_\
        );

    \I__4248\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26899\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__26899\,
            I => \N__26896\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__26896\,
            I => \ALU.a1_b_5\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__26893\,
            I => \N__26890\
        );

    \I__4244\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26886\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26883\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__26886\,
            I => \ALU.a2_b_4\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26883\,
            I => \ALU.a2_b_4\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__26878\,
            I => \ALU.a1_b_5_cascade_\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26871\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26868\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__26871\,
            I => \N__26865\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__26868\,
            I => \b_fastZ0Z_1\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__26865\,
            I => \b_fastZ0Z_1\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__26860\,
            I => \N__26853\
        );

    \I__4233\ : CascadeMux
    port map (
            O => \N__26859\,
            I => \N__26847\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__26858\,
            I => \N__26841\
        );

    \I__4231\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26834\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26834\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26834\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26829\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26824\
        );

    \I__4226\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26821\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26816\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26816\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26809\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26809\
        );

    \I__4221\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26809\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__26834\,
            I => \N__26806\
        );

    \I__4219\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26803\
        );

    \I__4218\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26800\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26794\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26791\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26788\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__26824\,
            I => \N__26783\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__26821\,
            I => \N__26783\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26816\,
            I => \N__26780\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__26809\,
            I => \N__26775\
        );

    \I__4210\ : Span4Mux_v
    port map (
            O => \N__26806\,
            I => \N__26775\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__26803\,
            I => \N__26772\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__26800\,
            I => \N__26769\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26762\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26762\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26762\
        );

    \I__4204\ : Sp12to4
    port map (
            O => \N__26794\,
            I => \N__26757\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26791\,
            I => \N__26757\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__26788\,
            I => \N__26752\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__26783\,
            I => \N__26752\
        );

    \I__4200\ : Span4Mux_h
    port map (
            O => \N__26780\,
            I => \N__26747\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__26775\,
            I => \N__26747\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__26772\,
            I => \b_2_repZ0Z2\
        );

    \I__4197\ : Odrv12
    port map (
            O => \N__26769\,
            I => \b_2_repZ0Z2\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26762\,
            I => \b_2_repZ0Z2\
        );

    \I__4195\ : Odrv12
    port map (
            O => \N__26757\,
            I => \b_2_repZ0Z2\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__26752\,
            I => \b_2_repZ0Z2\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__26747\,
            I => \b_2_repZ0Z2\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__26734\,
            I => \ALU.r4_RNIMTDQZ0Z_1_cascade_\
        );

    \I__4191\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26728\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26728\,
            I => \ALU.b_7_ns_1_1\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26719\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26719\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26715\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26712\
        );

    \I__4185\ : Odrv4
    port map (
            O => \N__26715\,
            I => \ALU.madd_46\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__26712\,
            I => \ALU.madd_46\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__26707\,
            I => \N__26704\
        );

    \I__4182\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26701\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__26701\,
            I => \N__26698\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__26698\,
            I => \ALU.a5_b_1\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__26695\,
            I => \ALU.madd_18_cascade_\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__26692\,
            I => \ALU.madd_43_cascade_\
        );

    \I__4177\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26683\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26688\,
            I => \N__26683\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26683\,
            I => \ALU.a2_b_3\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26676\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26673\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26676\,
            I => \ALU.madd_332\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__26673\,
            I => \ALU.madd_332\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__26665\,
            I => \ALU.madd_94\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26658\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26655\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__26658\,
            I => \ALU.madd_33\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26655\,
            I => \ALU.madd_33\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26647\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26647\,
            I => \ALU.madd_38\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26640\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26637\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__26640\,
            I => \ALU.a0_b_6\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26637\,
            I => \ALU.a0_b_6\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__26632\,
            I => \N__26629\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26629\,
            I => \N__26625\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26622\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26625\,
            I => \N__26619\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__26622\,
            I => \ALU.madd_51\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__26619\,
            I => \ALU.madd_51\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__26614\,
            I => \ALU.madd_51_cascade_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26607\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26604\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26607\,
            I => \ALU.madd_43\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26604\,
            I => \ALU.madd_43\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26593\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26593\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26593\,
            I => \ALU.madd_331\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26584\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26584\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__26584\,
            I => \ALU.a1_b_4\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26578\,
            I => \ALU.madd_87\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26572\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26572\,
            I => \N__26569\
        );

    \I__4137\ : Span4Mux_s1_v
    port map (
            O => \N__26569\,
            I => \N__26565\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26562\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__26565\,
            I => \ALU.madd_110\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26562\,
            I => \ALU.madd_110\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26553\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26550\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__26553\,
            I => \ALU.madd_115\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26550\,
            I => \ALU.madd_115\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26539\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26539\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26539\,
            I => \ALU.madd_124\
        );

    \I__4126\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \ALU.madd_124_cascade_\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26528\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26523\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26523\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26528\,
            I => \N__26518\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26523\,
            I => \N__26518\
        );

    \I__4120\ : Odrv12
    port map (
            O => \N__26518\,
            I => \ALU.madd_160\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__26515\,
            I => \N__26509\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26505\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26513\,
            I => \N__26501\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26498\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26495\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26492\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26489\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26486\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26483\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__26498\,
            I => \N__26480\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__26495\,
            I => \N__26477\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26492\,
            I => \N__26474\
        );

    \I__4107\ : Span12Mux_s7_v
    port map (
            O => \N__26489\,
            I => \N__26471\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26466\
        );

    \I__4105\ : Span4Mux_v
    port map (
            O => \N__26483\,
            I => \N__26466\
        );

    \I__4104\ : Span12Mux_s7_v
    port map (
            O => \N__26480\,
            I => \N__26463\
        );

    \I__4103\ : Span12Mux_s4_h
    port map (
            O => \N__26477\,
            I => \N__26458\
        );

    \I__4102\ : Span12Mux_s1_v
    port map (
            O => \N__26474\,
            I => \N__26458\
        );

    \I__4101\ : Odrv12
    port map (
            O => \N__26471\,
            I => \ALU.r6_RNIE0JB2Z0Z_6\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__26466\,
            I => \ALU.r6_RNIE0JB2Z0Z_6\
        );

    \I__4099\ : Odrv12
    port map (
            O => \N__26463\,
            I => \ALU.r6_RNIE0JB2Z0Z_6\
        );

    \I__4098\ : Odrv12
    port map (
            O => \N__26458\,
            I => \ALU.r6_RNIE0JB2Z0Z_6\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26444\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26448\,
            I => \N__26441\
        );

    \I__4095\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26438\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26444\,
            I => \N__26432\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26441\,
            I => \N__26429\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26426\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26423\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26420\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26417\
        );

    \I__4088\ : Span4Mux_v
    port map (
            O => \N__26432\,
            I => \N__26414\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__26429\,
            I => \N__26411\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__26426\,
            I => \N__26406\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__26423\,
            I => \N__26406\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__26420\,
            I => \N__26403\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26417\,
            I => \N__26400\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__26414\,
            I => \N__26395\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__26411\,
            I => \N__26395\
        );

    \I__4080\ : Span4Mux_v
    port map (
            O => \N__26406\,
            I => \N__26390\
        );

    \I__4079\ : Span4Mux_v
    port map (
            O => \N__26403\,
            I => \N__26390\
        );

    \I__4078\ : Odrv12
    port map (
            O => \N__26400\,
            I => \ALU.r4_RNI68Q22Z0Z_6\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__26395\,
            I => \ALU.r4_RNI68Q22Z0Z_6\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__26390\,
            I => \ALU.r4_RNI68Q22Z0Z_6\
        );

    \I__4075\ : CascadeMux
    port map (
            O => \N__26383\,
            I => \N__26380\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26377\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26377\,
            I => \ALU.a3_b_1\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__26374\,
            I => \ALU.a3_b_1_cascade_\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__26371\,
            I => \N__26368\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26365\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__26365\,
            I => \N__26362\
        );

    \I__4068\ : Odrv12
    port map (
            O => \N__26362\,
            I => \ALU.r5_RNIK81F5Z0Z_13\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26356\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26356\,
            I => \N__26353\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__26353\,
            I => \ALU.r0_12_prm_5_13_s0_c_RNOZ0\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__26350\,
            I => \N__26347\
        );

    \I__4063\ : InMux
    port map (
            O => \N__26347\,
            I => \N__26344\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26344\,
            I => \N__26341\
        );

    \I__4061\ : Span4Mux_v
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26338\,
            I => \ALU.r0_12_prm_6_13_s0_c_RNOZ0\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__26335\,
            I => \N__26332\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26329\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__26326\,
            I => \ALU.r0_12_prm_7_13_s0_c_RNOZ0\
        );

    \I__4055\ : CascadeMux
    port map (
            O => \N__26323\,
            I => \N__26320\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26316\
        );

    \I__4053\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26313\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__26316\,
            I => \N__26310\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__26313\,
            I => \ALU.madd_334\
        );

    \I__4050\ : Odrv12
    port map (
            O => \N__26310\,
            I => \ALU.madd_334\
        );

    \I__4049\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26301\
        );

    \I__4048\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26298\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__26301\,
            I => \N__26295\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__26298\,
            I => \ALU.madd_333\
        );

    \I__4045\ : Odrv12
    port map (
            O => \N__26295\,
            I => \ALU.madd_333\
        );

    \I__4044\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26287\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__26287\,
            I => \ALU.r0_12_prm_3_13_s0_sf\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26284\,
            I => \ALU.r0_12_s0_13\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26274\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26271\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26268\
        );

    \I__4038\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26265\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26262\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26274\,
            I => \N__26258\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__26271\,
            I => \N__26255\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__26268\,
            I => \N__26252\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__26265\,
            I => \N__26249\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26246\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26243\
        );

    \I__4030\ : Span4Mux_h
    port map (
            O => \N__26258\,
            I => \N__26232\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26232\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__26252\,
            I => \N__26232\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__26249\,
            I => \N__26232\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__26246\,
            I => \N__26227\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__26243\,
            I => \N__26227\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26224\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26221\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__26232\,
            I => \ALU.r0_12_13\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__26227\,
            I => \ALU.r0_12_13\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__26224\,
            I => \ALU.r0_12_13\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__26221\,
            I => \ALU.r0_12_13\
        );

    \I__4018\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26208\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26205\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26202\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__26205\,
            I => \N__26199\
        );

    \I__4014\ : Span4Mux_h
    port map (
            O => \N__26202\,
            I => \N__26193\
        );

    \I__4013\ : Span4Mux_h
    port map (
            O => \N__26199\,
            I => \N__26193\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26190\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__26193\,
            I => r0_13
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__26190\,
            I => r0_13
        );

    \I__4009\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26180\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26177\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26173\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26169\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__26177\,
            I => \N__26166\
        );

    \I__4004\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26163\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26173\,
            I => \N__26160\
        );

    \I__4002\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26157\
        );

    \I__4001\ : Span4Mux_v
    port map (
            O => \N__26169\,
            I => \N__26149\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__26166\,
            I => \N__26149\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26146\
        );

    \I__3998\ : Span4Mux_h
    port map (
            O => \N__26160\,
            I => \N__26141\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26141\
        );

    \I__3996\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26138\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26135\
        );

    \I__3994\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26132\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__26149\,
            I => \ALU.r0_12_11\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__26146\,
            I => \ALU.r0_12_11\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__26141\,
            I => \ALU.r0_12_11\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__26138\,
            I => \ALU.r0_12_11\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__26135\,
            I => \ALU.r0_12_11\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__26132\,
            I => \ALU.r0_12_11\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26115\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26112\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26108\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__26105\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26102\
        );

    \I__3982\ : Span4Mux_v
    port map (
            O => \N__26108\,
            I => \N__26099\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__26105\,
            I => \N__26094\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26094\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__26099\,
            I => \N__26091\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__26094\,
            I => \N__26088\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__26091\,
            I => r5_11
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__26088\,
            I => r5_11
        );

    \I__3975\ : InMux
    port map (
            O => \N__26083\,
            I => \N__26080\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__26080\,
            I => \N__26075\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26072\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26069\
        );

    \I__3971\ : Span4Mux_s1_h
    port map (
            O => \N__26075\,
            I => \N__26064\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__26072\,
            I => \N__26064\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__26069\,
            I => \N__26061\
        );

    \I__3968\ : Span4Mux_h
    port map (
            O => \N__26064\,
            I => \N__26058\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__26061\,
            I => \N__26055\
        );

    \I__3966\ : Odrv4
    port map (
            O => \N__26058\,
            I => r5_12
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__26055\,
            I => r5_12
        );

    \I__3964\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26046\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26042\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__26046\,
            I => \N__26039\
        );

    \I__3961\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26036\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26042\,
            I => \N__26029\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__26039\,
            I => \N__26029\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__26036\,
            I => \N__26029\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__26029\,
            I => r5_13
        );

    \I__3956\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26022\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26018\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__26015\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26012\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26018\,
            I => \N__26009\
        );

    \I__3951\ : Span4Mux_s3_h
    port map (
            O => \N__26015\,
            I => \N__26006\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26003\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__26009\,
            I => \N__25998\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__26006\,
            I => \N__25998\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__26003\,
            I => r5_14
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__25998\,
            I => r5_14
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__3944\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25983\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25980\
        );

    \I__3942\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25977\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25973\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__25986\,
            I => \N__25969\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25965\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__25980\,
            I => \N__25962\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__25977\,
            I => \N__25959\
        );

    \I__3936\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25956\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__25973\,
            I => \N__25953\
        );

    \I__3934\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25950\
        );

    \I__3933\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25947\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25944\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__25965\,
            I => \ALU.r0_12_15\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__25962\,
            I => \ALU.r0_12_15\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__25959\,
            I => \ALU.r0_12_15\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__25956\,
            I => \ALU.r0_12_15\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__25953\,
            I => \ALU.r0_12_15\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__25950\,
            I => \ALU.r0_12_15\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__25947\,
            I => \ALU.r0_12_15\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__25944\,
            I => \ALU.r0_12_15\
        );

    \I__3923\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25923\
        );

    \I__3922\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25919\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__25923\,
            I => \N__25916\
        );

    \I__3920\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25913\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25910\
        );

    \I__3918\ : Span4Mux_h
    port map (
            O => \N__25916\,
            I => \N__25907\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25904\
        );

    \I__3916\ : Span12Mux_s5_h
    port map (
            O => \N__25910\,
            I => \N__25901\
        );

    \I__3915\ : Span4Mux_v
    port map (
            O => \N__25907\,
            I => \N__25898\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__25904\,
            I => r5_5
        );

    \I__3913\ : Odrv12
    port map (
            O => \N__25901\,
            I => r5_5
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__25898\,
            I => r5_5
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__25891\,
            I => \ALU.a_3_ns_1_14_cascade_\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25884\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25887\,
            I => \N__25881\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__25884\,
            I => \N__25877\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__25881\,
            I => \N__25874\
        );

    \I__3906\ : InMux
    port map (
            O => \N__25880\,
            I => \N__25871\
        );

    \I__3905\ : Span4Mux_v
    port map (
            O => \N__25877\,
            I => \N__25866\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__25874\,
            I => \N__25866\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__25871\,
            I => r4_14
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__25866\,
            I => r4_14
        );

    \I__3901\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25858\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25854\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25851\
        );

    \I__3898\ : Span4Mux_v
    port map (
            O => \N__25854\,
            I => \N__25848\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__25851\,
            I => \N__25845\
        );

    \I__3896\ : Span4Mux_h
    port map (
            O => \N__25848\,
            I => \N__25839\
        );

    \I__3895\ : Span4Mux_h
    port map (
            O => \N__25845\,
            I => \N__25839\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25836\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__25839\,
            I => r2_14
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__25836\,
            I => r2_14
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__25831\,
            I => \N__25827\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25824\
        );

    \I__3889\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25821\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__25824\,
            I => \N__25817\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25814\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25811\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__25817\,
            I => \N__25808\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__25814\,
            I => \N__25805\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__25811\,
            I => r3_14
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__25808\,
            I => r3_14
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__25805\,
            I => r3_14
        );

    \I__3880\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25793\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25790\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25787\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25793\,
            I => \N__25784\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25790\,
            I => \N__25781\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25776\
        );

    \I__3874\ : Span4Mux_s3_h
    port map (
            O => \N__25784\,
            I => \N__25776\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__25781\,
            I => \N__25773\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__25776\,
            I => r7_14
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__25773\,
            I => r7_14
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__25768\,
            I => \ALU.a_6_ns_1_14_cascade_\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25765\,
            I => \N__25760\
        );

    \I__3868\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25757\
        );

    \I__3867\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25754\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__25760\,
            I => \N__25751\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25757\,
            I => \N__25748\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__25754\,
            I => \N__25745\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__25751\,
            I => \N__25742\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__25748\,
            I => r6_14
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__25745\,
            I => r6_14
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25742\,
            I => r6_14
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__25735\,
            I => \ALU.r6_RNID4772Z0Z_14_cascade_\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__25729\,
            I => \N__25726\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__25726\,
            I => \ALU.r5_RNI54M52Z0Z_14\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25716\
        );

    \I__3853\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25713\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__25716\,
            I => \N__25710\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__25713\,
            I => \N__25707\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__25710\,
            I => \N__25701\
        );

    \I__3849\ : Span4Mux_v
    port map (
            O => \N__25707\,
            I => \N__25701\
        );

    \I__3848\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25698\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__25701\,
            I => r0_14
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__25698\,
            I => r0_14
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__25693\,
            I => \N__25688\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__25692\,
            I => \N__25685\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25665\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25665\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25665\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25665\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25665\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25665\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25657\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25657\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25652\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25652\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25644\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25637\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25637\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25637\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25634\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25652\,
            I => \N__25631\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25620\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25620\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25620\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25648\,
            I => \N__25620\
        );

    \I__3823\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25620\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__25644\,
            I => \N__25615\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__25637\,
            I => \N__25615\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__25634\,
            I => \N__25610\
        );

    \I__3819\ : Span4Mux_h
    port map (
            O => \N__25631\,
            I => \N__25610\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25620\,
            I => \aZ0Z_0\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__25615\,
            I => \aZ0Z_0\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__25610\,
            I => \aZ0Z_0\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25591\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25591\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25586\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25600\,
            I => \N__25586\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25581\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25581\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25572\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__25596\,
            I => \N__25566\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__25591\,
            I => \N__25560\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25586\,
            I => \N__25557\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25581\,
            I => \N__25554\
        );

    \I__3804\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25541\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25541\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25541\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25541\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25576\,
            I => \N__25541\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25541\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25572\,
            I => \N__25538\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25531\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25531\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25531\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25522\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25522\
        );

    \I__3792\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25522\
        );

    \I__3791\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25522\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__25560\,
            I => \N__25519\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__25557\,
            I => \N__25512\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__25554\,
            I => \N__25512\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25512\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__25538\,
            I => \N__25509\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__25531\,
            I => \N__25506\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25522\,
            I => \aZ0Z_2\
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__25519\,
            I => \aZ0Z_2\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__25512\,
            I => \aZ0Z_2\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__25509\,
            I => \aZ0Z_2\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__25506\,
            I => \aZ0Z_2\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__25495\,
            I => \ALU.a_3_ns_1_15_cascade_\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25489\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25489\,
            I => \N__25486\
        );

    \I__3776\ : Odrv12
    port map (
            O => \N__25486\,
            I => \ALU.r5_RNI98M52Z0Z_15\
        );

    \I__3775\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25480\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25475\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25472\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25469\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__25475\,
            I => \N__25464\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__25472\,
            I => \N__25464\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25469\,
            I => \N__25461\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__25464\,
            I => \N__25458\
        );

    \I__3767\ : Odrv12
    port map (
            O => \N__25461\,
            I => r4_10
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__25458\,
            I => r4_10
        );

    \I__3765\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25449\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25445\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25442\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25439\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25445\,
            I => \N__25436\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__25442\,
            I => \N__25431\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25431\
        );

    \I__3758\ : Odrv12
    port map (
            O => \N__25436\,
            I => r4_12
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__25431\,
            I => r4_12
        );

    \I__3756\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25423\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__25420\,
            I => \N__25416\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25413\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__25416\,
            I => \N__25407\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25413\,
            I => \N__25407\
        );

    \I__3750\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25404\
        );

    \I__3749\ : Span4Mux_h
    port map (
            O => \N__25407\,
            I => \N__25401\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__25404\,
            I => \N__25398\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__25401\,
            I => r4_13
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__25398\,
            I => r4_13
        );

    \I__3745\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25388\
        );

    \I__3744\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25385\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25382\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25388\,
            I => \N__25379\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__25385\,
            I => \N__25376\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__25382\,
            I => \N__25373\
        );

    \I__3739\ : Span4Mux_h
    port map (
            O => \N__25379\,
            I => \N__25370\
        );

    \I__3738\ : Span12Mux_v
    port map (
            O => \N__25376\,
            I => \N__25365\
        );

    \I__3737\ : Span12Mux_s11_v
    port map (
            O => \N__25373\,
            I => \N__25365\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__25370\,
            I => r4_5
        );

    \I__3735\ : Odrv12
    port map (
            O => \N__25365\,
            I => r4_5
        );

    \I__3734\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25357\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__25357\,
            I => \N__25353\
        );

    \I__3732\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25349\
        );

    \I__3731\ : Span4Mux_h
    port map (
            O => \N__25353\,
            I => \N__25346\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25343\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25349\,
            I => \N__25340\
        );

    \I__3728\ : Span4Mux_v
    port map (
            O => \N__25346\,
            I => \N__25337\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25343\,
            I => \N__25334\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__25340\,
            I => \N__25329\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__25337\,
            I => \N__25329\
        );

    \I__3724\ : Sp12to4
    port map (
            O => \N__25334\,
            I => \N__25326\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__25329\,
            I => r4_6
        );

    \I__3722\ : Odrv12
    port map (
            O => \N__25326\,
            I => r4_6
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__25321\,
            I => \ALU.r6_RNI7L2O1Z0Z_4_cascade_\
        );

    \I__3720\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25314\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25311\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25308\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__25311\,
            I => \N__25305\
        );

    \I__3716\ : Span4Mux_h
    port map (
            O => \N__25308\,
            I => \N__25301\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__25305\,
            I => \N__25298\
        );

    \I__3714\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25295\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__25301\,
            I => r2_12
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__25298\,
            I => r2_12
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__25295\,
            I => r2_12
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__25288\,
            I => \N__25284\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__25287\,
            I => \N__25281\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25276\
        );

    \I__3707\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25276\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25276\,
            I => \N__25272\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25269\
        );

    \I__3704\ : Odrv12
    port map (
            O => \N__25272\,
            I => r2_4
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__25269\,
            I => r2_4
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__25264\,
            I => \TXbuffer_18_6_ns_1_4_cascade_\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25258\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25254\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25250\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__25254\,
            I => \N__25247\
        );

    \I__3697\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25244\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__25250\,
            I => \N__25241\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__25247\,
            I => \N__25236\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25236\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__25241\,
            I => r6_12
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__25236\,
            I => r6_12
        );

    \I__3691\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25228\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__25228\,
            I => \N__25225\
        );

    \I__3689\ : Span4Mux_v
    port map (
            O => \N__25225\,
            I => \N__25222\
        );

    \I__3688\ : Sp12to4
    port map (
            O => \N__25222\,
            I => \N__25219\
        );

    \I__3687\ : Odrv12
    port map (
            O => \N__25219\,
            I => \TXbuffer_RNO_6Z0Z_4\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__3685\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25209\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__25212\,
            I => \N__25206\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__25209\,
            I => \N__25203\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25200\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__25203\,
            I => \N__25197\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25200\,
            I => \N__25193\
        );

    \I__3679\ : Span4Mux_s2_h
    port map (
            O => \N__25197\,
            I => \N__25190\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__25196\,
            I => \N__25187\
        );

    \I__3677\ : Span12Mux_v
    port map (
            O => \N__25193\,
            I => \N__25184\
        );

    \I__3676\ : Span4Mux_h
    port map (
            O => \N__25190\,
            I => \N__25181\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25187\,
            I => \N__25178\
        );

    \I__3674\ : Odrv12
    port map (
            O => \N__25184\,
            I => r1_11
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__25181\,
            I => r1_11
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__25178\,
            I => r1_11
        );

    \I__3671\ : InMux
    port map (
            O => \N__25171\,
            I => \N__25167\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25164\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25167\,
            I => \N__25160\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__25164\,
            I => \N__25157\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__25163\,
            I => \N__25154\
        );

    \I__3666\ : Span12Mux_s5_h
    port map (
            O => \N__25160\,
            I => \N__25151\
        );

    \I__3665\ : Span4Mux_v
    port map (
            O => \N__25157\,
            I => \N__25148\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25145\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__25151\,
            I => r1_12
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__25148\,
            I => r1_12
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__25145\,
            I => r1_12
        );

    \I__3660\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25133\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__25137\,
            I => \N__25130\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25127\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25124\
        );

    \I__3656\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25121\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__25127\,
            I => \N__25118\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__25124\,
            I => \N__25113\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25121\,
            I => \N__25113\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__25118\,
            I => \N__25110\
        );

    \I__3651\ : Span4Mux_v
    port map (
            O => \N__25113\,
            I => \N__25107\
        );

    \I__3650\ : Odrv4
    port map (
            O => \N__25110\,
            I => r1_13
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__25107\,
            I => r1_13
        );

    \I__3648\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25093\
        );

    \I__3647\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25080\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25080\
        );

    \I__3645\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25080\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25080\
        );

    \I__3643\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25080\
        );

    \I__3642\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25080\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__25093\,
            I => \N__25068\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25080\,
            I => \N__25068\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25061\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25061\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25052\
        );

    \I__3636\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25052\
        );

    \I__3635\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25052\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25052\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__25073\,
            I => \N__25048\
        );

    \I__3632\ : Span12Mux_v
    port map (
            O => \N__25068\,
            I => \N__25043\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25040\
        );

    \I__3630\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25037\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__25061\,
            I => \N__25032\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25032\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25023\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25023\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25023\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25023\
        );

    \I__3623\ : Odrv12
    port map (
            O => \N__25043\,
            I => \bZ0Z_0\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__25040\,
            I => \bZ0Z_0\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__25037\,
            I => \bZ0Z_0\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__25032\,
            I => \bZ0Z_0\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25023\,
            I => \bZ0Z_0\
        );

    \I__3618\ : InMux
    port map (
            O => \N__25012\,
            I => \N__25008\
        );

    \I__3617\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25005\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__25008\,
            I => \N__24995\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24992\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24989\
        );

    \I__3613\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24984\
        );

    \I__3612\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24984\
        );

    \I__3611\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24975\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24975\
        );

    \I__3609\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24975\
        );

    \I__3608\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24975\
        );

    \I__3607\ : Span4Mux_v
    port map (
            O => \N__24995\,
            I => \N__24972\
        );

    \I__3606\ : Odrv12
    port map (
            O => \N__24992\,
            I => \a_0_repZ0Z1\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__24989\,
            I => \a_0_repZ0Z1\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__24984\,
            I => \a_0_repZ0Z1\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24975\,
            I => \a_0_repZ0Z1\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__24972\,
            I => \a_0_repZ0Z1\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__24961\,
            I => \ALU.a_6_ns_1_4_cascade_\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__24958\,
            I => \N__24954\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__24957\,
            I => \N__24950\
        );

    \I__3598\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24947\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24942\
        );

    \I__3596\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24942\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24939\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__24942\,
            I => \N__24936\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__24939\,
            I => \N__24933\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__24936\,
            I => \N__24930\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__24933\,
            I => r3_4
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__24930\,
            I => r3_4
        );

    \I__3589\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24919\
        );

    \I__3588\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24916\
        );

    \I__3587\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24913\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__24922\,
            I => \N__24910\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24902\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__24916\,
            I => \N__24899\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__24913\,
            I => \N__24896\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24893\
        );

    \I__3581\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24882\
        );

    \I__3580\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24882\
        );

    \I__3579\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24882\
        );

    \I__3578\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24882\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24882\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__24902\,
            I => \N__24879\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__24899\,
            I => \N__24874\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__24896\,
            I => \N__24874\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__24893\,
            I => \b_0_repZ0Z1\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__24882\,
            I => \b_0_repZ0Z1\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__24879\,
            I => \b_0_repZ0Z1\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__24874\,
            I => \b_0_repZ0Z1\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__24865\,
            I => \ALU.b_6_ns_1_4_cascade_\
        );

    \I__3568\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24859\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__24859\,
            I => \N__24856\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__24856\,
            I => \N__24853\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__24853\,
            I => \ALU.r6_RNI7L2O1Z0Z_4\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__24850\,
            I => \TXbuffer_18_3_ns_1_3_cascade_\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__24847\,
            I => \TXbuffer_RNO_5Z0Z_3_cascade_\
        );

    \I__3562\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24841\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__24841\,
            I => \N__24838\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__3559\ : Span4Mux_v
    port map (
            O => \N__24835\,
            I => \N__24832\
        );

    \I__3558\ : Sp12to4
    port map (
            O => \N__24832\,
            I => \N__24829\
        );

    \I__3557\ : Span12Mux_s5_h
    port map (
            O => \N__24829\,
            I => \N__24826\
        );

    \I__3556\ : Odrv12
    port map (
            O => \N__24826\,
            I => \TXbuffer_18_15_ns_1_3\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24823\,
            I => \N__24820\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__24820\,
            I => \N__24817\
        );

    \I__3553\ : Span4Mux_h
    port map (
            O => \N__24817\,
            I => \N__24812\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24809\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24815\,
            I => \N__24806\
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__24812\,
            I => r2_11
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24809\,
            I => r2_11
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__24806\,
            I => r2_11
        );

    \I__3547\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24796\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__24796\,
            I => \N__24791\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24788\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24785\
        );

    \I__3543\ : Span4Mux_h
    port map (
            O => \N__24791\,
            I => \N__24780\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__24788\,
            I => \N__24780\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__24785\,
            I => \N__24777\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__24780\,
            I => r2_3
        );

    \I__3539\ : Odrv12
    port map (
            O => \N__24777\,
            I => r2_3
        );

    \I__3538\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24769\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24769\,
            I => \N__24764\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24761\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24758\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__24764\,
            I => \N__24751\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24751\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__24758\,
            I => \N__24751\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__24751\,
            I => \N__24748\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__24748\,
            I => r6_11
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__24745\,
            I => \TXbuffer_18_6_ns_1_3_cascade_\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24739\,
            I => \TXbuffer_RNO_6Z0Z_3\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24736\,
            I => \N__24731\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24735\,
            I => \N__24728\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24734\,
            I => \N__24725\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24722\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__24728\,
            I => \N__24717\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24725\,
            I => \N__24717\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__24722\,
            I => r4_11
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__24717\,
            I => r4_11
        );

    \I__3518\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24707\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24702\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24696\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24693\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24688\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24688\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__24702\,
            I => \N__24685\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24680\
        );

    \I__3510\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24680\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24677\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24696\,
            I => \N__24674\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__24693\,
            I => \N__24671\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24688\,
            I => \N__24664\
        );

    \I__3505\ : Span4Mux_h
    port map (
            O => \N__24685\,
            I => \N__24664\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24664\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__24677\,
            I => \b_1_repZ0Z1\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__24674\,
            I => \b_1_repZ0Z1\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__24671\,
            I => \b_1_repZ0Z1\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__24664\,
            I => \b_1_repZ0Z1\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__24655\,
            I => \N__24650\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24646\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__24653\,
            I => \N__24643\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24638\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24635\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24632\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24627\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24624\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24620\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24638\,
            I => \N__24617\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__24635\,
            I => \N__24614\
        );

    \I__3488\ : Span4Mux_v
    port map (
            O => \N__24632\,
            I => \N__24611\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24608\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24605\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24627\,
            I => \N__24602\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__24624\,
            I => \N__24599\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24596\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24620\,
            I => \N__24593\
        );

    \I__3481\ : Span4Mux_v
    port map (
            O => \N__24617\,
            I => \N__24582\
        );

    \I__3480\ : Span4Mux_v
    port map (
            O => \N__24614\,
            I => \N__24582\
        );

    \I__3479\ : Span4Mux_s2_h
    port map (
            O => \N__24611\,
            I => \N__24582\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24582\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24605\,
            I => \N__24582\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__24602\,
            I => \N__24578\
        );

    \I__3475\ : Sp12to4
    port map (
            O => \N__24599\,
            I => \N__24573\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24573\
        );

    \I__3473\ : Span4Mux_v
    port map (
            O => \N__24593\,
            I => \N__24568\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__24582\,
            I => \N__24568\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24565\
        );

    \I__3470\ : Sp12to4
    port map (
            O => \N__24578\,
            I => \N__24562\
        );

    \I__3469\ : Span12Mux_s6_v
    port map (
            O => \N__24573\,
            I => \N__24559\
        );

    \I__3468\ : Span4Mux_h
    port map (
            O => \N__24568\,
            I => \N__24556\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24565\,
            I => \b_1_repZ0Z2\
        );

    \I__3466\ : Odrv12
    port map (
            O => \N__24562\,
            I => \b_1_repZ0Z2\
        );

    \I__3465\ : Odrv12
    port map (
            O => \N__24559\,
            I => \b_1_repZ0Z2\
        );

    \I__3464\ : Odrv4
    port map (
            O => \N__24556\,
            I => \b_1_repZ0Z2\
        );

    \I__3463\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24544\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24544\,
            I => \N__24540\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24536\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__24540\,
            I => \N__24533\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24530\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24527\
        );

    \I__3457\ : Span4Mux_s2_h
    port map (
            O => \N__24533\,
            I => \N__24524\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24521\
        );

    \I__3455\ : Span4Mux_v
    port map (
            O => \N__24527\,
            I => \N__24518\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__24524\,
            I => r0_11
        );

    \I__3453\ : Odrv12
    port map (
            O => \N__24521\,
            I => r0_11
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__24518\,
            I => r0_11
        );

    \I__3451\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24508\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__24505\,
            I => \N__24502\
        );

    \I__3448\ : Span4Mux_h
    port map (
            O => \N__24502\,
            I => \N__24499\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__24499\,
            I => \ALU.madd_368\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__24496\,
            I => \N__24493\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24490\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__24490\,
            I => \ALU.a12_b_2\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \ALU.a12_b_2_cascade_\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__3439\ : Span4Mux_h
    port map (
            O => \N__24475\,
            I => \N__24472\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__24472\,
            I => \ALU.madd_372\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__24469\,
            I => \N__24466\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24463\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24459\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24456\
        );

    \I__3433\ : Span4Mux_s3_v
    port map (
            O => \N__24459\,
            I => \N__24453\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24450\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__24453\,
            I => \ALU.g1_2\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__24450\,
            I => \ALU.g1_2\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24442\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__3427\ : Span4Mux_s2_h
    port map (
            O => \N__24439\,
            I => \N__24436\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__24436\,
            I => \ALU.madd_311_0\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__24433\,
            I => \ALU.a_3_cascade_\
        );

    \I__3424\ : InMux
    port map (
            O => \N__24430\,
            I => \N__24427\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24424\
        );

    \I__3422\ : Span4Mux_h
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__24421\,
            I => \ALU.g1_1\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__24418\,
            I => \ALU.b_4_cascade_\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24412\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__3417\ : Odrv12
    port map (
            O => \N__24409\,
            I => \ALU.madd_214_0\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__24406\,
            I => \ALU.b_2_cascade_\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24400\,
            I => \N__24397\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__24397\,
            I => \ALU.madd_134_0_tz_0\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24388\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24388\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__3409\ : Span4Mux_s2_h
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__24382\,
            I => \N__24379\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__24379\,
            I => \ALU.madd_172_0\
        );

    \I__3406\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24373\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__24373\,
            I => \N__24370\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__24370\,
            I => \N__24367\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__24367\,
            I => \N__24364\
        );

    \I__3402\ : Span4Mux_v
    port map (
            O => \N__24364\,
            I => \N__24361\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__24361\,
            I => \ALU.r6_RNIA0841Z0Z_0\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__24355\,
            I => \ALU.madd_92\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24348\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24345\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24348\,
            I => \N__24342\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__24345\,
            I => \ALU.madd_120\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__24342\,
            I => \ALU.madd_120\
        );

    \I__3393\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24333\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24330\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24324\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24330\,
            I => \N__24324\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24321\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__24324\,
            I => \N__24318\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24315\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__24318\,
            I => \ALU.r6_RNII9FT1Z0Z_3\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__24315\,
            I => \ALU.r6_RNII9FT1Z0Z_3\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__24310\,
            I => \ALU.b_3_cascade_\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24304\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24304\,
            I => \N__24301\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__24301\,
            I => \N__24298\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__24298\,
            I => \N__24295\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__24295\,
            I => \ALU.un2_addsub_axb_3\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__24292\,
            I => \ALU.b_1_cascade_\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24286\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__24283\,
            I => \ALU.a4_b_1\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__24280\,
            I => \ALU.madd_38_cascade_\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__24277\,
            I => \ALU.madd_87_cascade_\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__24274\,
            I => \ALU.madd_92_cascade_\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__24268\,
            I => \ALU.madd_78_0\
        );

    \I__3369\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24259\
        );

    \I__3368\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24259\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24256\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__24256\,
            I => \ALU.madd_68\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__24253\,
            I => \ALU.madd_78_0_cascade_\
        );

    \I__3364\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24244\
        );

    \I__3363\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24244\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__24244\,
            I => \ALU.madd_60\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__24241\,
            I => \ALU.madd_332_cascade_\
        );

    \I__3360\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24234\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24231\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24234\,
            I => \ALU.madd_68_0\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__24231\,
            I => \ALU.madd_68_0\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24223\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24223\,
            I => \N__24220\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__24220\,
            I => \ALU.madd_46_0\
        );

    \I__3353\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24213\
        );

    \I__3352\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24210\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__24213\,
            I => \ALU.madd_100\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__24210\,
            I => \ALU.madd_100\
        );

    \I__3349\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24201\
        );

    \I__3348\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24198\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__24201\,
            I => \ALU.madd_105\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__24198\,
            I => \ALU.madd_105\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__24193\,
            I => \ALU.madd_46_0_cascade_\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24187\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__24187\,
            I => \ALU.madd_82_0\
        );

    \I__3342\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24178\
        );

    \I__3341\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24178\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__24178\,
            I => \ALU.a5_b_3\
        );

    \I__3339\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24172\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__24172\,
            I => \N__24169\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__24169\,
            I => \ALU.g2_0_0_0\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24162\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24159\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24156\
        );

    \I__3333\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24153\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__24156\,
            I => \ALU.a0_b_7\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24153\,
            I => \ALU.a0_b_7\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__24148\,
            I => \N__24145\
        );

    \I__3329\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24142\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24142\,
            I => \ALU.a5_b_0\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__24139\,
            I => \N__24135\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24132\
        );

    \I__3325\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24129\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__24132\,
            I => \N__24123\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__24129\,
            I => \N__24123\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__24128\,
            I => \N__24120\
        );

    \I__3321\ : Span4Mux_v
    port map (
            O => \N__24123\,
            I => \N__24117\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24114\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__24117\,
            I => \N__24111\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__24114\,
            I => r3_5
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__24111\,
            I => r3_5
        );

    \I__3316\ : InMux
    port map (
            O => \N__24106\,
            I => \N__24103\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__24103\,
            I => \N__24098\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__24102\,
            I => \N__24095\
        );

    \I__3313\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24092\
        );

    \I__3312\ : Span4Mux_h
    port map (
            O => \N__24098\,
            I => \N__24089\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24086\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__24092\,
            I => r3_13
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__24089\,
            I => r3_13
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24086\,
            I => r3_13
        );

    \I__3307\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24075\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24072\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__24068\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24072\,
            I => \N__24065\
        );

    \I__3303\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24062\
        );

    \I__3302\ : Span4Mux_v
    port map (
            O => \N__24068\,
            I => \N__24057\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__24065\,
            I => \N__24057\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24062\,
            I => \N__24054\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__24057\,
            I => r6_13
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__24054\,
            I => r6_13
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__24049\,
            I => \N__24046\
        );

    \I__3296\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24043\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__24043\,
            I => \N__24040\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__24040\,
            I => \TXbuffer_18_6_ns_1_5\
        );

    \I__3293\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24033\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24029\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__24033\,
            I => \N__24026\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24023\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24020\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__24026\,
            I => \N__24017\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__24023\,
            I => \N__24014\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__24020\,
            I => \N__24011\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__24017\,
            I => \N__24008\
        );

    \I__3284\ : Span4Mux_v
    port map (
            O => \N__24014\,
            I => \N__24005\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__24011\,
            I => r6_5
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__24008\,
            I => r6_5
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__24005\,
            I => r6_5
        );

    \I__3280\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__23995\,
            I => \TXbuffer_RNO_5Z0Z_5\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__23992\,
            I => \TXbuffer_RNO_6Z0Z_5_cascade_\
        );

    \I__3277\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23985\
        );

    \I__3276\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23982\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__23985\,
            I => \N__23978\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23982\,
            I => \N__23975\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23972\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__23978\,
            I => r7_13
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__23975\,
            I => r7_13
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__23972\,
            I => r7_13
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__23965\,
            I => \N__23961\
        );

    \I__3268\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23958\
        );

    \I__3267\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23954\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__23958\,
            I => \N__23951\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23948\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__23954\,
            I => \N__23945\
        );

    \I__3263\ : Span4Mux_h
    port map (
            O => \N__23951\,
            I => \N__23940\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23940\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__23945\,
            I => \N__23935\
        );

    \I__3260\ : Span4Mux_v
    port map (
            O => \N__23940\,
            I => \N__23935\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__23935\,
            I => r7_5
        );

    \I__3258\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23929\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__23929\,
            I => \TXbuffer_18_13_ns_1_5\
        );

    \I__3256\ : InMux
    port map (
            O => \N__23926\,
            I => \N__23923\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__23923\,
            I => \TXbuffer_18_10_ns_1_5\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__23920\,
            I => \ALU.a_3_ns_1_13_cascade_\
        );

    \I__3253\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23913\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23910\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23907\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23903\
        );

    \I__3249\ : Span4Mux_v
    port map (
            O => \N__23907\,
            I => \N__23900\
        );

    \I__3248\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23897\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__23903\,
            I => \N__23894\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__23900\,
            I => r2_13
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__23897\,
            I => r2_13
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__23894\,
            I => r2_13
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__23887\,
            I => \ALU.a_6_ns_1_13_cascade_\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__23884\,
            I => \ALU.r6_RNI90772Z0Z_13_cascade_\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23878\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23878\,
            I => \ALU.r5_RNI10M52Z0Z_13\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__23875\,
            I => \ALU.r5_RNIPV8A9Z0Z_13_cascade_\
        );

    \I__3238\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23867\
        );

    \I__3237\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23864\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__23870\,
            I => \N__23861\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__23867\,
            I => \N__23858\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23855\
        );

    \I__3233\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23852\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__23858\,
            I => \N__23849\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__23855\,
            I => \N__23846\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23843\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__23849\,
            I => r3_12
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__23846\,
            I => r3_12
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__23843\,
            I => r3_12
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__23836\,
            I => \N__23833\
        );

    \I__3225\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__3223\ : Span4Mux_v
    port map (
            O => \N__23827\,
            I => \N__23824\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__23824\,
            I => \ALU.r0_12_prm_7_15_s1_c_RNOZ0\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__23821\,
            I => \N__23818\
        );

    \I__3220\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23815\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23812\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__23812\,
            I => \N__23809\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__23809\,
            I => \ALU.r0_12_prm_6_15_s1_c_RNOZ0\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23800\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23797\
        );

    \I__3213\ : Span4Mux_h
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__23794\,
            I => \ALU.r0_12_prm_4_15_s1_c_RNOZ0\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23788\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23788\,
            I => \N__23785\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__23782\,
            I => \ALU.madd_axb_14\
        );

    \I__3207\ : InMux
    port map (
            O => \N__23779\,
            I => \ALU.r0_12_s1_15\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23771\
        );

    \I__3205\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23768\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23765\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23771\,
            I => \N__23762\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23757\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23765\,
            I => \N__23757\
        );

    \I__3200\ : Span4Mux_v
    port map (
            O => \N__23762\,
            I => \N__23752\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__23757\,
            I => \N__23752\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__23752\,
            I => r2_5
        );

    \I__3197\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23746\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23746\,
            I => \N__23742\
        );

    \I__3195\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23738\
        );

    \I__3194\ : Span4Mux_h
    port map (
            O => \N__23742\,
            I => \N__23735\
        );

    \I__3193\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23732\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23729\
        );

    \I__3191\ : Span4Mux_s3_v
    port map (
            O => \N__23735\,
            I => \N__23726\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__23732\,
            I => \N__23723\
        );

    \I__3189\ : Span4Mux_h
    port map (
            O => \N__23729\,
            I => \N__23720\
        );

    \I__3188\ : Span4Mux_v
    port map (
            O => \N__23726\,
            I => \N__23715\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__23723\,
            I => \N__23715\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__23720\,
            I => r2_6
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__23715\,
            I => r2_6
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__23710\,
            I => \N__23707\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23702\
        );

    \I__3182\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23699\
        );

    \I__3181\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23696\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__23702\,
            I => \N__23693\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__23699\,
            I => \N__23690\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23696\,
            I => \N__23687\
        );

    \I__3177\ : Span4Mux_v
    port map (
            O => \N__23693\,
            I => \N__23684\
        );

    \I__3176\ : Span4Mux_h
    port map (
            O => \N__23690\,
            I => \N__23679\
        );

    \I__3175\ : Span4Mux_h
    port map (
            O => \N__23687\,
            I => \N__23679\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__23684\,
            I => r2_9
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__23679\,
            I => r2_9
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__23674\,
            I => \ALU.a_3_ns_1_11_cascade_\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__23668\,
            I => \ALU.r5_RNI3VN52Z0Z_11\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__23665\,
            I => \N__23662\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23659\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23659\,
            I => \N__23654\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23651\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23648\
        );

    \I__3164\ : Span4Mux_v
    port map (
            O => \N__23654\,
            I => \N__23645\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23651\,
            I => \N__23642\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__23648\,
            I => \N__23639\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__23645\,
            I => \N__23636\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__23642\,
            I => r3_3
        );

    \I__3159\ : Odrv12
    port map (
            O => \N__23639\,
            I => r3_3
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__23636\,
            I => r3_3
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__23629\,
            I => \ALU.a_6_ns_1_3_cascade_\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__23626\,
            I => \ALU.a_3_ns_1_12_cascade_\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23618\
        );

    \I__3154\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23615\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23612\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23609\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23606\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23603\
        );

    \I__3149\ : Span4Mux_s3_h
    port map (
            O => \N__23609\,
            I => \N__23600\
        );

    \I__3148\ : Span4Mux_s3_h
    port map (
            O => \N__23606\,
            I => \N__23595\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__23603\,
            I => \N__23595\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__23600\,
            I => r7_12
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__23595\,
            I => r7_12
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__23590\,
            I => \ALU.a_6_ns_1_12_cascade_\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__23587\,
            I => \ALU.r6_RNI5S672Z0Z_12_cascade_\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23581\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__23581\,
            I => \ALU.r5_RNIS3672Z0Z_12\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23575\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23575\,
            I => \N__23572\
        );

    \I__3138\ : Span4Mux_h
    port map (
            O => \N__23572\,
            I => \N__23568\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__23571\,
            I => \N__23565\
        );

    \I__3136\ : Span4Mux_v
    port map (
            O => \N__23568\,
            I => \N__23561\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23558\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23555\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__23561\,
            I => r2_8
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23558\,
            I => r2_8
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23555\,
            I => r2_8
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__23548\,
            I => \N__23543\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23540\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23535\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23535\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23540\,
            I => \N__23532\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23535\,
            I => \N__23529\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__23532\,
            I => \N__23526\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__23529\,
            I => \N__23523\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__23526\,
            I => r3_8
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__23523\,
            I => r3_8
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__23518\,
            I => \ALU.b_6_ns_1_8_cascade_\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23515\,
            I => \N__23512\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23512\,
            I => \N__23509\
        );

    \I__3117\ : Odrv12
    port map (
            O => \N__23509\,
            I => \ALU.r6_RNIN53O1Z0Z_8\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__23506\,
            I => \ALU.a_6_ns_1_1_cascade_\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__23503\,
            I => \ALU.a_3_ns_1_10_cascade_\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__23500\,
            I => \ALU.r5_RNIVQN52Z0Z_10_cascade_\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23493\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23490\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23493\,
            I => \N__23487\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23484\
        );

    \I__3109\ : Sp12to4
    port map (
            O => \N__23487\,
            I => \N__23480\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__23484\,
            I => \N__23477\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23474\
        );

    \I__3106\ : Odrv12
    port map (
            O => \N__23480\,
            I => r0_6
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__23477\,
            I => r0_6
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__23474\,
            I => r0_6
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__23467\,
            I => \ALU.a_6_ns_1_5_cascade_\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__23464\,
            I => \N__23460\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23457\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23454\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23450\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23447\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__23453\,
            I => \N__23444\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__23450\,
            I => \N__23441\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__23447\,
            I => \N__23438\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23435\
        );

    \I__3093\ : Span4Mux_v
    port map (
            O => \N__23441\,
            I => \N__23432\
        );

    \I__3092\ : Span4Mux_v
    port map (
            O => \N__23438\,
            I => \N__23429\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23435\,
            I => r3_6
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__23432\,
            I => r3_6
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__23429\,
            I => r3_6
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__23422\,
            I => \ALU.a_6_ns_1_6_cascade_\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__23416\,
            I => \ALU.a_6_ns_1_9\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__23413\,
            I => \ALU.a_6_ns_1_8_cascade_\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23410\,
            I => \N__23407\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23407\,
            I => \N__23401\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23394\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23394\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23394\
        );

    \I__3079\ : Span4Mux_h
    port map (
            O => \N__23401\,
            I => \N__23389\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23389\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__23389\,
            I => \ALU.r6_RNIKG3D2Z0Z_8\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23380\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__23380\,
            I => \N__23375\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23370\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23370\
        );

    \I__3071\ : Span4Mux_h
    port map (
            O => \N__23375\,
            I => \N__23367\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__23370\,
            I => r2_2
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__23367\,
            I => r2_2
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__23362\,
            I => \N__23358\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__23361\,
            I => \N__23354\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23351\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23346\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23346\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__23351\,
            I => \N__23343\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23340\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__23343\,
            I => \N__23337\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__23340\,
            I => r3_2
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__23337\,
            I => r3_2
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__23332\,
            I => \ALU.b_6_ns_1_2_cascade_\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__23329\,
            I => \ALU.b_6_ns_1_3_cascade_\
        );

    \I__3056\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23322\
        );

    \I__3055\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23319\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23315\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__23319\,
            I => \N__23312\
        );

    \I__3052\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23309\
        );

    \I__3051\ : Span4Mux_s3_h
    port map (
            O => \N__23315\,
            I => \N__23306\
        );

    \I__3050\ : Span4Mux_v
    port map (
            O => \N__23312\,
            I => \N__23303\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__23309\,
            I => \N__23300\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__23306\,
            I => r7_0
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__23303\,
            I => r7_0
        );

    \I__3046\ : Odrv12
    port map (
            O => \N__23300\,
            I => r7_0
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__23293\,
            I => \ALU.b_6_ns_1_0_cascade_\
        );

    \I__3044\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23287\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23284\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__23284\,
            I => \N__23279\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23274\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23274\
        );

    \I__3039\ : Span4Mux_v
    port map (
            O => \N__23279\,
            I => \N__23271\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__23274\,
            I => r6_0
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__23271\,
            I => r6_0
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__23266\,
            I => \ALU.a_3_ns_1_6_cascade_\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23257\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23257\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23257\,
            I => \N__23253\
        );

    \I__3032\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23250\
        );

    \I__3031\ : Span4Mux_h
    port map (
            O => \N__23253\,
            I => \N__23247\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23244\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__23247\,
            I => \ALU.a8_b_4\
        );

    \I__3028\ : Odrv12
    port map (
            O => \N__23244\,
            I => \ALU.a8_b_4\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__23239\,
            I => \ALU.g0_7_x1_cascade_\
        );

    \I__3026\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__23233\,
            I => \ALU.madd_76_1\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__23230\,
            I => \N__23225\
        );

    \I__3023\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23221\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23218\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23215\
        );

    \I__3020\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23212\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__23221\,
            I => \N__23207\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__23218\,
            I => \N__23207\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__23215\,
            I => \N__23202\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23202\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__23207\,
            I => \ALU.r6_RNIPK3D2Z0Z_9\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__23202\,
            I => \ALU.r6_RNIPK3D2Z0Z_9\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__23197\,
            I => \N__23193\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__23196\,
            I => \N__23190\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23185\
        );

    \I__3010\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23185\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23182\
        );

    \I__3008\ : Span4Mux_s1_h
    port map (
            O => \N__23182\,
            I => \N__23179\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__23179\,
            I => \ALU.a9_b_4\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__23176\,
            I => \ALU.a_8_cascade_\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23170\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23167\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__23167\,
            I => \ALU.madd_224_0\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__23164\,
            I => \N__23160\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23163\,
            I => \N__23155\
        );

    \I__3000\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23155\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__23149\,
            I => \ALU.madd_224\
        );

    \I__2996\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23143\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__23143\,
            I => \ALU.madd_121\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23137\,
            I => \N__23134\
        );

    \I__2992\ : Odrv12
    port map (
            O => \N__23134\,
            I => \ALU.b_3_ns_1_8\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__23131\,
            I => \ALU.a_9_cascade_\
        );

    \I__2990\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23125\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__2988\ : Span4Mux_h
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__23119\,
            I => \ALU.N_675_1\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__23116\,
            I => \ALU.bZ0Z_0_cascade_\
        );

    \I__2985\ : InMux
    port map (
            O => \N__23113\,
            I => \N__23110\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23110\,
            I => \ALU.madd_130_0_0\
        );

    \I__2983\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23103\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23097\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23103\,
            I => \N__23094\
        );

    \I__2980\ : InMux
    port map (
            O => \N__23102\,
            I => \N__23091\
        );

    \I__2979\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23088\
        );

    \I__2978\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23085\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__23097\,
            I => \N__23082\
        );

    \I__2976\ : Span4Mux_v
    port map (
            O => \N__23094\,
            I => \N__23077\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23077\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__23088\,
            I => \N__23074\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23085\,
            I => \N__23071\
        );

    \I__2972\ : Span4Mux_s3_h
    port map (
            O => \N__23082\,
            I => \N__23068\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__23077\,
            I => \N__23063\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__23074\,
            I => \N__23063\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__23071\,
            I => \N__23060\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__23068\,
            I => \ALU.r6_RNIGC3D2Z0Z_7\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__23063\,
            I => \ALU.r6_RNIGC3D2Z0Z_7\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__23060\,
            I => \ALU.r6_RNIGC3D2Z0Z_7\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__23053\,
            I => \ALU.a_7_cascade_\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__23050\,
            I => \N__23046\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__23049\,
            I => \N__23043\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23038\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23038\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__23034\
        );

    \I__2959\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23031\
        );

    \I__2958\ : Span4Mux_s2_h
    port map (
            O => \N__23034\,
            I => \N__23026\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__23026\
        );

    \I__2956\ : Span4Mux_v
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__23023\,
            I => \ALU.madd_76\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__23020\,
            I => \N__23017\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__23014\,
            I => \ALU.madd_213_0_tz\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23008\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__2949\ : Span4Mux_v
    port map (
            O => \N__23005\,
            I => \N__23002\
        );

    \I__2948\ : Odrv4
    port map (
            O => \N__23002\,
            I => \ALU.madd_209_0\
        );

    \I__2947\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22996\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__22996\,
            I => \ALU.madd_223_0_tz\
        );

    \I__2945\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22990\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__2943\ : Span4Mux_s1_v
    port map (
            O => \N__22987\,
            I => \N__22984\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__22984\,
            I => \ALU.madd_105_0\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__22978\,
            I => \ALU.r4_RNIU5NK1Z0Z_8\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__22975\,
            I => \ALU.un9_addsub_axb_1_cascade_\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22969\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__22969\,
            I => \ALU.a7_b_3\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__22966\,
            I => \ALU.a_1_cascade_\
        );

    \I__2935\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22960\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__22957\,
            I => \ALU.madd_228_0_tz\
        );

    \I__2932\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__22951\,
            I => \ALU.g3\
        );

    \I__2930\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__22945\,
            I => \ALU.madd_72_0_tz\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__22942\,
            I => \ALU.madd_40_cascade_\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__2926\ : InMux
    port map (
            O => \N__22936\,
            I => \N__22930\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22930\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22930\,
            I => \ALU.madd_72\
        );

    \I__2923\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22924\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__22924\,
            I => \N__22919\
        );

    \I__2921\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22914\
        );

    \I__2920\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22914\
        );

    \I__2919\ : Odrv12
    port map (
            O => \N__22919\,
            I => \ALU.madd_95\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__22914\,
            I => \ALU.madd_95\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__22909\,
            I => \ALU.madd_72_cascade_\
        );

    \I__2916\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22901\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22896\
        );

    \I__2914\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22896\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__22901\,
            I => \ALU.madd_77\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__22896\,
            I => \ALU.madd_77\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__22891\,
            I => \ALU.b_8_cascade_\
        );

    \I__2910\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22885\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22882\
        );

    \I__2908\ : Span4Mux_s2_v
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__22879\,
            I => \ALU.madd_82\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__22876\,
            I => \ALU.madd_127_cascade_\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22868\
        );

    \I__2904\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22865\
        );

    \I__2903\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22862\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22857\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22865\,
            I => \N__22857\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__22862\,
            I => \N__22854\
        );

    \I__2899\ : Span4Mux_v
    port map (
            O => \N__22857\,
            I => \N__22851\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__22854\,
            I => \ALU.madd_223\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__22851\,
            I => \ALU.madd_223\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__22846\,
            I => \ALU.a4_b_4_cascade_\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22838\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22833\
        );

    \I__2893\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22833\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__22838\,
            I => \N__22830\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22827\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__22830\,
            I => \ALU.madd_104\
        );

    \I__2889\ : Odrv12
    port map (
            O => \N__22827\,
            I => \ALU.madd_104\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__22822\,
            I => \ALU.madd_68_cascade_\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__22819\,
            I => \ALU.madd_82_0_cascade_\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22807\
        );

    \I__2885\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22807\
        );

    \I__2884\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22807\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__22807\,
            I => \N__22804\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__22804\,
            I => \ALU.madd_119\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \ALU.a_6_cascade_\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22795\,
            I => \ALU.r0_12_prm_6_11_s0_c_RNOZ0\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__2877\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22786\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__22786\,
            I => \ALU.r0_12_prm_7_11_s0_c_RNOZ0\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__2874\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22777\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__22777\,
            I => \N__22774\
        );

    \I__2872\ : Span4Mux_v
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__22771\,
            I => \ALU.r0_12_prm_6_11_s1_c_RNOZ0\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22762\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__2867\ : Odrv4
    port map (
            O => \N__22759\,
            I => \TXbuffer_18_3_ns_1_5\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__22756\,
            I => \TXbuffer_18_10_ns_1_6_cascade_\
        );

    \I__2865\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22750\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__2863\ : Sp12to4
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__2862\ : Odrv12
    port map (
            O => \N__22744\,
            I => \TXbuffer_RNO_1Z0Z_6\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__22741\,
            I => \TXbuffer_RNO_0Z0Z_6_cascade_\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22735\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22732\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__22732\,
            I => \TXbuffer_18_6_ns_1_6\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__22729\,
            I => \TXbuffer_RNO_6Z0Z_6_cascade_\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__22723\,
            I => \TXbuffer_18_15_ns_1_6\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__22720\,
            I => \TXbuffer_18_3_ns_1_6_cascade_\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22714\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__22714\,
            I => \TXbuffer_RNO_5Z0Z_6\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__22711\,
            I => \N__22708\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22705\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22702\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__22702\,
            I => \N__22699\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__22699\,
            I => \ALU.r0_12_prm_4_11_s1_c_RNOZ0\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22693\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__22693\,
            I => \ALU.r5_RNIAFVE5Z0Z_11\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22687\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__22687\,
            I => \ALU.r0_12_prm_5_11_s0_c_RNOZ0\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22681\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__22681\,
            I => \N__22676\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22680\,
            I => \N__22673\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22670\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__22676\,
            I => \N__22667\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__22673\,
            I => \N__22662\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22670\,
            I => \N__22662\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__22667\,
            I => \N__22659\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__22662\,
            I => \N__22656\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__22659\,
            I => r7_10
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__22656\,
            I => r7_10
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__22651\,
            I => \N__22646\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22643\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22640\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22646\,
            I => \N__22637\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22643\,
            I => \N__22632\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22640\,
            I => \N__22632\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22629\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__22632\,
            I => \N__22626\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__22629\,
            I => r7_11
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__22626\,
            I => r7_11
        );

    \I__2821\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22614\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22614\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22611\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22614\,
            I => r7_15
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22611\,
            I => r7_15
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \TXbuffer_18_3_ns_1_2_cascade_\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__2812\ : Span4Mux_v
    port map (
            O => \N__22594\,
            I => \N__22591\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__22591\,
            I => \TXbuffer_RNO_5Z0Z_2\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__22588\,
            I => \N__22585\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22582\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__22582\,
            I => \N__22579\
        );

    \I__2807\ : Sp12to4
    port map (
            O => \N__22579\,
            I => \N__22576\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__22576\,
            I => \TXbuffer_18_3_ns_1_4\
        );

    \I__2805\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22569\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22565\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22569\,
            I => \N__22562\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22559\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22556\
        );

    \I__2800\ : Span4Mux_s3_h
    port map (
            O => \N__22562\,
            I => \N__22551\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22551\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__22556\,
            I => \N__22548\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__22551\,
            I => \N__22545\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__22548\,
            I => \N__22542\
        );

    \I__2795\ : Span4Mux_s3_h
    port map (
            O => \N__22545\,
            I => \N__22539\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__22542\,
            I => r6_10
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__22539\,
            I => r6_10
        );

    \I__2792\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22526\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22521\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22521\
        );

    \I__2788\ : Span4Mux_h
    port map (
            O => \N__22526\,
            I => \N__22516\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22516\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__22516\,
            I => r6_15
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__22513\,
            I => \N__22508\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22503\
        );

    \I__2783\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22503\
        );

    \I__2782\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22500\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22497\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__22500\,
            I => \N__22494\
        );

    \I__2779\ : Span4Mux_s2_h
    port map (
            O => \N__22497\,
            I => \N__22489\
        );

    \I__2778\ : Span4Mux_v
    port map (
            O => \N__22494\,
            I => \N__22489\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__22489\,
            I => r3_15
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__22486\,
            I => \N__22483\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22478\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__22482\,
            I => \N__22475\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__22481\,
            I => \N__22472\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__22478\,
            I => \N__22469\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22466\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22463\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22469\,
            I => r3_7
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__22466\,
            I => r3_7
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22463\,
            I => r3_7
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__22456\,
            I => \TXbuffer_18_13_ns_1_6_cascade_\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__22453\,
            I => \ALU.a_6_ns_1_7_cascade_\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__22450\,
            I => \ALU.b_6_ns_1_7_cascade_\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22444\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22444\,
            I => \N__22441\
        );

    \I__2761\ : Span4Mux_v
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__22438\,
            I => \ALU.r6_RNIJ13O1Z0Z_7\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22428\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22425\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__22428\,
            I => \N__22419\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22425\,
            I => \N__22419\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22416\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__22419\,
            I => r2_15
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22416\,
            I => r2_15
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22403\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22398\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22398\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__22403\,
            I => r2_7
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__22398\,
            I => r2_7
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__22393\,
            I => \TXbuffer_18_6_ns_1_7_cascade_\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22386\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__22389\,
            I => \N__22382\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22379\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22376\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22373\
        );

    \I__2739\ : Span4Mux_s3_h
    port map (
            O => \N__22379\,
            I => \N__22366\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22366\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__22373\,
            I => \N__22366\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__22366\,
            I => r3_10
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \N__22358\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22355\
        );

    \I__2733\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22352\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22349\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__22355\,
            I => \N__22346\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22343\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22340\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__22346\,
            I => r3_11
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__22343\,
            I => r3_11
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__22340\,
            I => r3_11
        );

    \I__2725\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22330\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__2723\ : Span4Mux_s3_h
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__22324\,
            I => \N__22320\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22317\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__22320\,
            I => \N__22313\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__22317\,
            I => \N__22310\
        );

    \I__2718\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22307\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__22313\,
            I => r0_5
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__22310\,
            I => r0_5
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__22307\,
            I => r0_5
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__22300\,
            I => \ALU.a_3_ns_1_5_cascade_\
        );

    \I__2713\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22294\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__2711\ : Span4Mux_s2_h
    port map (
            O => \N__22291\,
            I => \N__22286\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22283\
        );

    \I__2709\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22280\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__22286\,
            I => r2_10
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22283\,
            I => r2_10
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__22280\,
            I => r2_10
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__22273\,
            I => \ALU.a_6_ns_1_10_cascade_\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__22270\,
            I => \ALU.a_6_ns_1_11_cascade_\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__22267\,
            I => \ALU.r6_RNIT7372Z0Z_11_cascade_\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__22264\,
            I => \ALU.b_5_cascade_\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__22261\,
            I => \TXbuffer_18_3_ns_1_1_cascade_\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__22258\,
            I => \TXbuffer_RNO_5Z0Z_1_cascade_\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22250\
        );

    \I__2698\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22245\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22245\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__22250\,
            I => r6_9
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__22245\,
            I => r6_9
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__22240\,
            I => \TXbuffer_18_6_ns_1_1_cascade_\
        );

    \I__2693\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__22234\,
            I => \TXbuffer_RNO_6Z0Z_1\
        );

    \I__2691\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22228\,
            I => \N__22221\
        );

    \I__2689\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22212\
        );

    \I__2688\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22212\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22212\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22212\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__22221\,
            I => \ALU.madd_213\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__22212\,
            I => \ALU.madd_213\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22202\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22197\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22197\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22194\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22197\,
            I => \ALU.a9_b_3\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__22194\,
            I => \ALU.a9_b_3\
        );

    \I__2677\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__22186\,
            I => \N__22183\
        );

    \I__2675\ : Span4Mux_s1_h
    port map (
            O => \N__22183\,
            I => \N__22180\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__22180\,
            I => \N__22177\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__22177\,
            I => \ALU.madd_167_0\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__22174\,
            I => \ALU.b_6_ns_1_5_cascade_\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__22171\,
            I => \ALU.b_3_ns_1_5_cascade_\
        );

    \I__2670\ : InMux
    port map (
            O => \N__22168\,
            I => \N__22165\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__22165\,
            I => \ALU.r6_RNIBP2O1Z0Z_5\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__22162\,
            I => \ALU.r4_RNI0QNE1Z0Z_5_cascade_\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22154\
        );

    \I__2666\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22149\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22149\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__22154\,
            I => \N__22146\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__22149\,
            I => \N__22143\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__22146\,
            I => \N__22138\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__22143\,
            I => \N__22138\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__22138\,
            I => \ALU.a0_b_14\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__22132\,
            I => \ALU.g2_0\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__22126\,
            I => \ALU.g0_2_N_4L5\
        );

    \I__2655\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22117\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22117\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__22117\,
            I => \N__22114\
        );

    \I__2652\ : Span4Mux_h
    port map (
            O => \N__22114\,
            I => \N__22110\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22107\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__22110\,
            I => \ALU.madd_134_0_tz\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22107\,
            I => \ALU.madd_134_0_tz\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22099\,
            I => \ALU.madd_130_0\
        );

    \I__2646\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__22093\,
            I => \N__22088\
        );

    \I__2644\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22083\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22083\
        );

    \I__2642\ : Span4Mux_s1_v
    port map (
            O => \N__22088\,
            I => \N__22080\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__22083\,
            I => \N__22077\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__22080\,
            I => \N__22074\
        );

    \I__2639\ : Span4Mux_s1_v
    port map (
            O => \N__22077\,
            I => \N__22071\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__22074\,
            I => \ALU.madd_130\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__22071\,
            I => \ALU.madd_130\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__22066\,
            I => \N__22063\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__2633\ : Span4Mux_s1_h
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__22054\,
            I => \ALU.madd_171_sx\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__22048\,
            I => \ALU.a5_b_8\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__22045\,
            I => \N__22042\
        );

    \I__2628\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22036\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22036\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__22036\,
            I => \ALU.a6_b_7\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22029\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22026\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__22029\,
            I => \N__22021\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__22021\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__22021\,
            I => \ALU.madd_321\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__22018\,
            I => \ALU.b_6_ns_1_6_cascade_\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__22015\,
            I => \ALU.r6_RNIIH042Z0Z_6_cascade_\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__22012\,
            I => \ALU.b_6_cascade_\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__22003\,
            I => \ALU.g0_2_N_3L3\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__22000\,
            I => \N__21996\
        );

    \I__2613\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21986\
        );

    \I__2612\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21986\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__21995\,
            I => \N__21981\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__21994\,
            I => \N__21976\
        );

    \I__2609\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21971\
        );

    \I__2608\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21971\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__21991\,
            I => \N__21965\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21960\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21947\
        );

    \I__2604\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21947\
        );

    \I__2603\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21947\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21947\
        );

    \I__2601\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21947\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21947\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21944\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21936\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21936\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21936\
        );

    \I__2595\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21929\
        );

    \I__2594\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21929\
        );

    \I__2593\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21926\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__21960\,
            I => \N__21921\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21921\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__21944\,
            I => \N__21918\
        );

    \I__2589\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21915\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__21936\,
            I => \N__21912\
        );

    \I__2587\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21907\
        );

    \I__2586\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21907\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__21929\,
            I => \bZ0Z_2\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__21926\,
            I => \bZ0Z_2\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__21921\,
            I => \bZ0Z_2\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__21918\,
            I => \bZ0Z_2\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__21915\,
            I => \bZ0Z_2\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__21912\,
            I => \bZ0Z_2\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__21907\,
            I => \bZ0Z_2\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__21892\,
            I => \ALU.b_3_ns_1_6_cascade_\
        );

    \I__2577\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21886\,
            I => \ALU.r4_RNIAP7R1Z0Z_6\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__21880\,
            I => \N__21877\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__21877\,
            I => \ALU.madd_144_0_tz\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21868\
        );

    \I__2571\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21865\
        );

    \I__2570\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21860\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21860\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__21868\,
            I => \N__21857\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__21865\,
            I => \ALU.a4_b_5\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21860\,
            I => \ALU.a4_b_5\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__21857\,
            I => \ALU.a4_b_5\
        );

    \I__2564\ : InMux
    port map (
            O => \N__21850\,
            I => \N__21847\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21844\
        );

    \I__2562\ : Span4Mux_s0_v
    port map (
            O => \N__21844\,
            I => \N__21841\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__21841\,
            I => \ALU.g0_6_1\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21835\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__21835\,
            I => \N__21831\
        );

    \I__2558\ : InMux
    port map (
            O => \N__21834\,
            I => \N__21828\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__21831\,
            I => \N__21825\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21822\
        );

    \I__2555\ : Odrv4
    port map (
            O => \N__21825\,
            I => \ALU.r6_RNIUC0U1Z0Z_10\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__21822\,
            I => \ALU.r6_RNIUC0U1Z0Z_10\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21814\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__21811\,
            I => \N__21807\
        );

    \I__2550\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21804\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__21807\,
            I => \ALU.r5_RNIMCFS1Z0Z_10\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__21804\,
            I => \ALU.r5_RNIMCFS1Z0Z_10\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21796\,
            I => \ALU.a0_b_10\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__21793\,
            I => \ALU.a5_b_8_cascade_\
        );

    \I__2544\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21783\
        );

    \I__2542\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21780\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__21783\,
            I => \N__21777\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21774\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__21777\,
            I => \N__21771\
        );

    \I__2538\ : Span4Mux_s3_h
    port map (
            O => \N__21774\,
            I => \N__21768\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__21771\,
            I => \ALU.madd_325\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__21768\,
            I => \ALU.madd_325\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__21763\,
            I => \ALU.b_7_cascade_\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__21760\,
            I => \N__21756\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21753\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21750\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21753\,
            I => \ALU.a5_b_7\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21750\,
            I => \ALU.a5_b_7\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__21745\,
            I => \ALU.a5_b_5_cascade_\
        );

    \I__2528\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21736\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21736\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__21736\,
            I => \N__21731\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21726\
        );

    \I__2524\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21726\
        );

    \I__2523\ : Span4Mux_s2_v
    port map (
            O => \N__21731\,
            I => \N__21721\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21721\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__21721\,
            I => \ALU.madd_176\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__21718\,
            I => \ALU.madd_43_0_cascade_\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__21712\,
            I => \ALU.madd_77_0_tz\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21705\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21702\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21705\,
            I => \N__21699\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__21702\,
            I => \N__21696\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__21699\,
            I => \ALU.madd_278\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__21696\,
            I => \ALU.madd_278\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21688\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21688\,
            I => \N__21684\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21687\,
            I => \N__21681\
        );

    \I__2508\ : Span4Mux_s3_h
    port map (
            O => \N__21684\,
            I => \N__21678\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__21681\,
            I => \ALU.madd_273\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__21678\,
            I => \ALU.madd_273\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__21673\,
            I => \N__21669\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21665\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21662\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21659\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21656\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__21662\,
            I => \N__21653\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21650\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__21656\,
            I => \N__21647\
        );

    \I__2497\ : Span4Mux_s3_h
    port map (
            O => \N__21653\,
            I => \N__21642\
        );

    \I__2496\ : Span4Mux_s3_h
    port map (
            O => \N__21650\,
            I => \N__21642\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__21647\,
            I => \N__21639\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__21642\,
            I => \N__21636\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__21639\,
            I => \ALU.madd_345\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__21636\,
            I => \ALU.madd_345\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__21628\,
            I => \ALU.madd_159_N_3L3\
        );

    \I__2489\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__21622\,
            I => \ALU.madd_61\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__2486\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21613\,
            I => \ALU.madd_140_0\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__21610\,
            I => \ALU.madd_140_0_cascade_\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21604\,
            I => \ALU.madd_155_1\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21597\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__21600\,
            I => \N__21594\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21597\,
            I => \N__21591\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21588\
        );

    \I__2477\ : Odrv12
    port map (
            O => \N__21591\,
            I => \ALU.a_i_11\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__21588\,
            I => \ALU.a_i_11\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21580\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21580\,
            I => \ALU.r0_12_prm_3_11_s0_sf\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21577\,
            I => \ALU.r0_12_s0_11\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21571\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__21565\,
            I => \ALU.r0_12_s0_11_THRU_CO\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__21562\,
            I => \ALU.g1_7_cascade_\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21556\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__21556\,
            I => \ALU.a4_b_0_0_5\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__21553\,
            I => \ALU.N_663_0_cascade_\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21543\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21543\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21540\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21543\,
            I => \ALU.madd_109\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__21540\,
            I => \ALU.madd_109\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21532\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__21529\,
            I => \ALU.N_683_0_0_0\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \TXbuffer_18_6_ns_1_0_cascade_\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21520\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__21520\,
            I => \N__21517\
        );

    \I__2453\ : Span4Mux_s2_h
    port map (
            O => \N__21517\,
            I => \N__21514\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__21514\,
            I => \TXbuffer_RNO_6Z0Z_0\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21508\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__21502\,
            I => \TXbuffer_18_13_ns_1_7\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21495\
        );

    \I__2446\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21492\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21495\,
            I => \N__21489\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__21492\,
            I => \N__21486\
        );

    \I__2443\ : Span4Mux_h
    port map (
            O => \N__21489\,
            I => \N__21483\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__21486\,
            I => \ALU.r5_RNIE0AK8_0Z0Z_11\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__21483\,
            I => \ALU.r5_RNIE0AK8_0Z0Z_11\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21472\,
            I => \N__21468\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21465\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__21468\,
            I => \N__21462\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21465\,
            I => \ALU.r5_RNIE0AK8_1Z0Z_11\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__21462\,
            I => \ALU.r5_RNIE0AK8_1Z0Z_11\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__21457\,
            I => \ALU.b_6_ns_1_12_cascade_\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21451\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21451\,
            I => \N__21448\
        );

    \I__2430\ : Odrv12
    port map (
            O => \N__21448\,
            I => \ALU.r6_RNI85GA2Z0Z_12\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21442\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__21442\,
            I => \N__21439\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__21439\,
            I => \N__21435\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21432\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__21435\,
            I => \ALU.r5_RNI05V82Z0Z_12\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__21432\,
            I => \ALU.r5_RNI05V82Z0Z_12\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__21427\,
            I => \ALU.r6_RNI85GA2Z0Z_12_cascade_\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__21424\,
            I => \ALU.b_3_ns_1_13_cascade_\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21418\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21418\,
            I => \ALU.r5_RNI49V82Z0Z_13\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__21415\,
            I => \ALU.a_6_ns_1_15_cascade_\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21409\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21409\,
            I => \ALU.r6_RNIH8772Z0Z_15\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21403\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__21403\,
            I => \N__21400\
        );

    \I__2414\ : Span4Mux_s3_h
    port map (
            O => \N__21400\,
            I => \N__21397\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__21397\,
            I => \ALU.r6_RNINRNUZ0Z_15\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__21394\,
            I => \N__21391\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21388\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21388\,
            I => \ALU.r0_12_prm_1_11_s1_c_RNOZ0\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21385\,
            I => \ALU.r0_12_s1_11\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__21382\,
            I => \ALU.b_3_ns_1_12_cascade_\
        );

    \I__2407\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21376\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__21376\,
            I => \ALU.r5_RNIH9VTZ0Z_14\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__21373\,
            I => \ALU.r1_RNI8DSRZ0Z_14_cascade_\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21367\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__21367\,
            I => \ALU.r2_RNIDP6TZ0Z_14\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__21364\,
            I => \ALU.b_7_ns_1_14_cascade_\
        );

    \I__2401\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21358\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21358\,
            I => \ALU.r6_RNILPNUZ0Z_14\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__21355\,
            I => \ALU.b_14_cascade_\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__21352\,
            I => \N__21349\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21346\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21346\,
            I => \N__21343\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__21343\,
            I => \ALU.r0_12_prm_7_11_s1_c_RNOZ0\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__21340\,
            I => \N__21337\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21337\,
            I => \N__21334\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21334\,
            I => \N__21331\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__21331\,
            I => \ALU.r0_12_prm_5_11_s1_c_RNOZ0\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__21328\,
            I => \ALU.b_6_ns_1_11_cascade_\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21322\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__21322\,
            I => \N__21319\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__21319\,
            I => \ALU.r6_RNI2H0U1Z0Z_11\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__21316\,
            I => \ALU.b_6_ns_1_9_cascade_\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21310\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__21310\,
            I => \N__21307\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__21307\,
            I => \N__21303\
        );

    \I__2382\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21300\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__21303\,
            I => \ALU.r6_RNIUT042Z0Z_9\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__21300\,
            I => \ALU.r6_RNIUT042Z0Z_9\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \ALU.b_3_ns_1_9_cascade_\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21289\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21289\,
            I => \N__21285\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21282\
        );

    \I__2375\ : Odrv12
    port map (
            O => \N__21285\,
            I => \ALU.r4_RNIM58R1Z0Z_9\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21282\,
            I => \ALU.r4_RNIM58R1Z0Z_9\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__21277\,
            I => \ALU.b_3_ns_1_10_cascade_\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__21274\,
            I => \ALU.b_3_ns_1_11_cascade_\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__21271\,
            I => \ALU.r5_RNIQGFS1Z0Z_11_cascade_\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__21268\,
            I => \ALU.b_6_ns_1_10_cascade_\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__21265\,
            I => \ALU.a12_b_0_cascade_\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21258\
        );

    \I__2367\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21255\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21250\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__21255\,
            I => \N__21250\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__21250\,
            I => \ALU.madd_263\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__21247\,
            I => \ALU.madd_264_cascade_\
        );

    \I__2362\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21238\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21238\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21238\,
            I => \ALU.madd_288\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21232\,
            I => \ALU.a12_b_0\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__21229\,
            I => \N__21225\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21220\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21220\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__21220\,
            I => \ALU.a10_b_2\
        );

    \I__2353\ : InMux
    port map (
            O => \N__21217\,
            I => \N__21214\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21214\,
            I => \ALU.madd_259\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__21211\,
            I => \N__21207\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21203\
        );

    \I__2349\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21198\
        );

    \I__2348\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21198\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N__21195\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__21198\,
            I => \ALU.a7_b_5\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__21195\,
            I => \ALU.a7_b_5\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__21190\,
            I => \ALU.madd_259_cascade_\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__21187\,
            I => \N__21184\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21180\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21177\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__21180\,
            I => \N__21174\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21171\
        );

    \I__2338\ : Span4Mux_s2_h
    port map (
            O => \N__21174\,
            I => \N__21166\
        );

    \I__2337\ : Span4Mux_s3_v
    port map (
            O => \N__21171\,
            I => \N__21166\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__21166\,
            I => \ALU.madd_284_0\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21154\
        );

    \I__2334\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21154\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21154\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21154\,
            I => \ALU.madd_336\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__21151\,
            I => \N__21147\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__21150\,
            I => \N__21144\
        );

    \I__2329\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21136\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21136\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21136\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__21136\,
            I => \N__21133\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__21133\,
            I => \ALU.madd_335\
        );

    \I__2324\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21127\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__21127\,
            I => \ALU.madd_283\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21121\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21118\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__21118\,
            I => \ALU.madd_124_0\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__21115\,
            I => \N__21112\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21109\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__21109\,
            I => \N__21106\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__21106\,
            I => \ALU.madd_218_0_tz\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__21103\,
            I => \ALU.madd_218_cascade_\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21097\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21097\,
            I => \ALU.madd_346_1\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21088\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21088\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__21088\,
            I => \N__21085\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__21085\,
            I => \ALU.a2_b_10\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__21082\,
            I => \ALU.a0_b_12_cascade_\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21075\
        );

    \I__2306\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21072\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21075\,
            I => \N__21069\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__21072\,
            I => \ALU.madd_279_0\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__21069\,
            I => \ALU.madd_279_0\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21060\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21056\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21060\,
            I => \N__21053\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21050\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__21056\,
            I => \ALU.madd_331_0\
        );

    \I__2297\ : Odrv12
    port map (
            O => \N__21053\,
            I => \ALU.madd_331_0\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__21050\,
            I => \ALU.madd_331_0\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__21043\,
            I => \N__21040\
        );

    \I__2294\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21037\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__21037\,
            I => \N__21033\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__21036\,
            I => \N__21030\
        );

    \I__2291\ : Span4Mux_s2_h
    port map (
            O => \N__21033\,
            I => \N__21025\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21022\
        );

    \I__2289\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21017\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21028\,
            I => \N__21017\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__21025\,
            I => \ALU.a0_b_12\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__21022\,
            I => \ALU.a0_b_12\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__21017\,
            I => \ALU.a0_b_12\
        );

    \I__2284\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21003\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21009\,
            I => \N__21003\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21008\,
            I => \N__20998\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__20995\
        );

    \I__2280\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20990\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20990\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__20998\,
            I => \ALU.madd_218\
        );

    \I__2277\ : Odrv12
    port map (
            O => \N__20995\,
            I => \ALU.madd_218\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20990\,
            I => \ALU.madd_218\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20979\
        );

    \I__2274\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20976\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__20979\,
            I => \ALU.madd_202\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__20976\,
            I => \ALU.madd_202\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20967\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20964\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__20967\,
            I => \ALU.madd_228\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__20964\,
            I => \ALU.madd_228\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20956\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20952\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20955\,
            I => \N__20949\
        );

    \I__2264\ : Odrv12
    port map (
            O => \N__20952\,
            I => \ALU.madd_338\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__20949\,
            I => \ALU.madd_338\
        );

    \I__2262\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20941\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20941\,
            I => \N__20937\
        );

    \I__2260\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20934\
        );

    \I__2259\ : Odrv12
    port map (
            O => \N__20937\,
            I => \ALU.madd_337\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__20934\,
            I => \ALU.madd_337\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20926\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20926\,
            I => \ALU.a0_b_13\
        );

    \I__2255\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20919\
        );

    \I__2254\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20916\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__20919\,
            I => \ALU.madd_335_0\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__20916\,
            I => \ALU.madd_335_0\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20908\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__20908\,
            I => \N__20904\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20901\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__20904\,
            I => \ALU.madd_233\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__20901\,
            I => \ALU.madd_233\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__20896\,
            I => \N__20893\
        );

    \I__2245\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20889\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__20892\,
            I => \N__20886\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20882\
        );

    \I__2242\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20877\
        );

    \I__2241\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20877\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__20882\,
            I => \N__20874\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20877\,
            I => \N__20871\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__20874\,
            I => \ALU.madd_238\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__20871\,
            I => \ALU.madd_238\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20860\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20860\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__20860\,
            I => \ALU.madd_294\
        );

    \I__2233\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20852\
        );

    \I__2232\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20849\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20846\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__20852\,
            I => \ALU.madd_304\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__20849\,
            I => \ALU.madd_304\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__20846\,
            I => \ALU.madd_304\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20833\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20833\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20829\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20832\,
            I => \N__20826\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__20829\,
            I => \ALU.madd_253\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__20826\,
            I => \ALU.madd_253\
        );

    \I__2221\ : InMux
    port map (
            O => \N__20821\,
            I => \N__20817\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__20820\,
            I => \N__20814\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__20817\,
            I => \N__20811\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20808\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__20811\,
            I => \ALU.madd_341\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__20808\,
            I => \ALU.madd_341\
        );

    \I__2215\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20800\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20800\,
            I => \ALU.a4_b_8\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__20797\,
            I => \ALU.a4_b_8_cascade_\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20791\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__20791\,
            I => \ALU.madd_269\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__20788\,
            I => \N__20784\
        );

    \I__2209\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20781\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20778\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__20781\,
            I => \ALU.madd_274\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20778\,
            I => \ALU.madd_274\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__20773\,
            I => \ALU.madd_269_cascade_\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20765\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20760\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20760\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20757\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__20760\,
            I => \ALU.madd_289\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__20757\,
            I => \ALU.madd_289\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__20752\,
            I => \ALU.madd_185_1_cascade_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20743\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__20743\,
            I => \N__20740\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__20740\,
            I => \ALU.madd_106\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__20737\,
            I => \ALU.g0_2_N_2L1_cascade_\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__20734\,
            I => \N__20731\
        );

    \I__2191\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20725\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20725\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__20725\,
            I => \ALU.madd_186_0\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20715\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20712\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__20715\,
            I => \ALU.a6_b_2\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__20712\,
            I => \ALU.a6_b_2\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__20707\,
            I => \ALU.a6_b_2_cascade_\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20700\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20697\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20700\,
            I => \ALU.a7_b_1\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__20697\,
            I => \ALU.a7_b_1\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__20692\,
            I => \ALU.madd_99_cascade_\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20681\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20681\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20676\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20676\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20681\,
            I => \ALU.madd_149\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__20676\,
            I => \ALU.madd_149\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20668\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__20668\,
            I => \ALU.madd_99\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20659\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20659\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20659\,
            I => \ALU.madd_145\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20653\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20653\,
            I => \ALU.madd_244\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \N__20647\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20644\,
            I => \ALU.madd_201\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20636\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20633\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20630\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20636\,
            I => \N__20627\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20633\,
            I => \ALU.madd_239\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__20630\,
            I => \ALU.madd_239\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__20627\,
            I => \ALU.madd_239\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__20620\,
            I => \ALU.a3_b_9_cascade_\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20614\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20614\,
            I => \ALU.a3_b_9\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__20611\,
            I => \ALU.madd_155_cascade_\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__20608\,
            I => \ALU.madd_109_0_tz_cascade_\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__20605\,
            I => \ALU.madd_109_cascade_\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20599\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20599\,
            I => \ALU.N_687_0\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20593\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20590\
        );

    \I__2144\ : Span4Mux_s0_v
    port map (
            O => \N__20590\,
            I => \N__20587\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__20587\,
            I => \ALU.madd_159_N_2L1\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20575\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20575\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__20575\,
            I => \ALU.madd_159\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \N__20569\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20563\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20563\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20560\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__20560\,
            I => \ALU.madd_150\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20551\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20551\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20551\,
            I => \ALU.madd_155\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__20548\,
            I => \ALU.a7_b_1_cascade_\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__20545\,
            I => \ALU.r6_RNIC9GA2Z0Z_13_cascade_\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__20542\,
            I => \ALU.b_13_cascade_\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__20539\,
            I => \TXbuffer_18_13_ns_1_4_cascade_\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20533\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20533\,
            I => \N__20530\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__20530\,
            I => \N__20527\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__20527\,
            I => \TXbuffer_RNO_1Z0Z_4\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__20524\,
            I => \N__20521\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20518\,
            I => \N__20515\
        );

    \I__2119\ : Odrv12
    port map (
            O => \N__20515\,
            I => \ALU.N_661_0\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__20512\,
            I => \ALU.a_15_cascade_\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__20509\,
            I => \ALU.lshift_3_ns_1_15_cascade_\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__20506\,
            I => \ALU.b_6_ns_1_13_cascade_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20497\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__20497\,
            I => \TXbuffer_18_13_ns_1_3\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__20491\,
            I => \ALU.r1_RNIAFSRZ0Z_15\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__20488\,
            I => \ALU.r5_RNIJBVTZ0Z_15_cascade_\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20482\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20482\,
            I => \ALU.b_7_ns_1_15\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20476\,
            I => \N__20473\
        );

    \I__2105\ : Span4Mux_v
    port map (
            O => \N__20473\,
            I => \N__20470\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__20467\,
            I => \ALU.madd_490_1\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__2100\ : Span4Mux_v
    port map (
            O => \N__20458\,
            I => \N__20455\
        );

    \I__2099\ : Span4Mux_s1_h
    port map (
            O => \N__20455\,
            I => \N__20452\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__20452\,
            I => \ALU.madd_490_9\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__20449\,
            I => \ALU.madd_490_0_cascade_\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20443\,
            I => \ALU.madd_490_13\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20437\,
            I => \N__20434\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__20434\,
            I => \ALU.madd_490_14\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__20431\,
            I => \ALU.r2_RNIFR6TZ0Z_15_cascade_\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__20428\,
            I => \ALU.b_15_cascade_\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20422\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__20422\,
            I => \N__20418\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20415\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__20418\,
            I => \ALU.a5_b_9\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__20415\,
            I => \ALU.a5_b_9\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__20410\,
            I => \ALU.a6_b_8_cascade_\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20401\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20401\,
            I => \N__20398\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__20398\,
            I => \ALU.madd_378\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__20395\,
            I => \ALU.b_i_3_cascade_\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__2076\ : Odrv12
    port map (
            O => \N__20386\,
            I => \ALU.a3_b_11\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__20380\,
            I => \ALU.madd_382\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20370\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20367\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__20370\,
            I => \ALU.a4_b_10\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20367\,
            I => \ALU.a4_b_10\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__20362\,
            I => \ALU.a11_b_3_cascade_\
        );

    \I__2067\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20356\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20356\,
            I => \ALU.madd_373\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__20353\,
            I => \N__20350\
        );

    \I__2064\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20347\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__20347\,
            I => \ALU.a11_b_3\
        );

    \I__2062\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20341\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20338\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__20338\,
            I => \N__20335\
        );

    \I__2059\ : Span4Mux_s0_h
    port map (
            O => \N__20335\,
            I => \N__20332\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__20332\,
            I => \ALU.madd_392\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20326\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20326\,
            I => \ALU.madd_490_16\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__20323\,
            I => \ALU.madd_490_15_cascade_\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20317\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20317\,
            I => \ALU.madd_490_19\
        );

    \I__2052\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20311\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__20311\,
            I => \N__20308\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__20308\,
            I => \N__20305\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__20305\,
            I => \ALU.madd_339\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__20302\,
            I => \N__20299\
        );

    \I__2047\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20296\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__20296\,
            I => \ALU.madd_340_0\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__20293\,
            I => \ALU.a7_b_7_cascade_\
        );

    \I__2044\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20287\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20282\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20277\
        );

    \I__2041\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20277\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__20282\,
            I => \ALU.madd_383\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__20277\,
            I => \ALU.madd_383\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__20272\,
            I => \ALU.b_9_cascade_\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__20269\,
            I => \N__20266\
        );

    \I__2036\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__20263\,
            I => \ALU.madd_326_0\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__20260\,
            I => \ALU.a5_b_9_cascade_\
        );

    \I__2033\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20254\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__20254\,
            I => \N__20251\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__20251\,
            I => \ALU.a6_b_8\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20242\
        );

    \I__2029\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20242\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__20242\,
            I => \ALU.madd_413_0\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__20239\,
            I => \ALU.madd_418_cascade_\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__20236\,
            I => \N__20233\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20227\
        );

    \I__2024\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20227\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__20224\,
            I => \ALU.madd_293\
        );

    \I__2021\ : InMux
    port map (
            O => \N__20221\,
            I => \N__20215\
        );

    \I__2020\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20215\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__20215\,
            I => \ALU.madd_336_0\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20208\
        );

    \I__2017\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20205\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__20208\,
            I => \ALU.madd_351\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__20205\,
            I => \ALU.madd_351\
        );

    \I__2014\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__20197\,
            I => \ALU.madd_346\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20190\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20187\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__20190\,
            I => \ALU.madd_172\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__20187\,
            I => \ALU.madd_172\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__20182\,
            I => \ALU.madd_346_cascade_\
        );

    \I__2007\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20175\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20172\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__20175\,
            I => \ALU.madd_298_0\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20172\,
            I => \ALU.madd_298_0\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20161\
        );

    \I__2002\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20161\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__20161\,
            I => \ALU.madd_360\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20155\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20155\,
            I => \ALU.madd_190\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__20152\,
            I => \N__20149\
        );

    \I__1997\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20146\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__20146\,
            I => \ALU.madd_330_0_tz\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20140\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20140\,
            I => \ALU.madd_326\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__20137\,
            I => \ALU.madd_326_cascade_\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20131\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20131\,
            I => \ALU.madd_350_0\
        );

    \I__1990\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20125\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__20125\,
            I => \ALU.madd_355\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20118\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20115\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__20118\,
            I => \ALU.madd_408\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20115\,
            I => \ALU.madd_408\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__20110\,
            I => \ALU.madd_350_0_cascade_\
        );

    \I__1983\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20104\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20101\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__20101\,
            I => \ALU.madd_422\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20095\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__20095\,
            I => \ALU.madd_356\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20083\
        );

    \I__1976\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20083\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__20083\,
            I => \ALU.madd_303_0\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__20080\,
            I => \ALU.madd_356_cascade_\
        );

    \I__1973\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20071\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20071\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20071\,
            I => \ALU.madd_175\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20065\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20065\,
            I => \N__20062\
        );

    \I__1968\ : Span4Mux_s2_h
    port map (
            O => \N__20062\,
            I => \N__20059\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__20059\,
            I => \ALU.madd_388_0\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20053\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__20053\,
            I => \N__20050\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__20050\,
            I => \ALU.madd_393\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20044\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__20044\,
            I => \N__20040\
        );

    \I__1961\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20037\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__20040\,
            I => \N__20032\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20032\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__20032\,
            I => \ALU.madd_340\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__20029\,
            I => \ALU.madd_355_cascade_\
        );

    \I__1956\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20023\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__20023\,
            I => \ALU.madd_418\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__20020\,
            I => \N__20017\
        );

    \I__1953\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20010\
        );

    \I__1951\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20007\
        );

    \I__1950\ : Odrv12
    port map (
            O => \N__20010\,
            I => \ALU.madd_181_0\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__20007\,
            I => \ALU.madd_181_0\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__20002\,
            I => \N__19999\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19995\
        );

    \I__1946\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19992\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__19995\,
            I => \N__19989\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19986\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__19989\,
            I => \N__19983\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__19986\,
            I => \ALU.madd_315_0\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__19983\,
            I => \ALU.madd_315_0\
        );

    \I__1940\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19974\
        );

    \I__1939\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19971\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19968\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__19971\,
            I => \N__19965\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__19968\,
            I => \ALU.madd_320\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__19965\,
            I => \ALU.madd_320\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__19960\,
            I => \ALU.madd_393_cascade_\
        );

    \I__1933\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19954\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__19948\,
            I => \ALU.madd_412\
        );

    \I__1929\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19939\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19939\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19936\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__19936\,
            I => \ALU.madd_308_0_tz_0\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__1924\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19924\
        );

    \I__1923\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19924\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__19924\,
            I => \ALU.madd_299\
        );

    \I__1921\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19917\
        );

    \I__1920\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19914\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__19917\,
            I => \ALU.madd_209\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__19914\,
            I => \ALU.madd_209\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19903\
        );

    \I__1916\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19903\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__19903\,
            I => \ALU.madd_243\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__19900\,
            I => \ALU.a0_b_13_cascade_\
        );

    \I__1913\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19891\
        );

    \I__1911\ : Sp12to4
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__19888\,
            I => \ALU.g2_0_1\
        );

    \I__1909\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19880\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__19884\,
            I => \N__19877\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__19883\,
            I => \N__19874\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19871\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19866\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19866\
        );

    \I__1903\ : Span4Mux_s1_v
    port map (
            O => \N__19871\,
            I => \N__19863\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__19866\,
            I => \N__19860\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__19863\,
            I => \ALU.madd_182_0\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__19860\,
            I => \ALU.madd_182_0\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__19855\,
            I => \N__19851\
        );

    \I__1898\ : InMux
    port map (
            O => \N__19854\,
            I => \N__19847\
        );

    \I__1897\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19842\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19842\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19847\,
            I => \ALU.a3_b_7\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__19842\,
            I => \ALU.a3_b_7\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__19837\,
            I => \N__19834\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19830\
        );

    \I__1891\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19827\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__19830\,
            I => \N__19824\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__19827\,
            I => \ALU.a2_b_8\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__19824\,
            I => \ALU.a2_b_8\
        );

    \I__1887\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19816\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19810\
        );

    \I__1885\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19803\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19803\
        );

    \I__1883\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19803\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__19810\,
            I => \ALU.madd_177\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19803\,
            I => \ALU.madd_177\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19792\
        );

    \I__1879\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19792\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__19792\,
            I => \ALU.madd_229\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__19789\,
            I => \ALU.madd_243_cascade_\
        );

    \I__1876\ : InMux
    port map (
            O => \N__19786\,
            I => \N__19778\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19778\
        );

    \I__1874\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19773\
        );

    \I__1873\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19773\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__19778\,
            I => \ALU.madd_219_0\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19773\,
            I => \ALU.madd_219_0\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__19768\,
            I => \N__19764\
        );

    \I__1869\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19759\
        );

    \I__1868\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19759\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__19759\,
            I => \ALU.madd_192_0\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19747\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19747\
        );

    \I__1864\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19747\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__19747\,
            I => \ALU.madd_144\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19741\,
            I => \ALU.g0_1\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__19738\,
            I => \N__19735\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19732\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__19729\,
            I => \ALU.N_695_0\
        );

    \I__1856\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19723\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__19723\,
            I => \ALU.g0_4\
        );

    \I__1854\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19714\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19714\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__19714\,
            I => \ALU.madd_197\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19707\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19704\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19707\,
            I => \ALU.madd_112\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__19704\,
            I => \ALU.madd_112\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19692\
        );

    \I__1846\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19692\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19689\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__19692\,
            I => \N__19686\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19689\,
            I => \ALU.madd_191\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__19686\,
            I => \ALU.madd_191\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__19675\,
            I => \ALU.madd_234\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__19672\,
            I => \ALU.madd_112_cascade_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19665\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19660\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19657\
        );

    \I__1834\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19654\
        );

    \I__1833\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19651\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19660\,
            I => \ALU.madd_196_0\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__19657\,
            I => \ALU.madd_196_0\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__19654\,
            I => \ALU.madd_196_0\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19651\,
            I => \ALU.madd_196_0\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19636\
        );

    \I__1827\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19631\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19631\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19628\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19636\,
            I => \ALU.madd_187\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__19631\,
            I => \ALU.madd_187\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19628\,
            I => \ALU.madd_187\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19615\
        );

    \I__1820\ : InMux
    port map (
            O => \N__19620\,
            I => \N__19615\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__19615\,
            I => \ALU.madd_154\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19606\
        );

    \I__1817\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19606\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19606\,
            I => \ALU.madd_134\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19603\,
            I => clkdiv_cry_22
        );

    \I__1814\ : IoInMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19594\
        );

    \I__1812\ : Span12Mux_s8_v
    port map (
            O => \N__19594\,
            I => \N__19590\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19587\
        );

    \I__1810\ : Odrv12
    port map (
            O => \N__19590\,
            I => \GPIO3_c\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19587\,
            I => \GPIO3_c\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__19582\,
            I => \ALU.madd_154_cascade_\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__19579\,
            I => \ALU.N_703_1_cascade_\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__19576\,
            I => \ALU.g0_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19573\,
            I => \N__19567\
        );

    \I__1804\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19567\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__19567\,
            I => \ALU.madd_206\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__19564\,
            I => \ALU.madd_334_cascade_\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19558\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19558\,
            I => \ALU.N_724_0_0_0\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19552\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__19552\,
            I => \clkdivZ0Z_14\
        );

    \I__1797\ : InMux
    port map (
            O => \N__19549\,
            I => clkdiv_cry_13
        );

    \I__1796\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19543\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19543\,
            I => \clkdivZ0Z_15\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19540\,
            I => clkdiv_cry_14
        );

    \I__1793\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19534\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19534\,
            I => \clkdivZ0Z_16\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19531\,
            I => \bfn_1_17_0_\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19525\,
            I => \clkdivZ0Z_17\
        );

    \I__1788\ : InMux
    port map (
            O => \N__19522\,
            I => clkdiv_cry_16
        );

    \I__1787\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19516\,
            I => \clkdivZ0Z_18\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19513\,
            I => clkdiv_cry_17
        );

    \I__1784\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19507\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19507\,
            I => \clkdivZ0Z_19\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19504\,
            I => clkdiv_cry_18
        );

    \I__1781\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19498\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__19498\,
            I => \clkdivZ0Z_20\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19495\,
            I => clkdiv_cry_19
        );

    \I__1778\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19489\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19489\,
            I => \clkdivZ0Z_21\
        );

    \I__1776\ : InMux
    port map (
            O => \N__19486\,
            I => clkdiv_cry_20
        );

    \I__1775\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19480\,
            I => \clkdivZ0Z_22\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19477\,
            I => clkdiv_cry_21
        );

    \I__1772\ : InMux
    port map (
            O => \N__19474\,
            I => clkdiv_cry_5
        );

    \I__1771\ : InMux
    port map (
            O => \N__19471\,
            I => clkdiv_cry_6
        );

    \I__1770\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19465\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__19465\,
            I => \clkdivZ0Z_8\
        );

    \I__1768\ : InMux
    port map (
            O => \N__19462\,
            I => \bfn_1_16_0_\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19456\,
            I => \clkdivZ0Z_9\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19453\,
            I => clkdiv_cry_8
        );

    \I__1764\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19447\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__19447\,
            I => \clkdivZ0Z_10\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19444\,
            I => clkdiv_cry_9
        );

    \I__1761\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__19438\,
            I => \clkdivZ0Z_11\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19435\,
            I => clkdiv_cry_10
        );

    \I__1758\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19429\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19429\,
            I => \clkdivZ0Z_12\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19426\,
            I => clkdiv_cry_11
        );

    \I__1755\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__19420\,
            I => \clkdivZ0Z_13\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19417\,
            I => clkdiv_cry_12
        );

    \I__1752\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__19411\,
            I => \TXbuffer_RNO_1Z0Z_3\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19408\,
            I => \bfn_1_15_0_\
        );

    \I__1749\ : InMux
    port map (
            O => \N__19405\,
            I => clkdiv_cry_0
        );

    \I__1748\ : InMux
    port map (
            O => \N__19402\,
            I => clkdiv_cry_1
        );

    \I__1747\ : InMux
    port map (
            O => \N__19399\,
            I => clkdiv_cry_2
        );

    \I__1746\ : InMux
    port map (
            O => \N__19396\,
            I => clkdiv_cry_3
        );

    \I__1745\ : InMux
    port map (
            O => \N__19393\,
            I => clkdiv_cry_4
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__19390\,
            I => \TXbuffer_RNO_5Z0Z_4_cascade_\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__19387\,
            I => \TXbuffer_18_15_ns_1_4_cascade_\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19381\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19381\,
            I => \TXbuffer_RNO_1Z0Z_0\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__19378\,
            I => \TXbuffer_18_15_ns_1_0_cascade_\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__19375\,
            I => \TXbuffer_18_10_ns_1_3_cascade_\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__19372\,
            I => \TXbuffer_RNO_0Z0Z_3_cascade_\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__19369\,
            I => \TXbuffer_18_10_ns_1_4_cascade_\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19363\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19363\,
            I => \N__19360\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__19360\,
            I => \TXbuffer_RNO_0Z0Z_4\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__19357\,
            I => \ALU.a6_b_9_cascade_\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__19354\,
            I => \ALU.madd_490_10_cascade_\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__19351\,
            I => \ALU.madd_490_7_cascade_\
        );

    \I__1730\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19345\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__19345\,
            I => \ALU.madd_490_11\
        );

    \I__1728\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19339\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__19339\,
            I => \ALU.a2_b_13\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__19336\,
            I => \TXbuffer_18_13_ns_1_0_cascade_\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__19333\,
            I => \TXbuffer_18_6_ns_1_2_cascade_\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__19330\,
            I => \TXbuffer_RNO_6Z0Z_2_cascade_\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__19321\,
            I => \ALU.madd_417\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__19318\,
            I => \ALU.madd_490_1_0_cascade_\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__19315\,
            I => \N__19312\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19309\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__19306\,
            I => \N__19303\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__19303\,
            I => \ALU.madd_378_0\
        );

    \I__1714\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19297\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__19297\,
            I => \N__19294\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__19294\,
            I => \ALU.madd_388\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__19291\,
            I => \ALU.madd_402_cascade_\
        );

    \I__1710\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19285\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__19285\,
            I => \N__19280\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19275\
        );

    \I__1707\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19275\
        );

    \I__1706\ : Odrv12
    port map (
            O => \N__19280\,
            I => \ALU.madd_330\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__19275\,
            I => \ALU.madd_330\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19267\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__19267\,
            I => \ALU.madd_490_21\
        );

    \I__1702\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19258\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__19258\,
            I => \ALU.madd_397\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \ALU.madd_388_cascade_\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__19252\,
            I => \ALU.madd_403_cascade_\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__19249\,
            I => \N__19246\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19243\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__19243\,
            I => \ALU.a1_b_13\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__19240\,
            I => \ALU.madd_403_0_cascade_\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__19237\,
            I => \ALU.a_6_ns_1_2_cascade_\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__19234\,
            I => \TXbuffer_18_13_ns_1_2_cascade_\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__19231\,
            I => \ALU.madd_311_cascade_\
        );

    \I__1690\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__19225\,
            I => \ALU.madd_268\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__19222\,
            I => \ALU.madd_268_cascade_\
        );

    \I__1687\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19216\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__19216\,
            I => \ALU.madd_311\
        );

    \I__1685\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19207\
        );

    \I__1684\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19207\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__19207\,
            I => \ALU.madd_316\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19198\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19198\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__19198\,
            I => \ALU.a8_b_5\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__19195\,
            I => \ALU.a1_b_13_cascade_\
        );

    \I__1678\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__19189\,
            I => \ALU.madd_171_0_tz\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__19186\,
            I => \ALU.madd_171_cascade_\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__19183\,
            I => \ALU.madd_315_0_tz_cascade_\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19176\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19173\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19176\,
            I => \ALU.madd_214\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__19173\,
            I => \ALU.madd_214\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__19168\,
            I => \ALU.madd_234_cascade_\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__19165\,
            I => \ALU.a7_b_8_cascade_\
        );

    \I__1668\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__19159\,
            I => \ALU.madd_490_3\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__19156\,
            I => \ALU.madd_171_0_tz_cascade_\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19150\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__19150\,
            I => \ALU.madd_97\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__19147\,
            I => \ALU.madd_171_x_cascade_\
        );

    \I__1662\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__19141\,
            I => \ALU.g0_2\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__19138\,
            I => \ALU.a5_b_4_cascade_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19126\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19126\
        );

    \I__1657\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19126\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__19126\,
            I => \ALU.madd_139\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__19123\,
            I => \ALU.a2_b_8_cascade_\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__19120\,
            I => \ALU.madd_181_cascade_\
        );

    \I__1653\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19110\
        );

    \I__1652\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19110\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19107\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__19110\,
            I => \ALU.a3_b_8\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19107\,
            I => \ALU.a3_b_8\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__19102\,
            I => \ALU.a3_b_8_cascade_\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \N__19095\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19092\
        );

    \I__1645\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19089\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__19092\,
            I => \ALU.madd_181\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__19089\,
            I => \ALU.madd_181\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__19084\,
            I => \ALU.N_675_0_0_cascade_\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__19081\,
            I => \ALU.N_703_0_0_0_cascade_\
        );

    \I__1640\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19075\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__19072\,
            I => \ALU.N_681_0_0_0\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \ALU.g0_0_2_cascade_\
        );

    \I__1636\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19063\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__19063\,
            I => \ALU.N_699_0\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__19060\,
            I => \ALU.madd_167_cascade_\
        );

    \I__1633\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__1632\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19051\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__19051\,
            I => \ALU.madd_167\
        );

    \INVFTDI.baudAcc_0C\ : INV
    port map (
            O => \INVFTDI.baudAcc_0C_net\,
            I => \N__56247\
        );

    \INVFTDI.TXstate_3C\ : INV
    port map (
            O => \INVFTDI.TXstate_3C_net\,
            I => \N__56244\
        );

    \INVFTDI.TXstate_0C\ : INV
    port map (
            O => \INVFTDI.TXstate_0C_net\,
            I => \N__56238\
        );

    \INVFTDI.TXshift_0C\ : INV
    port map (
            O => \INVFTDI.TXshift_0C_net\,
            I => \N__56243\
        );

    \INVFTDI.TXstate_2C\ : INV
    port map (
            O => \INVFTDI.TXstate_2C_net\,
            I => \N__56237\
        );

    \INVFTDI.TXstate_1C\ : INV
    port map (
            O => \INVFTDI.TXstate_1C_net\,
            I => \N__56235\
        );

    \INVFTDI.TXshift_4C\ : INV
    port map (
            O => \INVFTDI.TXshift_4C_net\,
            I => \N__56239\
        );

    \INVFTDI.TXshift_1C\ : INV
    port map (
            O => \INVFTDI.TXshift_1C_net\,
            I => \N__56236\
        );

    \INVFTDI.TXshift_7C\ : INV
    port map (
            O => \INVFTDI.TXshift_7C_net\,
            I => \N__56233\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_7_s1\,
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_7_s0\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_11_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_1_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_6_s1\,
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_13_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_3_0_\
        );

    \IN_MUX_bfv_13_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_6_s0\,
            carryinitout => \bfn_13_4_0_\
        );

    \IN_MUX_bfv_13_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_5_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_4\,
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_16_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_5_0_\
        );

    \IN_MUX_bfv_16_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_3\,
            carryinitout => \bfn_16_6_0_\
        );

    \IN_MUX_bfv_14_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_1_0_\
        );

    \IN_MUX_bfv_14_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_2\,
            carryinitout => \bfn_14_2_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_1\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_18_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_6_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_9_s1\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_9_s0\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_8_s1\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_8_s0\,
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_5_s1\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_5_s0\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_15_s1\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_15_s0\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_14_s1\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_14_s0\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_13_s1\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_6_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_13_s0\,
            carryinitout => \bfn_6_16_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_12_s1\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_12_s0\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_11_s1\,
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_11_s0\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_10_s1\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_prm_2_10_s0\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_12_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_2_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_s1_0\,
            carryinitout => \bfn_12_3_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.r0_12_s0_0\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.madd_cry_7\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_7,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_15,
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.un9_addsub_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.un2_addsub_cry_7\,
            carryinitout => \bfn_10_10_0_\
        );

    \clkdiv_RNIQAHO1_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26956\,
            GLOBALBUFFEROUTPUT => params5_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \ALU.mult_madd_159_N_2L1_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46375\,
            in2 => \_gnd_net_\,
            in3 => \N__48612\,
            lcout => \ALU.madd_159_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_134_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22123\,
            in1 => \N__38018\,
            in2 => \N__23050\,
            in3 => \N__52275\,
            lcout => \ALU.madd_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_17_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__47424\,
            in1 => \N__49003\,
            in2 => \N__20524\,
            in3 => \N__22096\,
            lcout => \ALU.N_681_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_20_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22122\,
            in1 => \N__38019\,
            in2 => \N__23049\,
            in3 => \N__52276\,
            lcout => OPEN,
            ltout => \ALU.N_675_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_15_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__19897\,
            in1 => \N__19639\,
            in2 => \N__19084\,
            in3 => \N__21535\,
            lcout => OPEN,
            ltout => \ALU.N_703_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_1_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20641\,
            in1 => \N__19066\,
            in2 => \N__19081\,
            in3 => \N__19144\,
            lcout => OPEN,
            ltout => \ALU.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_14_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111000"
        )
    port map (
            in0 => \N__19819\,
            in1 => \N__19078\,
            in2 => \N__19069\,
            in3 => \N__19668\,
            lcout => \ALU.N_724_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_18_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__19057\,
            in1 => \N__19135\,
            in2 => \_gnd_net_\,
            in3 => \N__19756\,
            lcout => \ALU.N_699_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_167_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22189\,
            in1 => \N__52253\,
            in2 => \_gnd_net_\,
            in3 => \N__46796\,
            lcout => \ALU.madd_167\,
            ltout => \ALU.madd_167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_187_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19133\,
            in2 => \N__19060\,
            in3 => \N__19754\,
            lcout => \ALU.madd_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_1_0_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19116\,
            in1 => \N__19785\,
            in2 => \_gnd_net_\,
            in3 => \N__21741\,
            lcout => \ALU.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_191_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__19056\,
            in1 => \N__19134\,
            in2 => \_gnd_net_\,
            in3 => \N__19755\,
            lcout => \ALU.madd_191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_2_0_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19117\,
            in1 => \N__19786\,
            in2 => \N__19099\,
            in3 => \N__21742\,
            lcout => \ALU.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_4_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__29101\,
            in1 => \N__29013\,
            in2 => \N__29245\,
            in3 => \N__40530\,
            lcout => OPEN,
            ltout => \ALU.a5_b_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_139_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__43393\,
            in1 => \N__21874\,
            in2 => \N__19138\,
            in3 => \N__44349\,
            lcout => \ALU.madd_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_10_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__42827\,
            in1 => \N__43637\,
            in2 => \N__19855\,
            in3 => \N__19833\,
            lcout => \ALU.N_695_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_7_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__44723\,
            in1 => \N__31922\,
            in2 => \N__36769\,
            in3 => \N__31834\,
            lcout => \ALU.a3_b_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_8_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32665\,
            in1 => \N__32590\,
            in2 => \N__29244\,
            in3 => \N__46334\,
            lcout => \ALU.a2_b_8\,
            ltout => \ALU.a2_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_181_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__43636\,
            in1 => \N__19850\,
            in2 => \N__19123\,
            in3 => \N__42826\,
            lcout => \ALU.madd_181\,
            ltout => \ALU.madd_181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_238_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011101000"
        )
    port map (
            in0 => \N__21734\,
            in1 => \N__19783\,
            in2 => \N__19120\,
            in3 => \N__19115\,
            lcout => \ALU.madd_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_8_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46335\,
            in1 => \N__31923\,
            in2 => \N__32262\,
            in3 => \N__31835\,
            lcout => \ALU.a3_b_8\,
            ltout => \ALU.a3_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_234_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21735\,
            in1 => \N__19784\,
            in2 => \N__19102\,
            in3 => \N__19098\,
            lcout => \ALU.madd_234\,
            ltout => \ALU.madd_234_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_248_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101000"
        )
    port map (
            in0 => \N__19697\,
            in1 => \N__19663\,
            in2 => \N__19168\,
            in3 => \N__19710\,
            lcout => \ALU.madd_308_0_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a7_b_8_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46433\,
            in1 => \N__23107\,
            in2 => \N__32278\,
            in3 => \N__30723\,
            lcout => OPEN,
            ltout => \ALU.a7_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_9_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19162\,
            in1 => \N__43631\,
            in2 => \N__19165\,
            in3 => \N__52199\,
            lcout => \ALU.madd_490_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_3_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__46795\,
            in1 => \N__44783\,
            in2 => \N__47071\,
            in3 => \N__46139\,
            lcout => \ALU.madd_490_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_1_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__43950\,
            in1 => \N__41570\,
            in2 => \N__45249\,
            in3 => \N__51810\,
            lcout => \ALU.madd_490_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_170_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46793\,
            in1 => \N__46135\,
            in2 => \N__52254\,
            in3 => \N__43949\,
            lcout => \ALU.madd_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_171_0_tz_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__43948\,
            in1 => \N__52198\,
            in2 => \N__46189\,
            in3 => \N__46794\,
            lcout => \ALU.madd_171_0_tz\,
            ltout => \ALU.madd_171_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_171_x_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__51809\,
            in1 => \_gnd_net_\,
            in2 => \N__19156\,
            in3 => \N__38017\,
            lcout => OPEN,
            ltout => \ALU.madd_171_x_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_229_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__19153\,
            in1 => \N__19179\,
            in2 => \N__19147\,
            in3 => \N__19920\,
            lcout => \ALU.madd_229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a8_b_5_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__45194\,
            in1 => \N__23410\,
            in2 => \N__36763\,
            in3 => \N__30622\,
            lcout => \ALU.a8_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_171_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__51811\,
            in1 => \N__19192\,
            in2 => \N__22066\,
            in3 => \N__37896\,
            lcout => OPEN,
            ltout => \ALU.madd_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_233_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__19180\,
            in1 => \_gnd_net_\,
            in2 => \N__19186\,
            in3 => \N__19921\,
            lcout => \ALU.madd_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_378_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__43376\,
            in1 => \N__46456\,
            in2 => \N__43666\,
            in3 => \N__46188\,
            lcout => \ALU.madd_378_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_315_0_tz_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__40987\,
            in1 => \N__43937\,
            in2 => \N__41364\,
            in3 => \N__46805\,
            lcout => OPEN,
            ltout => \ALU.madd_315_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_315_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41566\,
            in2 => \N__19183\,
            in3 => \N__37895\,
            lcout => \ALU.madd_315_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_214_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__45195\,
            in1 => \N__24415\,
            in2 => \_gnd_net_\,
            in3 => \N__43375\,
            lcout => \ALU.madd_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_314_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46806\,
            in1 => \N__41339\,
            in2 => \N__43954\,
            in3 => \N__40988\,
            lcout => \ALU.madd_181_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_297_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20885\,
            in1 => \N__21009\,
            in2 => \N__21043\,
            in3 => \N__22231\,
            lcout => \ALU.madd_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_311_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__46807\,
            in1 => \_gnd_net_\,
            in2 => \N__41365\,
            in3 => \N__24445\,
            lcout => \ALU.madd_311\,
            ltout => \ALU.madd_311_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_340_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19213\,
            in2 => \N__19231\,
            in3 => \N__19228\,
            lcout => \ALU.madd_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_268_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22207\,
            in1 => \N__23256\,
            in2 => \_gnd_net_\,
            in3 => \N__21210\,
            lcout => \ALU.madd_268\,
            ltout => \ALU.madd_268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_336_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19212\,
            in2 => \N__19222\,
            in3 => \N__19219\,
            lcout => \ALU.madd_336_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_316_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19203\,
            in1 => \N__51742\,
            in2 => \N__23196\,
            in3 => \N__44344\,
            lcout => \ALU.madd_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_298_0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101000"
        )
    port map (
            in0 => \N__20907\,
            in1 => \N__21010\,
            in2 => \N__20892\,
            in3 => \N__21079\,
            lcout => \ALU.madd_298_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_320_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__19204\,
            in1 => \N__51743\,
            in2 => \N__23197\,
            in3 => \N__44345\,
            lcout => \ALU.madd_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_330_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__20158\,
            in1 => \N__47352\,
            in2 => \N__20152\,
            in3 => \N__42843\,
            lcout => \ALU.madd_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a1_b_13_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__35374\,
            in1 => \N__31655\,
            in2 => \N__32202\,
            in3 => \N__31741\,
            lcout => \ALU.a1_b_13\,
            ltout => \ALU.a1_b_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_388_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__39863\,
            in1 => \N__22159\,
            in2 => \N__19195\,
            in3 => \N__48391\,
            lcout => \ALU.madd_388\,
            ltout => \ALU.madd_388_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_403_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__20286\,
            in1 => \N__19284\,
            in2 => \N__19255\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ALU.madd_403_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_417_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__27280\,
            in1 => \N__20407\,
            in2 => \N__19252\,
            in3 => \N__21672\,
            lcout => \ALU.madd_417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_392_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__48390\,
            in1 => \N__39862\,
            in2 => \N__19249\,
            in3 => \N__22158\,
            lcout => \ALU.madd_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_403_0_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22157\,
            in1 => \N__20068\,
            in2 => \_gnd_net_\,
            in3 => \N__20285\,
            lcout => OPEN,
            ltout => \ALU.madd_403_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_413_0_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20406\,
            in1 => \N__19283\,
            in2 => \N__19240\,
            in3 => \N__27279\,
            lcout => \ALU.madd_413_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIS0G71_2_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__23378\,
            in1 => \N__25012\,
            in2 => \N__23361\,
            in3 => \N__31096\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIBF8D2_2_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__28089\,
            in1 => \N__39167\,
            in2 => \N__19237\,
            in3 => \N__30926\,
            lcout => \ALU.r6_RNIBF8D2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_2_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40296\,
            lcout => r2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56279\,
            ce => \N__47712\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_2_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__30040\,
            in1 => \N__22390\,
            in2 => \N__30387\,
            in3 => \N__23357\,
            lcout => OPEN,
            ltout => \TXbuffer_18_13_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_2_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__22684\,
            in1 => \N__30041\,
            in2 => \N__19234\,
            in3 => \N__28090\,
            lcout => \TXbuffer_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_2_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__30042\,
            in1 => \N__22297\,
            in2 => \N__30388\,
            in3 => \N__23379\,
            lcout => OPEN,
            ltout => \TXbuffer_18_6_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_2_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__39168\,
            in1 => \N__30043\,
            in2 => \N__19333\,
            in3 => \N__22572\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_6Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_2_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__22603\,
            in1 => \N__29670\,
            in2 => \N__19330\,
            in3 => \N__49932\,
            lcout => \TXbuffer_18_15_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_1_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19264\,
            in1 => \N__19270\,
            in2 => \_gnd_net_\,
            in3 => \N__19957\,
            lcout => OPEN,
            ltout => \ALU.madd_490_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20107\,
            in1 => \N__19327\,
            in2 => \N__19318\,
            in3 => \N__20320\,
            lcout => \ALU.madd_340_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_402_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__20359\,
            in1 => \N__20425\,
            in2 => \N__19315\,
            in3 => \N__24511\,
            lcout => OPEN,
            ltout => \ALU.madd_402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_21_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__20290\,
            in1 => \N__19300\,
            in2 => \N__19291\,
            in3 => \N__19288\,
            lcout => \ALU.madd_490_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_397_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101000"
        )
    port map (
            in0 => \N__19978\,
            in1 => \N__21790\,
            in2 => \N__20020\,
            in3 => \N__19998\,
            lcout => \ALU.madd_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r3_2_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40300\,
            lcout => r3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56287\,
            ce => \N__47763\,
            sr => \_gnd_net_\
        );

    \ALU.r3_3_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50199\,
            lcout => r3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56287\,
            ce => \N__47763\,
            sr => \_gnd_net_\
        );

    \ALU.mult_a6_b_9_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__47425\,
            in1 => \N__26513\,
            in2 => \N__36767\,
            in3 => \N__26449\,
            lcout => OPEN,
            ltout => \ALU.a6_b_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_10_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__40113\,
            in1 => \N__31954\,
            in2 => \N__19357\,
            in3 => \N__38021\,
            lcout => OPEN,
            ltout => \ALU.madd_490_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_13_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19354\,
            in3 => \N__19348\,
            lcout => \ALU.madd_490_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_7_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__39925\,
            in1 => \N__49013\,
            in2 => \N__47139\,
            in3 => \N__48613\,
            lcout => OPEN,
            ltout => \ALU.madd_490_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_11_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__39837\,
            in1 => \N__19342\,
            in2 => \N__19351\,
            in3 => \N__49418\,
            lcout => \ALU.madd_490_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_13_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__35373\,
            in1 => \N__32655\,
            in2 => \N__36766\,
            in3 => \N__32578\,
            lcout => \ALU.a2_b_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29969\,
            in1 => \N__23547\,
            in2 => \N__30310\,
            in3 => \N__28838\,
            lcout => OPEN,
            ltout => \TXbuffer_18_13_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29971\,
            in1 => \N__27826\,
            in2 => \N__19336\,
            in3 => \N__23326\,
            lcout => \TXbuffer_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_4_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29970\,
            in1 => \N__25452\,
            in2 => \N__22588\,
            in3 => \N__34300\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_5Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_4_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__49937\,
            in1 => \N__29661\,
            in2 => \N__19390\,
            in3 => \N__25231\,
            lcout => OPEN,
            ltout => \TXbuffer_18_15_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_4_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__49939\,
            in1 => \N__20536\,
            in2 => \N__19387\,
            in3 => \N__19366\,
            lcout => \TXbufferZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56296\,
            ce => \N__56037\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_0_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__49936\,
            in1 => \N__21523\,
            in2 => \N__29674\,
            in3 => \N__27655\,
            lcout => OPEN,
            ltout => \TXbuffer_18_15_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__49938\,
            in1 => \N__19384\,
            in2 => \N__19378\,
            in3 => \N__27607\,
            lcout => \TXbufferZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56296\,
            ce => \N__56037\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_3_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__29887\,
            in1 => \N__33244\,
            in2 => \N__25212\,
            in3 => \N__30240\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_3_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__29885\,
            in1 => \N__33610\,
            in2 => \N__19375\,
            in3 => \N__26118\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_3_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__49902\,
            in1 => \N__19414\,
            in2 => \N__19372\,
            in3 => \N__24844\,
            lcout => \TXbufferZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56300\,
            ce => \N__56036\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_4_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29884\,
            in1 => \N__25171\,
            in2 => \N__30304\,
            in3 => \N__33478\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_4_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29886\,
            in1 => \N__26083\,
            in2 => \N__19369\,
            in3 => \N__33574\,
            lcout => \TXbuffer_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXstart_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27075\,
            in1 => \N__26976\,
            in2 => \N__27015\,
            in3 => \N__27051\,
            lcout => \TXstartZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI7AQC9_0_15_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40084\,
            in2 => \_gnd_net_\,
            in3 => \N__39973\,
            lcout => \ALU.r2_RNI7AQC9_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_3_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__29859\,
            in1 => \N__28060\,
            in2 => \N__22651\,
            in3 => \N__20503\,
            lcout => \TXbuffer_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_0_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26975\,
            in2 => \_gnd_net_\,
            in3 => \N__19408\,
            lcout => \clkdivZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => clkdiv_cry_0,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_1_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27074\,
            in2 => \_gnd_net_\,
            in3 => \N__19405\,
            lcout => \clkdivZ0Z_1\,
            ltout => OPEN,
            carryin => clkdiv_cry_0,
            carryout => clkdiv_cry_1,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_2_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27050\,
            in2 => \_gnd_net_\,
            in3 => \N__19402\,
            lcout => \clkdivZ0Z_2\,
            ltout => OPEN,
            carryin => clkdiv_cry_1,
            carryout => clkdiv_cry_2,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_3_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27008\,
            in2 => \_gnd_net_\,
            in3 => \N__19399\,
            lcout => \clkdivZ0Z_3\,
            ltout => OPEN,
            carryin => clkdiv_cry_2,
            carryout => clkdiv_cry_3,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_4_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49853\,
            in2 => \_gnd_net_\,
            in3 => \N__19396\,
            lcout => \clkdivZ0Z_4\,
            ltout => OPEN,
            carryin => clkdiv_cry_3,
            carryout => clkdiv_cry_4,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_5_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29622\,
            in2 => \_gnd_net_\,
            in3 => \N__19393\,
            lcout => \clkdivZ0Z_5\,
            ltout => OPEN,
            carryin => clkdiv_cry_4,
            carryout => clkdiv_cry_5,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_6_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29842\,
            in2 => \_gnd_net_\,
            in3 => \N__19474\,
            lcout => \clkdivZ0Z_6\,
            ltout => OPEN,
            carryin => clkdiv_cry_5,
            carryout => clkdiv_cry_6,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_7_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30209\,
            in2 => \_gnd_net_\,
            in3 => \N__19471\,
            lcout => \clkdivZ0Z_7\,
            ltout => OPEN,
            carryin => clkdiv_cry_6,
            carryout => clkdiv_cry_7,
            clk => \N__56303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_8_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19468\,
            in2 => \_gnd_net_\,
            in3 => \N__19462\,
            lcout => \clkdivZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => clkdiv_cry_8,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_9_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19459\,
            in2 => \_gnd_net_\,
            in3 => \N__19453\,
            lcout => \clkdivZ0Z_9\,
            ltout => OPEN,
            carryin => clkdiv_cry_8,
            carryout => clkdiv_cry_9,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_10_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19450\,
            in2 => \_gnd_net_\,
            in3 => \N__19444\,
            lcout => \clkdivZ0Z_10\,
            ltout => OPEN,
            carryin => clkdiv_cry_9,
            carryout => clkdiv_cry_10,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_11_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19441\,
            in2 => \_gnd_net_\,
            in3 => \N__19435\,
            lcout => \clkdivZ0Z_11\,
            ltout => OPEN,
            carryin => clkdiv_cry_10,
            carryout => clkdiv_cry_11,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_12_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19432\,
            in2 => \_gnd_net_\,
            in3 => \N__19426\,
            lcout => \clkdivZ0Z_12\,
            ltout => OPEN,
            carryin => clkdiv_cry_11,
            carryout => clkdiv_cry_12,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_13_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19423\,
            in2 => \_gnd_net_\,
            in3 => \N__19417\,
            lcout => \clkdivZ0Z_13\,
            ltout => OPEN,
            carryin => clkdiv_cry_12,
            carryout => clkdiv_cry_13,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_14_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19555\,
            in2 => \_gnd_net_\,
            in3 => \N__19549\,
            lcout => \clkdivZ0Z_14\,
            ltout => OPEN,
            carryin => clkdiv_cry_13,
            carryout => clkdiv_cry_14,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_15_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19546\,
            in2 => \_gnd_net_\,
            in3 => \N__19540\,
            lcout => \clkdivZ0Z_15\,
            ltout => OPEN,
            carryin => clkdiv_cry_14,
            carryout => clkdiv_cry_15,
            clk => \N__56304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_16_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19537\,
            in2 => \_gnd_net_\,
            in3 => \N__19531\,
            lcout => \clkdivZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => clkdiv_cry_16,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_17_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19528\,
            in2 => \_gnd_net_\,
            in3 => \N__19522\,
            lcout => \clkdivZ0Z_17\,
            ltout => OPEN,
            carryin => clkdiv_cry_16,
            carryout => clkdiv_cry_17,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_18_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19519\,
            in2 => \_gnd_net_\,
            in3 => \N__19513\,
            lcout => \clkdivZ0Z_18\,
            ltout => OPEN,
            carryin => clkdiv_cry_17,
            carryout => clkdiv_cry_18,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_19_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19510\,
            in2 => \_gnd_net_\,
            in3 => \N__19504\,
            lcout => \clkdivZ0Z_19\,
            ltout => OPEN,
            carryin => clkdiv_cry_18,
            carryout => clkdiv_cry_19,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_20_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19501\,
            in2 => \_gnd_net_\,
            in3 => \N__19495\,
            lcout => \clkdivZ0Z_20\,
            ltout => OPEN,
            carryin => clkdiv_cry_19,
            carryout => clkdiv_cry_20,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_21_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19492\,
            in2 => \_gnd_net_\,
            in3 => \N__19486\,
            lcout => \clkdivZ0Z_21\,
            ltout => OPEN,
            carryin => clkdiv_cry_20,
            carryout => clkdiv_cry_21,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_22_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19483\,
            in2 => \_gnd_net_\,
            in3 => \N__19477\,
            lcout => \clkdivZ0Z_22\,
            ltout => OPEN,
            carryin => clkdiv_cry_21,
            carryout => clkdiv_cry_22,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_23_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19593\,
            in2 => \_gnd_net_\,
            in3 => \N__19603\,
            lcout => \GPIO3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_154_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__22841\,
            in1 => \N__21871\,
            in2 => \N__31575\,
            in3 => \N__21549\,
            lcout => \ALU.madd_154\,
            ltout => \ALU.madd_154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_0_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__19885\,
            in1 => \N__23128\,
            in2 => \N__19582\,
            in3 => \N__19642\,
            lcout => OPEN,
            ltout => \ALU.N_703_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__19669\,
            in1 => \N__19711\,
            in2 => \N__19579\,
            in3 => \N__19726\,
            lcout => OPEN,
            ltout => \ALU.g0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_10_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19572\,
            in1 => \N__26319\,
            in2 => \N__19576\,
            in3 => \N__26304\,
            lcout => \ALU.madd_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_150_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22842\,
            in1 => \N__21872\,
            in2 => \N__31576\,
            in3 => \N__21550\,
            lcout => \ALU.madd_150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_206_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__20689\,
            in1 => \N__19767\,
            in2 => \N__20584\,
            in3 => \N__19720\,
            lcout => \ALU.madd_206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_202_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19719\,
            in1 => \N__20580\,
            in2 => \N__19768\,
            in3 => \N__20688\,
            lcout => \ALU.madd_334\,
            ltout => \ALU.madd_334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_13_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010000000"
        )
    port map (
            in0 => \N__19573\,
            in1 => \N__20602\,
            in2 => \N__19564\,
            in3 => \N__19561\,
            lcout => \ALU.g0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_192_0_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__19815\,
            in1 => \_gnd_net_\,
            in2 => \N__47269\,
            in3 => \N__24394\,
            lcout => \ALU.madd_192_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_144_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__21883\,
            in1 => \N__22888\,
            in2 => \N__43649\,
            in3 => \N__49361\,
            lcout => \ALU.madd_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_3_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19744\,
            in1 => \N__19698\,
            in2 => \N__19738\,
            in3 => \N__20639\,
            lcout => \ALU.g0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_197_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19640\,
            in1 => \N__19620\,
            in2 => \N__19883\,
            in3 => \N__19611\,
            lcout => \ALU.madd_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_195_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20686\,
            lcout => \ALU.madd_112\,
            ltout => \ALU.madd_112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_244_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__19699\,
            in1 => \N__19681\,
            in2 => \N__19672\,
            in3 => \N__19664\,
            lcout => \ALU.madd_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_196_0_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000101000"
        )
    port map (
            in0 => \N__19814\,
            in1 => \N__24393\,
            in2 => \N__47268\,
            in3 => \N__20687\,
            lcout => \ALU.madd_196_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_201_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011101000"
        )
    port map (
            in0 => \N__19641\,
            in1 => \N__19621\,
            in2 => \N__19884\,
            in3 => \N__19612\,
            lcout => \ALU.madd_201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_239_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__20748\,
            in1 => \N__19797\,
            in2 => \N__23164\,
            in3 => \N__20730\,
            lcout => \ALU.madd_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g2_0_1_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__51988\,
            in1 => \N__48928\,
            in2 => \N__47457\,
            in3 => \N__48570\,
            lcout => \ALU.g2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_182_0_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__48569\,
            in1 => \N__47423\,
            in2 => \N__48988\,
            in3 => \N__51987\,
            lcout => \ALU.madd_182_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_0_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__38020\,
            in1 => \N__48571\,
            in2 => \N__46823\,
            in3 => \N__48932\,
            lcout => \ALU.mult_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_177_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__42753\,
            in1 => \N__19854\,
            in2 => \N__19837\,
            in3 => \N__43635\,
            lcout => \ALU.madd_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_243_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101000"
        )
    port map (
            in0 => \N__19798\,
            in1 => \N__23163\,
            in2 => \N__20734\,
            in3 => \N__20749\,
            lcout => \ALU.madd_243\,
            ltout => \ALU.madd_243_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_299_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__21183\,
            in1 => \N__20770\,
            in2 => \N__19789\,
            in3 => \N__22871\,
            lcout => \ALU.madd_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_219_0_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__44766\,
            in1 => \N__45461\,
            in2 => \N__43664\,
            in3 => \N__42752\,
            lcout => \ALU.madd_219_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_304_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20865\,
            in1 => \N__19944\,
            in2 => \_gnd_net_\,
            in3 => \N__19929\,
            lcout => \ALU.madd_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_303_0_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__22873\,
            in1 => \N__20769\,
            in2 => \N__21187\,
            in3 => \N__19909\,
            lcout => \ALU.madd_303_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_293_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__20794\,
            in1 => \_gnd_net_\,
            in2 => \N__20788\,
            in3 => \N__20970\,
            lcout => \ALU.madd_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_393_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__20013\,
            in1 => \N__21786\,
            in2 => \N__20002\,
            in3 => \N__19977\,
            lcout => \ALU.madd_393\,
            ltout => \ALU.madd_393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_412_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20047\,
            in2 => \N__19960\,
            in3 => \N__20923\,
            lcout => \ALU.madd_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_308_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__19945\,
            in1 => \_gnd_net_\,
            in2 => \N__19933\,
            in3 => \N__20866\,
            lcout => \ALU.madd_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_209_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__51808\,
            in1 => \N__23011\,
            in2 => \_gnd_net_\,
            in3 => \N__46789\,
            lcout => \ALU.madd_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_302_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20768\,
            in2 => \_gnd_net_\,
            in3 => \N__19908\,
            lcout => \ALU.madd_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_365_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101000"
        )
    port map (
            in0 => \N__20212\,
            in1 => \N__20098\,
            in2 => \N__20092\,
            in3 => \N__20077\,
            lcout => \ALU.madd_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_13_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35387\,
            in2 => \_gnd_net_\,
            in3 => \N__49004\,
            lcout => \ALU.a0_b_13\,
            ltout => \ALU.a0_b_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_331_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__48608\,
            in1 => \N__39813\,
            in2 => \N__19900\,
            in3 => \N__21261\,
            lcout => \ALU.madd_331_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_356_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__20194\,
            in1 => \N__20200\,
            in2 => \N__20820\,
            in3 => \N__20178\,
            lcout => \ALU.madd_356\,
            ltout => \ALU.madd_356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_361_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__20088\,
            in1 => \N__20211\,
            in2 => \N__20080\,
            in3 => \N__20076\,
            lcout => \ALU.madd_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_388_0_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__48365\,
            in1 => \N__35388\,
            in2 => \N__39849\,
            in3 => \N__48609\,
            lcout => \ALU.madd_388_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_1_c_RNO_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41823\,
            lcout => \ALU.r0_12_prm_3_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_RNO_4_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__48366\,
            in1 => \N__53516\,
            in2 => \N__54478\,
            in3 => \N__48610\,
            lcout => \ALU.rshift_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_427_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111001001000"
        )
    port map (
            in0 => \N__20248\,
            in1 => \N__20026\,
            in2 => \N__21673\,
            in3 => \N__20167\,
            lcout => \ALU.madd_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_408_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20056\,
            in1 => \N__20922\,
            in2 => \_gnd_net_\,
            in3 => \N__20043\,
            lcout => \ALU.madd_408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_355_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__20220\,
            in1 => \N__20232\,
            in2 => \_gnd_net_\,
            in3 => \N__21243\,
            lcout => \ALU.madd_355\,
            ltout => \ALU.madd_355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_418_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__20982\,
            in1 => \N__20121\,
            in2 => \N__20029\,
            in3 => \N__20134\,
            lcout => \ALU.madd_418\,
            ltout => \ALU.madd_418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_423_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20247\,
            in1 => \N__21668\,
            in2 => \N__20239\,
            in3 => \N__20166\,
            lcout => \ALU.madd_338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_351_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__21244\,
            in1 => \_gnd_net_\,
            in2 => \N__20236\,
            in3 => \N__20221\,
            lcout => \ALU.madd_351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_346_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20143\,
            in1 => \N__21059\,
            in2 => \_gnd_net_\,
            in3 => \N__21100\,
            lcout => \ALU.madd_346\,
            ltout => \ALU.madd_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_360_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101000"
        )
    port map (
            in0 => \N__20821\,
            in1 => \N__20193\,
            in2 => \N__20182\,
            in3 => \N__20179\,
            lcout => \ALU.madd_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_329_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49364\,
            in1 => \N__51919\,
            in2 => \N__35540\,
            in3 => \N__48364\,
            lcout => \ALU.madd_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_330_0_tz_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__48363\,
            in1 => \N__35500\,
            in2 => \N__51958\,
            in3 => \N__49365\,
            lcout => \ALU.madd_330_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_326_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__35496\,
            in1 => \_gnd_net_\,
            in2 => \N__20269\,
            in3 => \N__48362\,
            lcout => \ALU.madd_326\,
            ltout => \ALU.madd_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_350_0_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21130\,
            in2 => \N__20137\,
            in3 => \N__21064\,
            lcout => \ALU.madd_350_0\,
            ltout => \ALU.madd_350_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_422_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101000"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__20122\,
            in2 => \N__20110\,
            in3 => \N__20983\,
            lcout => \ALU.madd_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a7_b_7_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__44776\,
            in1 => \N__23102\,
            in2 => \N__32201\,
            in3 => \N__30722\,
            lcout => \ALU.a7_b_7\,
            ltout => \ALU.a7_b_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_383_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__49363\,
            in1 => \N__35539\,
            in2 => \N__20293\,
            in3 => \N__20373\,
            lcout => \ALU.madd_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a4_b_10_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__51918\,
            in1 => \N__32464\,
            in2 => \N__32200\,
            in3 => \N__32372\,
            lcout => \ALU.a4_b_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIU2J74_9_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24630\,
            in1 => \N__21306\,
            in2 => \_gnd_net_\,
            in3 => \N__21288\,
            lcout => \ALU.b_9\,
            ltout => \ALU.b_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_326_0_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__42842\,
            in1 => \N__51917\,
            in2 => \N__20272\,
            in3 => \N__49362\,
            lcout => \ALU.madd_326_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_11_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__35501\,
            in1 => \N__31921\,
            in2 => \N__31833\,
            in3 => \N__32199\,
            lcout => \ALU.a3_b_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_9_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__29003\,
            in1 => \N__29077\,
            in2 => \N__32237\,
            in3 => \N__47342\,
            lcout => \ALU.a5_b_9\,
            ltout => \ALU.a5_b_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_382_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__43651\,
            in2 => \N__20260\,
            in3 => \N__46173\,
            lcout => \ALU.madd_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a6_b_8_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__26504\,
            in1 => \N__26435\,
            in2 => \N__32238\,
            in3 => \N__46432\,
            lcout => \ALU.a6_b_8\,
            ltout => \ALU.a6_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_378_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__20421\,
            in1 => \N__43650\,
            in2 => \N__20410\,
            in3 => \N__46172\,
            lcout => \ALU.madd_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNILIOQ3_3_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__32883\,
            in1 => \N__24336\,
            in2 => \_gnd_net_\,
            in3 => \N__33036\,
            lcout => \ALU.b_i_3\,
            ltout => \ALU.b_i_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNINFAJC_3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20395\,
            in3 => \N__24307\,
            lcout => \ALU.r4_RNINFAJCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_16_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001101100"
        )
    port map (
            in0 => \N__20392\,
            in1 => \N__20383\,
            in2 => \N__48061\,
            in3 => \N__20377\,
            lcout => \ALU.madd_490_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a11_b_3_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__24337\,
            in1 => \N__33037\,
            in2 => \N__32895\,
            in3 => \N__40892\,
            lcout => \ALU.a11_b_3\,
            ltout => \ALU.a11_b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_373_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__36486\,
            in1 => \N__45222\,
            in2 => \N__20362\,
            in3 => \N__52299\,
            lcout => \ALU.madd_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_15_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001101100"
        )
    port map (
            in0 => \N__27306\,
            in1 => \N__24484\,
            in2 => \N__20353\,
            in3 => \N__36487\,
            lcout => OPEN,
            ltout => \ALU.madd_490_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_19_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20344\,
            in1 => \N__20329\,
            in2 => \N__20323\,
            in3 => \N__20440\,
            lcout => \ALU.madd_490_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_14_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__20314\,
            in1 => \N__20959\,
            in2 => \N__20302\,
            in3 => \N__20944\,
            lcout => \ALU.madd_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIE0AK8_1_11_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__40957\,
            in1 => \_gnd_net_\,
            in2 => \N__35592\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r5_RNIE0AK8_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIAFSR_15_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30480\,
            in1 => \N__30117\,
            in2 => \_gnd_net_\,
            in3 => \N__29507\,
            lcout => \ALU.r1_RNIAFSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__40521\,
            in1 => \N__44361\,
            in2 => \N__41362\,
            in3 => \N__40956\,
            lcout => OPEN,
            ltout => \ALU.madd_490_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_14_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20479\,
            in1 => \N__20464\,
            in2 => \N__20449\,
            in3 => \N__20446\,
            lcout => \ALU.madd_490_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNISP2L9_2_12_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39826\,
            in1 => \_gnd_net_\,
            in2 => \N__41363\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r5_RNISP2L9_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIFR6T_15_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25079\,
            in1 => \N__22511\,
            in2 => \_gnd_net_\,
            in3 => \N__22431\,
            lcout => OPEN,
            ltout => \ALU.r2_RNIFR6TZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI418R4_15_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__32892\,
            in1 => \N__21406\,
            in2 => \N__20431\,
            in3 => \N__20485\,
            lcout => \ALU.b_15\,
            ltout => \ALU.b_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_15_s1_c_RNO_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101010101"
        )
    port map (
            in0 => \N__53254\,
            in1 => \_gnd_net_\,
            in2 => \N__20428\,
            in3 => \N__40114\,
            lcout => \ALU.r0_12_prm_7_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_7_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__22512\,
            in1 => \N__29975\,
            in2 => \N__22486\,
            in3 => \N__30281\,
            lcout => \TXbuffer_18_13_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_3_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29976\,
            in1 => \N__22362\,
            in2 => \N__30336\,
            in3 => \N__23658\,
            lcout => \TXbuffer_18_13_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIJBVT_15_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30447\,
            in1 => \N__25078\,
            in2 => \_gnd_net_\,
            in3 => \N__29721\,
            lcout => OPEN,
            ltout => \ALU.r5_RNIJBVTZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIJING2_15_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__24641\,
            in1 => \N__20494\,
            in2 => \N__20488\,
            in3 => \N__21963\,
            lcout => \ALU.b_7_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_11_s1_c_RNO_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__35568\,
            in1 => \N__53238\,
            in2 => \N__54780\,
            in3 => \N__40960\,
            lcout => \ALU.r0_12_prm_5_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIE0AK8_2_11_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__40961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35566\,
            lcout => \ALU.r5_RNIE0AK8_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_9_s0_c_RNO_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55968\,
            in2 => \_gnd_net_\,
            in3 => \N__42448\,
            lcout => \ALU.r0_12_prm_2_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIUF9K8_2_10_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51983\,
            in2 => \_gnd_net_\,
            in3 => \N__51836\,
            lcout => \ALU.r5_RNIUF9K8_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_11_s1_c_RNO_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__35567\,
            in1 => \N__53237\,
            in2 => \_gnd_net_\,
            in3 => \N__40959\,
            lcout => \ALU.r0_12_prm_7_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIAG9A9_15_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53680\,
            in1 => \N__40054\,
            in2 => \_gnd_net_\,
            in3 => \N__47046\,
            lcout => \ALU.r5_RNIAG9A9Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIE0AK8_0_11_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40958\,
            lcout => \ALU.r5_RNIE0AK8_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_15_s1_c_RNO_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__40086\,
            in1 => \N__53256\,
            in2 => \N__54778\,
            in3 => \N__53685\,
            lcout => \ALU.r0_12_prm_4_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_15_s1_c_RNO_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__39957\,
            in1 => \N__53255\,
            in2 => \N__53899\,
            in3 => \N__40085\,
            lcout => \ALU.r0_12_prm_6_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI39IH4_15_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25492\,
            in1 => \N__36764\,
            in2 => \_gnd_net_\,
            in3 => \N__21412\,
            lcout => \ALU.a_15\,
            ltout => \ALU.a_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNINNEH9_15_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__53681\,
            in1 => \N__47033\,
            in2 => \N__20512\,
            in3 => \N__54585\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIVF7TI_13_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__54586\,
            in1 => \N__41520\,
            in2 => \N__20509\,
            in3 => \N__41317\,
            lcout => \ALU.r5_RNIVF7TIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_11_s1_c_RNO_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__53686\,
            in1 => \N__55969\,
            in2 => \_gnd_net_\,
            in3 => \N__35768\,
            lcout => \ALU.r0_12_prm_1_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_13_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26281\,
            lcout => r2_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56301\,
            ce => \N__47707\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINFOB1_13_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__25066\,
            in1 => \N__24106\,
            in2 => \N__22000\,
            in3 => \N__23906\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIC9GA2_13_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__23988\,
            in1 => \N__24078\,
            in2 => \N__20506\,
            in3 => \N__21999\,
            lcout => OPEN,
            ltout => \ALU.r6_RNIC9GA2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIR9125_13_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__21421\,
            in1 => \_gnd_net_\,
            in2 => \N__20545\,
            in3 => \N__32896\,
            lcout => \ALU.b_13\,
            ltout => \ALU.b_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNID2JJ9_2_13_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__41544\,
            in1 => \_gnd_net_\,
            in2 => \N__20542\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r5_RNID2JJ9_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNID2JJ9_0_13_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35347\,
            in2 => \_gnd_net_\,
            in3 => \N__41542\,
            lcout => \ALU.r5_RNID2JJ9_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNID2JJ9_1_13_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35348\,
            in2 => \_gnd_net_\,
            in3 => \N__41543\,
            lcout => \ALU.r5_RNID2JJ9_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_4_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__29934\,
            in1 => \N__23872\,
            in2 => \N__24958\,
            in3 => \N__30208\,
            lcout => OPEN,
            ltout => \TXbuffer_18_13_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_4_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29844\,
            in1 => \N__23622\,
            in2 => \N__20539\,
            in3 => \N__28027\,
            lcout => \TXbuffer_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_6_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29843\,
            in1 => \N__25861\,
            in2 => \N__30268\,
            in3 => \N__23745\,
            lcout => \TXbuffer_18_6_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_5_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29903\,
            in1 => \N__26212\,
            in2 => \N__30360\,
            in3 => \N__22333\,
            lcout => \TXbuffer_18_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_4_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__46204\,
            in1 => \N__20704\,
            in2 => \N__20722\,
            in3 => \N__37964\,
            lcout => \ALU.N_661_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_155_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__21607\,
            in1 => \N__48576\,
            in2 => \N__46431\,
            in3 => \N__20665\,
            lcout => \ALU.madd_155\,
            ltout => \ALU.madd_155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_160_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20568\,
            in2 => \N__20611\,
            in3 => \N__22814\,
            lcout => \ALU.madd_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_109_0_tz_LC_3_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__44750\,
            in1 => \N__46383\,
            in2 => \N__48987\,
            in3 => \N__48575\,
            lcout => OPEN,
            ltout => \ALU.madd_109_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_109_LC_3_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__43570\,
            in1 => \N__48351\,
            in2 => \N__20608\,
            in3 => \N__21625\,
            lcout => \ALU.madd_109\,
            ltout => \ALU.madd_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_5_LC_3_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000101000"
        )
    port map (
            in0 => \N__22816\,
            in1 => \N__21850\,
            in2 => \N__20605\,
            in3 => \N__20557\,
            lcout => \ALU.N_687_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_159_LC_3_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001011101011"
        )
    port map (
            in0 => \N__20664\,
            in1 => \N__20596\,
            in2 => \N__21619\,
            in3 => \N__21631\,
            lcout => \ALU.madd_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_164_LC_3_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__22815\,
            in1 => \_gnd_net_\,
            in2 => \N__20572\,
            in3 => \N__20556\,
            lcout => \ALU.madd_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a4_b_5_LC_3_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32470\,
            in1 => \N__32376\,
            in2 => \N__29226\,
            in3 => \N__45180\,
            lcout => \ALU.a4_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a7_b_1_LC_3_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44549\,
            in2 => \_gnd_net_\,
            in3 => \N__46750\,
            lcout => \ALU.a7_b_1\,
            ltout => \ALU.a7_b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_95_LC_3_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__46153\,
            in1 => \N__20718\,
            in2 => \N__20548\,
            in3 => \N__37966\,
            lcout => \ALU.madd_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a6_b_2_LC_3_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__26512\,
            in1 => \N__26448\,
            in2 => \N__29227\,
            in3 => \N__43928\,
            lcout => \ALU.a6_b_2\,
            ltout => \ALU.a6_b_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_99_LC_3_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__46152\,
            in1 => \N__37965\,
            in2 => \N__20707\,
            in3 => \N__20703\,
            lcout => \ALU.madd_99\,
            ltout => \ALU.madd_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_149_LC_3_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__48926\,
            in1 => \N__47413\,
            in2 => \N__20692\,
            in3 => \N__22091\,
            lcout => \ALU.madd_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_145_LC_3_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__22092\,
            in1 => \N__20671\,
            in2 => \N__47455\,
            in3 => \N__48927\,
            lcout => \ALU.madd_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_253_LC_3_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__20656\,
            in1 => \_gnd_net_\,
            in2 => \N__20650\,
            in3 => \N__20640\,
            lcout => \ALU.madd_253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_9_LC_3_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__47436\,
            in1 => \N__31924\,
            in2 => \N__31840\,
            in3 => \N__36759\,
            lcout => \ALU.a3_b_9\,
            ltout => \ALU.a3_b_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_274_LC_3_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__21093\,
            in1 => \N__35573\,
            in2 => \N__20620\,
            in3 => \N__48568\,
            lcout => \ALU.madd_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_278_LC_3_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__48567\,
            in1 => \N__20617\,
            in2 => \N__35593\,
            in3 => \N__21094\,
            lcout => \ALU.madd_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_11_l_fx_LC_3_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20832\,
            in1 => \N__27480\,
            in2 => \_gnd_net_\,
            in3 => \N__20855\,
            lcout => \ALU.madd_axb_11_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_273_LC_3_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010000000"
        )
    port map (
            in0 => \N__43394\,
            in1 => \N__43639\,
            in2 => \N__21760\,
            in3 => \N__20803\,
            lcout => \ALU.madd_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a4_b_8_LC_3_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32471\,
            in1 => \N__32377\,
            in2 => \N__36778\,
            in3 => \N__46336\,
            lcout => \ALU.a4_b_8\,
            ltout => \ALU.a4_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_269_LC_3_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__43395\,
            in1 => \N__43638\,
            in2 => \N__20797\,
            in3 => \N__21759\,
            lcout => \ALU.madd_269\,
            ltout => \ALU.madd_269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_289_LC_3_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20787\,
            in2 => \N__20773\,
            in3 => \N__20971\,
            lcout => \ALU.madd_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_185_1_LC_3_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37973\,
            in2 => \_gnd_net_\,
            in3 => \N__52222\,
            lcout => OPEN,
            ltout => \ALU.madd_185_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_185_LC_3_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__21799\,
            in1 => \N__23037\,
            in2 => \N__20752\,
            in3 => \N__22113\,
            lcout => \ALU.madd_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_2_N_2L1_LC_3_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111111111"
        )
    port map (
            in0 => \N__21313\,
            in1 => \N__21292\,
            in2 => \N__24655\,
            in3 => \N__48553\,
            lcout => OPEN,
            ltout => \ALU.g0_2_N_2L1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_2_LC_3_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000001"
        )
    port map (
            in0 => \N__22129\,
            in1 => \N__22009\,
            in2 => \N__20737\,
            in3 => \N__22135\,
            lcout => \ALU.madd_186_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_218_0_tz_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__45206\,
            in1 => \N__40509\,
            in2 => \N__43425\,
            in3 => \N__44551\,
            lcout => \ALU.madd_218_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_228_LC_3_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__22963\,
            in1 => \N__22102\,
            in2 => \N__47456\,
            in3 => \N__48307\,
            lcout => \ALU.madd_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_217_LC_3_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__45205\,
            in1 => \N__40508\,
            in2 => \N__43424\,
            in3 => \N__44550\,
            lcout => \ALU.madd_124_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_13_l_ofx_LC_3_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20955\,
            in1 => \N__21163\,
            in2 => \N__21151\,
            in3 => \N__20940\,
            lcout => \ALU.madd_axb_13_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_335_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010001000"
        )
    port map (
            in0 => \N__20929\,
            in1 => \N__21262\,
            in2 => \N__39850\,
            in3 => \N__48611\,
            lcout => \ALU.madd_335_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_12_ma_LC_3_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20838\,
            in2 => \_gnd_net_\,
            in3 => \N__20856\,
            lcout => \ALU.madd_cry_12_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_294_LC_3_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20911\,
            in1 => \N__21008\,
            in2 => \N__20896\,
            in3 => \N__21078\,
            lcout => \ALU.madd_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_12_l_ofx_LC_3_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__20857\,
            in1 => \N__20839\,
            in2 => \N__21150\,
            in3 => \N__21161\,
            lcout => \ALU.madd_axb_12_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_5_s0_c_RNO_LC_3_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__47255\,
            in1 => \N__53145\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_7_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_341_LC_3_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21708\,
            in1 => \N__22032\,
            in2 => \_gnd_net_\,
            in3 => \N__21691\,
            lcout => \ALU.madd_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_13_ma_LC_3_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21143\,
            lcout => \ALU.madd_cry_13_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_283_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22226\,
            in1 => \N__21029\,
            in2 => \_gnd_net_\,
            in3 => \N__21001\,
            lcout => \ALU.madd_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_218_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__21124\,
            in1 => \N__46103\,
            in2 => \N__21115\,
            in3 => \N__44343\,
            lcout => \ALU.madd_218\,
            ltout => \ALU.madd_218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_346_1_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101011111"
        )
    port map (
            in0 => \N__22225\,
            in1 => \_gnd_net_\,
            in2 => \N__21103\,
            in3 => \N__21028\,
            lcout => \ALU.madd_346_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_10_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__51908\,
            in1 => \N__32666\,
            in2 => \N__36755\,
            in3 => \N__32570\,
            lcout => \ALU.a2_b_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_12_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__21445\,
            in1 => \N__21454\,
            in2 => \N__32894\,
            in3 => \N__48916\,
            lcout => \ALU.a0_b_12\,
            ltout => \ALU.a0_b_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_279_0_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21082\,
            in3 => \N__22224\,
            lcout => \ALU.madd_279_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_349_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010000000"
        )
    port map (
            in0 => \N__22227\,
            in1 => \N__21063\,
            in2 => \N__21036\,
            in3 => \N__21002\,
            lcout => \ALU.madd_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a7_b_5_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__45106\,
            in1 => \N__23106\,
            in2 => \N__36754\,
            in3 => \N__30724\,
            lcout => \ALU.a7_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a12_b_0_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__41276\,
            in1 => \N__32748\,
            in2 => \N__32864\,
            in3 => \N__32719\,
            lcout => \ALU.a12_b_0\,
            ltout => \ALU.a12_b_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_263_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__21228\,
            in1 => \N__40876\,
            in2 => \N__21265\,
            in3 => \N__46780\,
            lcout => \ALU.madd_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a10_b_2_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__29364\,
            in1 => \N__51747\,
            in2 => \N__32863\,
            in3 => \N__33348\,
            lcout => \ALU.a10_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_264_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22205\,
            in1 => \_gnd_net_\,
            in2 => \N__21211\,
            in3 => \N__23262\,
            lcout => OPEN,
            ltout => \ALU.madd_264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_288_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21217\,
            in2 => \N__21247\,
            in3 => \N__22872\,
            lcout => \ALU.madd_288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_259_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__21235\,
            in1 => \N__40877\,
            in2 => \N__21229\,
            in3 => \N__46781\,
            lcout => \ALU.madd_259\,
            ltout => \ALU.madd_259_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_284_0_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23263\,
            in1 => \N__21206\,
            in2 => \N__21190\,
            in3 => \N__22206\,
            lcout => \ALU.madd_284_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIUOP24_10_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24654\,
            in1 => \N__21834\,
            in2 => \_gnd_net_\,
            in3 => \N__21810\,
            lcout => \ALU.b_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIRP8Q_9_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__29486\,
            in1 => \N__31011\,
            in2 => \N__26858\,
            in3 => \N__31146\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIM58R1_9_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__33687\,
            in1 => \N__21968\,
            in2 => \N__21295\,
            in3 => \N__34405\,
            lcout => \ALU.r4_RNIM58R1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_0_rep2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b_0_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56270\,
            ce => \N__56043\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIB9GU_10_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__28123\,
            in1 => \N__26844\,
            in2 => \N__27973\,
            in3 => \N__29487\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIMCFS1_10_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21969\,
            in1 => \N__27937\,
            in2 => \N__21277\,
            in3 => \N__25483\,
            lcout => \ALU.r5_RNIMCFS1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIDBGU_11_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__24539\,
            in1 => \N__29488\,
            in2 => \N__25216\,
            in3 => \N__26845\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIQGFS1_11_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21970\,
            in1 => \N__26119\,
            in2 => \N__21274\,
            in3 => \N__24736\,
            lcout => OPEN,
            ltout => \ALU.r5_RNIQGFS1Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI61Q24_11_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24631\,
            in2 => \N__21271\,
            in3 => \N__21325\,
            lcout => \ALU.b_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIFP8V_10_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__22290\,
            in1 => \N__26856\,
            in2 => \N__29516\,
            in3 => \N__22385\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIUC0U1_10_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__22680\,
            in1 => \N__21943\,
            in2 => \N__21268\,
            in3 => \N__22573\,
            lcout => \ALU.r6_RNIUC0U1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_10_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28192\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r2_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56275\,
            ce => \N__47716\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIHR8V_11_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__29481\,
            in1 => \N__22361\,
            in2 => \N__26860\,
            in3 => \N__24816\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI2H0U1_11_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__24768\,
            in1 => \N__21934\,
            in2 => \N__21328\,
            in3 => \N__22649\,
            lcout => \ALU.r6_RNI2H0U1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_11_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26172\,
            lcout => r2_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56275\,
            ce => \N__47716\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIV5LU_9_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__27581\,
            in1 => \N__29482\,
            in2 => \N__23710\,
            in3 => \N__26857\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIUT042_9_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21935\,
            in1 => \N__27795\,
            in2 => \N__21316\,
            in3 => \N__22255\,
            lcout => \ALU.r6_RNIUT042Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIDP6T_14_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25830\,
            in1 => \N__25857\,
            in2 => \_gnd_net_\,
            in3 => \N__25076\,
            lcout => \ALU.r2_RNIDP6TZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNILPNU_14_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25075\,
            in1 => \N__25798\,
            in2 => \_gnd_net_\,
            in3 => \N__25763\,
            lcout => \ALU.r6_RNILPNUZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIH9VT_14_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26026\,
            in1 => \N__25887\,
            in2 => \_gnd_net_\,
            in3 => \N__25074\,
            lcout => \ALU.r5_RNIH9VTZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_RNI8DSR_14_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__28245\,
            in2 => \_gnd_net_\,
            in3 => \N__29508\,
            lcout => OPEN,
            ltout => \ALU.r1_RNI8DSRZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIFENG2_14_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__24649\,
            in1 => \N__21379\,
            in2 => \N__21373\,
            in3 => \N__21964\,
            lcout => OPEN,
            ltout => \ALU.b_7_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNISO7R4_14_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__32887\,
            in1 => \N__21370\,
            in2 => \N__21364\,
            in3 => \N__21361\,
            lcout => \ALU.b_14\,
            ltout => \ALU.b_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINPPC9_2_14_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21355\,
            in3 => \N__47045\,
            lcout => \ALU.r2_RNINPPC9_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_2_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__25077\,
            in1 => \_gnd_net_\,
            in2 => \N__21991\,
            in3 => \N__32893\,
            lcout => \bZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56280\,
            ce => \N__56041\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s1_c_RNO_0_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34234\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \ALU.r0_12_prm_8_11_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s1_c_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34444\,
            in2 => \N__31120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_11_s1_cy\,
            carryout => \ALU.r0_12_prm_8_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_11_s1_c_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21498\,
            in2 => \N__21352\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_11_s1\,
            carryout => \ALU.r0_12_prm_7_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_11_s1_c_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35145\,
            in2 => \N__22783\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_11_s1\,
            carryout => \ALU.r0_12_prm_6_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_11_s1_c_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21471\,
            in2 => \N__21340\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_11_s1\,
            carryout => \ALU.r0_12_prm_5_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_11_s1_c_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21601\,
            in2 => \N__22711\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_11_s1\,
            carryout => \ALU.r0_12_prm_4_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_11_s1_c_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56398\,
            in2 => \N__55259\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_11_s1\,
            carryout => \ALU.r0_12_prm_3_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_11_s1_c_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35844\,
            in2 => \N__35806\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_11_s1\,
            carryout => \ALU.r0_12_prm_2_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_11_s1_c_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35772\,
            in2 => \N__21394\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \ALU.r0_12_s1_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_11_s0_c_RNI9L4SLH1_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111010000010"
        )
    port map (
            in0 => \N__21574\,
            in1 => \N__27534\,
            in2 => \N__27508\,
            in3 => \N__21385\,
            lcout => \ALU.r0_12_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_11_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26154\,
            lcout => r0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56288\,
            ce => \N__49733\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIHTVA1_12_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__25047\,
            in1 => \N__25170\,
            in2 => \N__21995\,
            in3 => \N__28373\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI05V82_12_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26079\,
            in1 => \N__25453\,
            in2 => \N__21382\,
            in3 => \N__21984\,
            lcout => \ALU.r5_RNI05V82Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNILDOB1_12_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__21980\,
            in1 => \N__23871\,
            in2 => \N__25073\,
            in3 => \N__25317\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI85GA2_12_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__23623\,
            in1 => \N__25257\,
            in2 => \N__21457\,
            in3 => \N__21985\,
            lcout => \ALU.r6_RNI85GA2Z0Z_12\,
            ltout => \ALU.r6_RNI85GA2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIJ1125_12_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21438\,
            in2 => \N__21427\,
            in3 => \N__32891\,
            lcout => \ALU.b_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_0_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25051\,
            lcout => \bZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56292\,
            ce => \N__56040\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIJVVA1_13_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__25046\,
            in1 => \N__25136\,
            in2 => \N__21994\,
            in3 => \N__26211\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI49V82_13_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26050\,
            in1 => \N__25419\,
            in2 => \N__21424\,
            in3 => \N__21979\,
            lcout => \ALU.r5_RNI49V82Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIPDI91_15_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22424\,
            in1 => \N__25600\,
            in2 => \N__22513\,
            in3 => \N__25679\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIH8772_15_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25601\,
            in1 => \N__22619\,
            in2 => \N__21415\,
            in3 => \N__22529\,
            lcout => \ALU.r6_RNIH8772Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_15_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25987\,
            lcout => r2_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56297\,
            ce => \N__47706\,
            sr => \_gnd_net_\
        );

    \ALU.r6_RNINRNU_15_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22620\,
            in1 => \N__22530\,
            in2 => \_gnd_net_\,
            in3 => \N__25067\,
            lcout => \ALU.r6_RNINRNUZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIA0841_0_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23318\,
            in1 => \N__23282\,
            in2 => \_gnd_net_\,
            in3 => \N__25678\,
            lcout => \ALU.r6_RNIA0841Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_0_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29985\,
            in1 => \N__23578\,
            in2 => \N__30364\,
            in3 => \N__28741\,
            lcout => OPEN,
            ltout => \TXbuffer_18_6_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_0_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__39205\,
            in1 => \N__29986\,
            in2 => \N__21526\,
            in3 => \N__23283\,
            lcout => \TXbuffer_RNO_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_7_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__22621\,
            in1 => \N__21511\,
            in2 => \N__30048\,
            in3 => \N__27850\,
            lcout => \TXbuffer_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s0_c_RNO_0_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34549\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \ALU.r0_12_prm_8_11_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s0_c_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34443\,
            in2 => \N__31303\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_11_s0_cy\,
            carryout => \ALU.r0_12_prm_8_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_11_s0_c_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21499\,
            in2 => \N__22792\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_11_s0\,
            carryout => \ALU.r0_12_prm_7_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_11_s0_c_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22798\,
            in2 => \N__35149\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_11_s0\,
            carryout => \ALU.r0_12_prm_6_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_11_s0_c_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22690\,
            in2 => \N__21478\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_11_s0\,
            carryout => \ALU.r0_12_prm_5_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_11_s0_c_inv_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40969\,
            in1 => \N__22696\,
            in2 => \N__21600\,
            in3 => \_gnd_net_\,
            lcout => \ALU.a_i_11\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_11_s0\,
            carryout => \ALU.r0_12_prm_4_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_11_s0_c_inv_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55279\,
            in1 => \N__21583\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_11_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_11_s0\,
            carryout => \ALU.r0_12_prm_3_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_11_s0_c_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34216\,
            in2 => \N__35845\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_11_s0\,
            carryout => \ALU.r0_12_prm_2_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_11_s0_c_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35773\,
            in2 => \N__35731\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \ALU.r0_12_s0_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s0_11_THRU_LUT4_0_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21577\,
            lcout => \ALU.r0_12_s0_11_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_21_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__45188\,
            in1 => \N__32476\,
            in2 => \N__36784\,
            in3 => \N__32375\,
            lcout => \ALU.a4_b_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g1_7_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29220\,
            in1 => \N__29100\,
            in2 => \_gnd_net_\,
            in3 => \N__28978\,
            lcout => OPEN,
            ltout => \ALU.g1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_19_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__22954\,
            in1 => \N__44347\,
            in2 => \N__21562\,
            in3 => \N__24430\,
            lcout => OPEN,
            ltout => \ALU.N_663_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_16_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001100000"
        )
    port map (
            in0 => \N__24175\,
            in1 => \N__21559\,
            in2 => \N__21553\,
            in3 => \N__21548\,
            lcout => \ALU.N_683_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_76_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48291\,
            in1 => \N__40519\,
            in2 => \N__45230\,
            in3 => \N__49348\,
            lcout => OPEN,
            ltout => \ALU.madd_43_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_77_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__44348\,
            in1 => \N__21715\,
            in2 => \N__21718\,
            in3 => \N__42815\,
            lcout => \ALU.madd_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_77_0_tz_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__48290\,
            in1 => \N__40518\,
            in2 => \N__45229\,
            in3 => \N__49349\,
            lcout => \ALU.madd_77_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a6_b_7_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__44704\,
            in1 => \N__36625\,
            in2 => \N__26515\,
            in3 => \N__26437\,
            lcout => \ALU.a6_b_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_345_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__21709\,
            in1 => \N__22033\,
            in2 => \_gnd_net_\,
            in3 => \N__21687\,
            lcout => \ALU.madd_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_159_N_3L3_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101011111"
        )
    port map (
            in0 => \N__22905\,
            in1 => \_gnd_net_\,
            in2 => \N__22939\,
            in3 => \N__22923\,
            lcout => \ALU.madd_159_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_108_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48922\,
            in1 => \N__46307\,
            in2 => \N__44763\,
            in3 => \N__48512\,
            lcout => \ALU.madd_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_140_0_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__44705\,
            in1 => \N__48289\,
            in2 => \N__43643\,
            in3 => \N__49366\,
            lcout => \ALU.madd_140_0\,
            ltout => \ALU.madd_140_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_155_1_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__22922\,
            in1 => \N__22935\,
            in2 => \N__21610\,
            in3 => \N__22904\,
            lcout => \ALU.madd_155_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_144_0_tz_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__48511\,
            in1 => \N__44719\,
            in2 => \N__46348\,
            in3 => \N__48288\,
            lcout => \ALU.madd_144_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_6_1_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22843\,
            in1 => \N__21873\,
            in2 => \_gnd_net_\,
            in3 => \N__31563\,
            lcout => \ALU.g0_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_10_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__21838\,
            in1 => \N__21817\,
            in2 => \N__24653\,
            in3 => \N__48830\,
            lcout => \ALU.a0_b_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_8_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__28999\,
            in1 => \N__29096\,
            in2 => \N__36681\,
            in3 => \N__46308\,
            lcout => \ALU.a5_b_8\,
            ltout => \ALU.a5_b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_325_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__43589\,
            in1 => \N__22041\,
            in2 => \N__21793\,
            in3 => \N__44544\,
            lcout => \ALU.madd_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI435F3_7_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24711\,
            in1 => \N__22447\,
            in2 => \_gnd_net_\,
            in3 => \N__29533\,
            lcout => \ALU.b_7\,
            ltout => \ALU.b_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_7_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__29095\,
            in1 => \N__36621\,
            in2 => \N__21763\,
            in3 => \N__28998\,
            lcout => \ALU.a5_b_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_5_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__28997\,
            in1 => \N__29094\,
            in2 => \N__36680\,
            in3 => \N__45181\,
            lcout => \ALU.a5_b_5\,
            ltout => \ALU.a5_b_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_176_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__43280\,
            in1 => \N__22972\,
            in2 => \N__21745\,
            in3 => \N__40510\,
            lcout => \ALU.madd_176\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_321_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__44545\,
            in1 => \N__22051\,
            in2 => \N__22045\,
            in3 => \N__43590\,
            lcout => \ALU.madd_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIPVKU_6_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__29515\,
            in1 => \N__23463\,
            in2 => \N__26859\,
            in3 => \N__23749\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIIH042_6_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21993\,
            in1 => \N__27883\,
            in2 => \N__22018\,
            in3 => \N__38793\,
            lcout => OPEN,
            ltout => \ALU.r6_RNIIH042Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI6AI74_6_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24642\,
            in2 => \N__22015\,
            in3 => \N__21889\,
            lcout => \ALU.b_6\,
            ltout => \ALU.b_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2BKQ8_1_6_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__43396\,
            in1 => \_gnd_net_\,
            in2 => \N__22012\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r4_RNI2BKQ8_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_2_N_3L3_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37888\,
            in2 => \_gnd_net_\,
            in3 => \N__52139\,
            lcout => \ALU.g0_2_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNILJ8Q_6_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__23496\,
            in1 => \N__29514\,
            in2 => \N__38520\,
            in3 => \N__26846\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIAP7R1_6_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__33783\,
            in1 => \N__21992\,
            in2 => \N__21892\,
            in3 => \N__25360\,
            lcout => \ALU.r4_RNIAP7R1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a9_b_5_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__45128\,
            in1 => \N__30813\,
            in2 => \N__32265\,
            in3 => \N__23229\,
            lcout => \ALU.a9_b_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_14_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47112\,
            in2 => \_gnd_net_\,
            in3 => \N__48915\,
            lcout => \ALU.a0_b_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g2_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__48914\,
            in1 => \N__44489\,
            in2 => \N__51979\,
            in3 => \N__23236\,
            lcout => \ALU.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_2_N_4L5_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__44488\,
            in1 => \N__46009\,
            in2 => \N__43936\,
            in3 => \N__46779\,
            lcout => \ALU.g0_2_N_4L5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_134_0_tz_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__46777\,
            in1 => \N__43899\,
            in2 => \N__46074\,
            in3 => \N__44487\,
            lcout => \ALU.madd_134_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_227_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51940\,
            in1 => \N__48913\,
            in2 => \N__35588\,
            in3 => \N__48509\,
            lcout => \ALU.madd_130_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_130_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__46776\,
            in1 => \_gnd_net_\,
            in2 => \N__46073\,
            in3 => \N__23113\,
            lcout => \ALU.madd_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_171_sx_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43900\,
            in1 => \N__46778\,
            in2 => \N__52228\,
            in3 => \N__46008\,
            lcout => \ALU.madd_171_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_224_0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__51939\,
            in1 => \N__48342\,
            in2 => \N__47435\,
            in3 => \N__48514\,
            lcout => \ALU.madd_224_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_9_s0_c_RNO_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53676\,
            in1 => \N__52143\,
            in2 => \N__53232\,
            in3 => \N__47394\,
            lcout => \ALU.r0_12_prm_6_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_0_l_ofx_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__37828\,
            in1 => \N__48515\,
            in2 => \N__46832\,
            in3 => \N__48921\,
            lcout => \ALU.madd_axb_0_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_0_s1_c_RNO_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__37829\,
            in1 => \N__53675\,
            in2 => \N__53208\,
            in3 => \N__48920\,
            lcout => \ALU.r0_12_prm_6_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_213_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__40932\,
            in1 => \N__23146\,
            in2 => \N__23020\,
            in3 => \N__37827\,
            lcout => \ALU.madd_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a9_b_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__44342\,
            in1 => \N__30814\,
            in2 => \N__36783\,
            in3 => \N__23228\,
            lcout => \ALU.a9_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_167_0_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__45988\,
            in1 => \N__37826\,
            in2 => \N__51806\,
            in3 => \N__43920\,
            lcout => \ALU.madd_167_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNILTKU_5_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__23774\,
            in1 => \N__33140\,
            in2 => \N__24922\,
            in3 => \N__24138\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIBP2O1_5_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__24032\,
            in1 => \N__23964\,
            in2 => \N__22174\,
            in3 => \N__26832\,
            lcout => \ALU.r6_RNIBP2O1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIFAMP_5_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22316\,
            in1 => \N__33303\,
            in2 => \N__37129\,
            in3 => \N__33203\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI0QNE1_5_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__33141\,
            in1 => \N__25927\,
            in2 => \N__22171\,
            in3 => \N__25391\,
            lcout => OPEN,
            ltout => \ALU.r4_RNI0QNE1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKI4F3_5_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22168\,
            in2 => \N__22162\,
            in3 => \N__24710\,
            lcout => \ALU.b_5\,
            ltout => \ALU.b_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI8B628_1_5_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22264\,
            in3 => \N__45512\,
            lcout => \ALU.r4_RNI8B628_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_5_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37209\,
            lcout => r0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56263\,
            ce => \N__49739\,
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIPK3D2_9_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__22253\,
            in1 => \N__30927\,
            in2 => \N__27799\,
            in3 => \N__23419\,
            lcout => \ALU.r6_RNIPK3D2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_9_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34032\,
            lcout => r6_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56267\,
            ce => \N__45853\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_1_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__30386\,
            in1 => \N__31147\,
            in2 => \N__35092\,
            in3 => \N__30038\,
            lcout => OPEN,
            ltout => \TXbuffer_18_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_1_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30039\,
            in1 => \N__34401\,
            in2 => \N__22261\,
            in3 => \N__34369\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_1_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__29675\,
            in1 => \N__49969\,
            in2 => \N__22258\,
            in3 => \N__22237\,
            lcout => \TXbuffer_18_15_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_1_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__30036\,
            in1 => \N__28662\,
            in2 => \N__30398\,
            in3 => \N__23706\,
            lcout => OPEN,
            ltout => \TXbuffer_18_6_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_1_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__22254\,
            in1 => \N__30037\,
            in2 => \N__22240\,
            in3 => \N__29396\,
            lcout => \TXbuffer_RNO_6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__42163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56267\,
            ce => \N__45853\,
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIG3U21_5_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__28788\,
            in1 => \N__22323\,
            in2 => \N__37124\,
            in3 => \N__30557\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI24Q22_5_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__25926\,
            in1 => \N__25393\,
            in2 => \N__22300\,
            in3 => \N__25597\,
            lcout => \ALU.r4_RNI24Q22Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_0_rep2_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \a_0_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56271\,
            ce => \N__56044\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNICBU71_10_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__22289\,
            in2 => \N__22389\,
            in3 => \N__28789\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIP3372_10_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30912\,
            in1 => \N__22679\,
            in2 => \N__22273\,
            in3 => \N__22568\,
            lcout => \ALU.r6_RNIP3372Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIEDU71_11_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__30559\,
            in1 => \N__24815\,
            in2 => \N__22363\,
            in3 => \N__28790\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIT7372_11_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30913\,
            in1 => \N__22650\,
            in2 => \N__22270\,
            in3 => \N__24767\,
            lcout => OPEN,
            ltout => \ALU.r6_RNIT7372Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI8VFH4_11_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29202\,
            in2 => \N__22267\,
            in3 => \N__23671\,
            lcout => \ALU.a_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINJA71_7_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__22406\,
            in1 => \N__30570\,
            in2 => \N__22482\,
            in3 => \N__25004\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIGC3D2_7_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__27842\,
            in1 => \N__38681\,
            in2 => \N__22453\,
            in3 => \N__30885\,
            lcout => \ALU.r6_RNIGC3D2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_7_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38754\,
            lcout => r2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56276\,
            ce => \N__47690\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIP1LU_7_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__33139\,
            in1 => \N__24923\,
            in2 => \N__22481\,
            in3 => \N__22407\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIJ13O1_7_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__38682\,
            in1 => \N__27843\,
            in2 => \N__22450\,
            in3 => \N__26850\,
            lcout => \ALU.r6_RNIJ13O1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_7_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__30044\,
            in1 => \N__22435\,
            in2 => \N__22411\,
            in3 => \N__30305\,
            lcout => OPEN,
            ltout => \TXbuffer_18_6_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_7_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__38683\,
            in1 => \N__30045\,
            in2 => \N__22393\,
            in3 => \N__22534\,
            lcout => \TXbuffer_RNO_6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r3_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35018\,
            lcout => r3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_10_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28189\,
            lcout => r3_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_11_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26155\,
            lcout => r3_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_15_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25993\,
            in3 => \_gnd_net_\,
            lcout => r3_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_7_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38755\,
            lcout => r3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_8_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39525\,
            lcout => r3_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_9_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34026\,
            lcout => r3_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_1_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42155\,
            lcout => r3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56281\,
            ce => \N__47755\,
            sr => \_gnd_net_\
        );

    \ALU.r3_6_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38878\,
            lcout => r3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56285\,
            ce => \N__47762\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_6_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__29968\,
            in1 => \N__25820\,
            in2 => \N__23453\,
            in3 => \N__30303\,
            lcout => OPEN,
            ltout => \TXbuffer_18_13_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_6_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29974\,
            in1 => \N__25796\,
            in2 => \N__22456\,
            in3 => \N__27882\,
            lcout => \TXbuffer_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r3_14_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28312\,
            lcout => r3_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56285\,
            ce => \N__47762\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_2_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29972\,
            in1 => \N__28121\,
            in2 => \N__30354\,
            in3 => \N__33418\,
            lcout => OPEN,
            ltout => \TXbuffer_18_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_2_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29967\,
            in1 => \N__25478\,
            in2 => \N__22606\,
            in3 => \N__34333\,
            lcout => \TXbuffer_RNO_5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_4_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29973\,
            in1 => \N__28374\,
            in2 => \N__30355\,
            in3 => \N__33511\,
            lcout => \TXbuffer_18_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35025\,
            lcout => r6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_10_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28191\,
            lcout => r6_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_11_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r6_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_12_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28440\,
            lcout => r6_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_13_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26277\,
            lcout => r6_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_14_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28309\,
            lcout => r6_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_15_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25976\,
            lcout => r6_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r6_5_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37211\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56289\,
            ce => \N__45842\,
            sr => \_gnd_net_\
        );

    \ALU.r7_0_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35026\,
            lcout => r7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_10_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28190\,
            lcout => r7_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_11_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26176\,
            lcout => r7_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_12_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28446\,
            lcout => r7_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_13_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26279\,
            lcout => r7_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_14_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28311\,
            lcout => r7_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_15_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25972\,
            lcout => r7_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \ALU.r7_5_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37212\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56293\,
            ce => \N__45895\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_6_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29932\,
            in1 => \N__28246\,
            in2 => \N__30324\,
            in3 => \N__38524\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_6_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__33784\,
            in1 => \N__29933\,
            in2 => \N__22756\,
            in3 => \N__26025\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_6_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__49889\,
            in1 => \N__22753\,
            in2 => \N__22741\,
            in3 => \N__22726\,
            lcout => \TXbufferZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56298\,
            ce => \N__56038\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_6_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001010101"
        )
    port map (
            in0 => \N__22738\,
            in1 => \N__25764\,
            in2 => \N__38800\,
            in3 => \N__29931\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_6Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_6_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__29668\,
            in1 => \N__49888\,
            in2 => \N__22729\,
            in3 => \N__22717\,
            lcout => \TXbuffer_18_15_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_6_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23497\,
            in1 => \N__29929\,
            in2 => \N__25723\,
            in3 => \N__30269\,
            lcout => OPEN,
            ltout => \TXbuffer_18_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_6_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29930\,
            in1 => \N__25888\,
            in2 => \N__22720\,
            in3 => \N__25356\,
            lcout => \TXbuffer_RNO_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_11_s1_c_RNO_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54054\,
            in1 => \N__53003\,
            in2 => \N__54779\,
            in3 => \N__40968\,
            lcout => \ALU.r0_12_prm_4_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIAFVE5_11_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__40965\,
            in1 => \N__54596\,
            in2 => \N__53166\,
            in3 => \N__54052\,
            lcout => \ALU.r5_RNIAFVE5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_11_s0_c_RNO_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54595\,
            in1 => \N__35579\,
            in2 => \N__53169\,
            in3 => \N__40966\,
            lcout => \ALU.r0_12_prm_5_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNISP2L9_0_12_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39830\,
            in2 => \_gnd_net_\,
            in3 => \N__41329\,
            lcout => \ALU.r5_RNISP2L9_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_11_s0_c_RNO_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54051\,
            in1 => \N__35578\,
            in2 => \N__53168\,
            in3 => \N__40964\,
            lcout => \ALU.r0_12_prm_6_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_13_s1_c_RNO_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__52996\,
            in1 => \N__35392\,
            in2 => \_gnd_net_\,
            in3 => \N__41464\,
            lcout => \ALU.r0_12_prm_7_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_11_s0_c_RNO_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53004\,
            in1 => \N__35577\,
            in2 => \_gnd_net_\,
            in3 => \N__40963\,
            lcout => \ALU.r0_12_prm_7_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_11_s1_c_RNO_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__40967\,
            in1 => \N__54053\,
            in2 => \N__53167\,
            in3 => \N__35580\,
            lcout => \ALU.r0_12_prm_6_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_5_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__29989\,
            in1 => \N__25426\,
            in2 => \N__22768\,
            in3 => \N__25392\,
            lcout => \TXbuffer_RNO_5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_5_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__29988\,
            in1 => \N__23917\,
            in2 => \N__30359\,
            in3 => \N__23776\,
            lcout => \TXbuffer_18_6_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_5_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__30317\,
            in1 => \N__24101\,
            in2 => \N__24128\,
            in3 => \N__29990\,
            lcout => \TXbuffer_18_13_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_105_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__22993\,
            in1 => \N__48949\,
            in2 => \_gnd_net_\,
            in3 => \N__46363\,
            lcout => \ALU.madd_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a4_b_4_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32472\,
            in1 => \N__32373\,
            in2 => \N__36782\,
            in3 => \N__40520\,
            lcout => \ALU.a4_b_4\,
            ltout => \ALU.a4_b_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_104_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__24183\,
            in1 => \N__45232\,
            in2 => \N__22846\,
            in3 => \N__49350\,
            lcout => \ALU.madd_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_68_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__45504\,
            in1 => \N__24237\,
            in2 => \_gnd_net_\,
            in3 => \N__43930\,
            lcout => \ALU.madd_68\,
            ltout => \ALU.madd_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_82_0_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__24166\,
            in1 => \N__43644\,
            in2 => \N__22822\,
            in3 => \N__48513\,
            lcout => \ALU.madd_82_0\,
            ltout => \ALU.madd_82_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_119_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001000"
        )
    port map (
            in0 => \N__24226\,
            in1 => \N__24217\,
            in2 => \N__22819\,
            in3 => \N__24205\,
            lcout => \ALU.madd_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_100_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__24184\,
            in1 => \N__45233\,
            in2 => \N__38451\,
            in3 => \N__49351\,
            lcout => \ALU.madd_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_68_0_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__37897\,
            in1 => \N__44518\,
            in2 => \N__43355\,
            in3 => \N__46745\,
            lcout => \ALU.madd_68_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_0_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__29079\,
            in1 => \N__29005\,
            in2 => \N__32186\,
            in3 => \N__37898\,
            lcout => \ALU.a5_b_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIS02J4_6_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29219\,
            in1 => \N__26508\,
            in2 => \_gnd_net_\,
            in3 => \N__26436\,
            lcout => \ALU.a_6\,
            ltout => \ALU.a_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_72_0_tz_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__46744\,
            in1 => \N__45454\,
            in2 => \N__22801\,
            in3 => \N__43886\,
            lcout => \ALU.madd_72_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g3_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__49277\,
            in1 => \N__45201\,
            in2 => \N__24469\,
            in3 => \N__40485\,
            lcout => \ALU.g3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_71_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46746\,
            in1 => \N__43279\,
            in2 => \N__45495\,
            in3 => \N__43887\,
            lcout => OPEN,
            ltout => \ALU.madd_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_72_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__37899\,
            in1 => \N__22948\,
            in2 => \N__22942\,
            in3 => \N__44519\,
            lcout => \ALU.madd_72\,
            ltout => \ALU.madd_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_110_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22927\,
            in1 => \_gnd_net_\,
            in2 => \N__22909\,
            in3 => \N__22906\,
            lcout => \ALU.madd_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIVA4L3_8_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24623\,
            in1 => \N__23515\,
            in2 => \_gnd_net_\,
            in3 => \N__22981\,
            lcout => \ALU.b_8\,
            ltout => \ALU.b_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_143_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44675\,
            in1 => \N__48235\,
            in2 => \N__22891\,
            in3 => \N__48472\,
            lcout => \ALU.madd_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_8_s0_c_RNO_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__46317\,
            in1 => \N__53898\,
            in2 => \N__53068\,
            in3 => \N__46080\,
            lcout => \ALU.r0_12_prm_6_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_222_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44678\,
            in1 => \N__46316\,
            in2 => \N__42755\,
            in3 => \N__49236\,
            lcout => OPEN,
            ltout => \ALU.madd_127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_223_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__45505\,
            in1 => \N__43520\,
            in2 => \N__22876\,
            in3 => \N__22999\,
            lcout => \ALU.madd_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_223_0_tz_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__44677\,
            in1 => \N__46315\,
            in2 => \N__42754\,
            in3 => \N__49237\,
            lcout => \ALU.madd_223_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_105_0_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__48473\,
            in1 => \N__43521\,
            in2 => \N__48292\,
            in3 => \N__44676\,
            lcout => \ALU.madd_105_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIU5NK1_8_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__26852\,
            in1 => \N__34069\,
            in2 => \N__33727\,
            in3 => \N__23140\,
            lcout => \ALU.r4_RNIU5NK1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2THO8_0_3_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__31911\,
            in1 => \N__44252\,
            in2 => \N__32264\,
            in3 => \N__31824\,
            lcout => \ALU.un9_addsub_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIUES39_0_1_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001110101100"
        )
    port map (
            in0 => \N__31631\,
            in1 => \N__31721\,
            in2 => \N__32263\,
            in3 => \N__46672\,
            lcout => OPEN,
            ltout => \ALU.un9_addsub_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI90J9E_1_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22975\,
            in3 => \N__48505\,
            lcout => \ALU.r4_RNI90J9EZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a7_b_3_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__44251\,
            in1 => \N__23101\,
            in2 => \N__36685\,
            in3 => \N__30715\,
            lcout => \ALU.a7_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJPM55_2_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27754\,
            in1 => \N__32656\,
            in2 => \_gnd_net_\,
            in3 => \N__32574\,
            lcout => \ALU.a_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIBHM55_1_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31630\,
            in1 => \N__31720\,
            in2 => \_gnd_net_\,
            in3 => \N__27753\,
            lcout => \ALU.a_1\,
            ltout => \ALU.a_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_228_0_tz_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__35581\,
            in1 => \N__51975\,
            in2 => \N__22966\,
            in3 => \N__48759\,
            lcout => \ALU.madd_228_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIUES39_1_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31632\,
            in1 => \N__31722\,
            in2 => \N__46775\,
            in3 => \N__32245\,
            lcout => \ALU.r4_RNIUES39Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIURI55_9_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27751\,
            in1 => \N__30812\,
            in2 => \_gnd_net_\,
            in3 => \N__23224\,
            lcout => \ALU.a_9\,
            ltout => \ALU.a_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_9_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__24403\,
            in1 => \N__32995\,
            in2 => \N__23131\,
            in3 => \N__37831\,
            lcout => \ALU.N_675_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIR1GK3_0_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32744\,
            in1 => \N__24712\,
            in2 => \_gnd_net_\,
            in3 => \N__32708\,
            lcout => \ALU.bZ0Z_0\,
            ltout => \ALU.bZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_130_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__43822\,
            in1 => \N__52102\,
            in2 => \N__23116\,
            in3 => \N__44435\,
            lcout => \ALU.madd_130_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIDBI55_7_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27750\,
            in1 => \N__23100\,
            in2 => \_gnd_net_\,
            in3 => \N__30711\,
            lcout => \ALU.a_7\,
            ltout => \ALU.a_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_133_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46670\,
            in1 => \N__43837\,
            in2 => \N__23053\,
            in3 => \N__46055\,
            lcout => \ALU.madd_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_213_0_tz_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__52104\,
            in1 => \N__43823\,
            in2 => \N__51807\,
            in3 => \N__46671\,
            lcout => \ALU.madd_213_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_209_0_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__43821\,
            in1 => \N__52103\,
            in2 => \N__40970\,
            in3 => \N__37830\,
            lcout => \ALU.madd_209_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a8_b_4_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__36697\,
            in1 => \N__40429\,
            in2 => \N__30621\,
            in3 => \N__23406\,
            lcout => \ALU.a8_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_7_x1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__23405\,
            in1 => \N__30614\,
            in2 => \N__46754\,
            in3 => \N__27741\,
            lcout => OPEN,
            ltout => \ALU.g0_7_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_7_ns_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23239\,
            in3 => \N__43860\,
            lcout => \ALU.madd_76_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a9_b_4_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__40428\,
            in1 => \N__30811\,
            in2 => \N__23230\,
            in3 => \N__36698\,
            lcout => \ALU.a9_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNILJI55_8_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27740\,
            in1 => \N__23404\,
            in2 => \_gnd_net_\,
            in3 => \N__30613\,
            lcout => \ALU.a_8\,
            ltout => \ALU.a_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNICTFPA_9_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__54128\,
            in1 => \N__52122\,
            in2 => \N__23176\,
            in3 => \N__53811\,
            lcout => \ALU.lshift_3_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_224_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__48870\,
            in1 => \N__23173\,
            in2 => \_gnd_net_\,
            in3 => \N__35562\,
            lcout => \ALU.madd_224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_212_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46693\,
            in1 => \N__52121\,
            in2 => \N__43914\,
            in3 => \N__51732\,
            lcout => \ALU.madd_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI6GLV_8_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__39439\,
            in1 => \N__24906\,
            in2 => \N__30663\,
            in3 => \N__33288\,
            lcout => \ALU.b_3_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_0_rep1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24909\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56259\,
            ce => \N__56047\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIUF141_2_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__24905\,
            in2 => \N__23362\,
            in3 => \N__33289\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIE5FT1_2_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__26797\,
            in1 => \N__28088\,
            in2 => \N__23332\,
            in3 => \N__39169\,
            lcout => \ALU.r6_RNIE5FT1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI0I141_3_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__24794\,
            in1 => \N__24907\,
            in2 => \N__23665\,
            in3 => \N__33290\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNII9FT1_3_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__26798\,
            in1 => \N__28059\,
            in2 => \N__23329\,
            in3 => \N__39132\,
            lcout => \ALU.r6_RNII9FT1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIQB141_0_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__28740\,
            in1 => \N__24908\,
            in2 => \N__28839\,
            in3 => \N__33291\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI6TET1_0_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__26799\,
            in1 => \N__23325\,
            in2 => \N__23293\,
            in3 => \N__23290\,
            lcout => \ALU.r6_RNI6TET1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNII5U21_6_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__28781\,
            in1 => \N__38519\,
            in2 => \N__30563\,
            in3 => \N__23483\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI68Q22_6_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__25569\,
            in1 => \N__25352\,
            in2 => \N__23266\,
            in3 => \N__33770\,
            lcout => \ALU.r4_RNI68Q22Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_6_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56264\,
            ce => \N__49746\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIKFA71_5_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23775\,
            in1 => \N__30543\,
            in2 => \N__24139\,
            in3 => \N__28784\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIASIB2_5_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__23957\,
            in1 => \N__24037\,
            in2 => \N__23467\,
            in3 => \N__25571\,
            lcout => \ALU.r6_RNIASIB2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIMHA71_6_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23741\,
            in1 => \N__30541\,
            in2 => \N__23464\,
            in3 => \N__28782\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIE0JB2_6_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__27878\,
            in1 => \N__38786\,
            in2 => \N__23422\,
            in3 => \N__25570\,
            lcout => \ALU.r6_RNIE0JB2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNISNA71_9_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23705\,
            in1 => \N__30542\,
            in2 => \N__27588\,
            in3 => \N__28783\,
            lcout => \ALU.a_6_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIPLA71_8_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23564\,
            in1 => \N__30567\,
            in2 => \N__23548\,
            in3 => \N__25003\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIKG3D2_8_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__27824\,
            in1 => \N__39200\,
            in2 => \N__23413\,
            in3 => \N__30915\,
            lcout => \ALU.r6_RNIKG3D2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_8_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39526\,
            lcout => r2_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56268\,
            ce => \N__47708\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIR3LU_8_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__24924\,
            in1 => \N__33112\,
            in2 => \N__23571\,
            in3 => \N__23546\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIN53O1_8_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__39201\,
            in1 => \N__27825\,
            in2 => \N__23518\,
            in3 => \N__26851\,
            lcout => \ALU.r6_RNIN53O1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIQUF71_1_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__25002\,
            in1 => \N__28652\,
            in2 => \N__28700\,
            in3 => \N__31062\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI7B8D2_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30914\,
            in1 => \N__29439\,
            in2 => \N__23506\,
            in3 => \N__29406\,
            lcout => \ALU.r6_RNI7B8D2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42156\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56268\,
            ce => \N__47708\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIMIB71_10_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__28122\,
            in1 => \N__25000\,
            in2 => \N__27962\,
            in3 => \N__31061\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIVQN52_10_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__27932\,
            in1 => \N__25479\,
            in2 => \N__23503\,
            in3 => \N__30888\,
            lcout => \ALU.r5_RNIVQN52Z0Z_10\,
            ltout => \ALU.r5_RNIVQN52Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI0NFH4_10_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29156\,
            in2 => \N__23500\,
            in3 => \N__36795\,
            lcout => \ALU.a_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_0_rep1_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25001\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \a_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56272\,
            ce => \N__56045\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIOKB71_11_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__24543\,
            in1 => \N__24998\,
            in2 => \N__25196\,
            in3 => \N__31060\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI3VN52_11_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__24734\,
            in1 => \N__26111\,
            in2 => \N__23674\,
            in3 => \N__30886\,
            lcout => \ALU.r5_RNI3VN52Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIU2G71_3_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__24795\,
            in1 => \N__24999\,
            in2 => \N__31084\,
            in3 => \N__23657\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIFJ8D2_3_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__28046\,
            in1 => \N__39128\,
            in2 => \N__23629\,
            in3 => \N__30887\,
            lcout => \ALU.r6_RNIFJ8D2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIEV9A1_12_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__28375\,
            in1 => \N__30889\,
            in2 => \N__25163\,
            in3 => \N__25647\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIS3672_12_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25563\,
            in1 => \N__26078\,
            in2 => \N__23626\,
            in3 => \N__25448\,
            lcout => \ALU.r5_RNIS3672Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIJ7I91_12_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25304\,
            in1 => \N__25564\,
            in2 => \N__23870\,
            in3 => \N__25648\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI5S672_12_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25565\,
            in1 => \N__23621\,
            in2 => \N__23590\,
            in3 => \N__25253\,
            lcout => OPEN,
            ltout => \ALU.r6_RNI5S672Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI9O1J4_12_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29207\,
            in2 => \N__23587\,
            in3 => \N__23584\,
            lcout => \ALU.a_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_2_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__25650\,
            in1 => \_gnd_net_\,
            in2 => \N__25596\,
            in3 => \N__32161\,
            lcout => \aZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56277\,
            ce => \N__56042\,
            sr => \_gnd_net_\
        );

    \a_2_rep2_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32162\,
            in1 => \N__30890\,
            in2 => \_gnd_net_\,
            in3 => \N__25651\,
            lcout => \a_2_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56277\,
            ce => \N__56042\,
            sr => \_gnd_net_\
        );

    \a_0_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56277\,
            ce => \N__56042\,
            sr => \_gnd_net_\
        );

    \ALU.r2_12_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28441\,
            lcout => r2_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56282\,
            ce => \N__47686\,
            sr => \_gnd_net_\
        );

    \ALU.r2_14_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r2_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56282\,
            ce => \N__47686\,
            sr => \_gnd_net_\
        );

    \ALU.r2_5_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37210\,
            lcout => r2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56282\,
            ce => \N__47686\,
            sr => \_gnd_net_\
        );

    \ALU.r2_6_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38873\,
            lcout => r2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56282\,
            ce => \N__47686\,
            sr => \_gnd_net_\
        );

    \ALU.r2_9_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34033\,
            lcout => r2_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56282\,
            ce => \N__47686\,
            sr => \_gnd_net_\
        );

    \ALU.r2_3_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50200\,
            lcout => r2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56282\,
            ce => \N__47686\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s1_c_RNO_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37519\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \ALU.r0_12_prm_8_15_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s1_c_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36031\,
            in2 => \N__31201\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_15_s1_cy\,
            carryout => \ALU.r0_12_prm_8_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_15_s1_c_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35986\,
            in2 => \N__23836\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_15_s1\,
            carryout => \ALU.r0_12_prm_7_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_15_s1_c_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35949\,
            in2 => \N__23821\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_15_s1\,
            carryout => \ALU.r0_12_prm_6_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_15_s1_c_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35911\,
            in2 => \N__37540\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_15_s1\,
            carryout => \ALU.r0_12_prm_5_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_15_s1_c_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35881\,
            in2 => \N__23806\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_15_s1\,
            carryout => \ALU.r0_12_prm_4_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_15_s1_c_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55216\,
            in2 => \N__56413\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_15_s1\,
            carryout => \ALU.r0_12_prm_3_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_15_s1_c_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36259\,
            in2 => \N__31249\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_15_s1\,
            carryout => \ALU.r0_12_prm_2_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_15_s1_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37297\,
            in2 => \N__37252\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \ALU.r0_12_s1_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_15_s0_c_RNI2DJ0GB2_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111010000010"
        )
    port map (
            in0 => \N__36190\,
            in1 => \N__23791\,
            in2 => \N__27358\,
            in3 => \N__23779\,
            lcout => \ALU.r0_12_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_15_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25968\,
            lcout => r0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56290\,
            ce => \N__49717\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIHPP81_13_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__26198\,
            in1 => \N__25598\,
            in2 => \N__25137\,
            in3 => \N__25680\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI10M52_13_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__26045\,
            in1 => \N__25412\,
            in2 => \N__23920\,
            in3 => \N__25602\,
            lcout => \ALU.r5_RNI10M52Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIL9I91_13_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__23916\,
            in1 => \N__25599\,
            in2 => \N__24102\,
            in3 => \N__25681\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI90772_13_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__23981\,
            in1 => \N__24071\,
            in2 => \N__23887\,
            in3 => \N__25603\,
            lcout => OPEN,
            ltout => \ALU.r6_RNI90772Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIIOHH4_13_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29206\,
            in2 => \N__23884\,
            in3 => \N__23881\,
            lcout => \ALU.a_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIPV8A9_13_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53900\,
            in1 => \N__47003\,
            in2 => \_gnd_net_\,
            in3 => \N__41445\,
            lcout => OPEN,
            ltout => \ALU.r5_RNIPV8A9Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNILM5AE_15_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__53955\,
            in1 => \N__54383\,
            in2 => \N__23875\,
            in3 => \N__40142\,
            lcout => \ALU.r5_RNILM5AEZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r3_4_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39091\,
            lcout => r3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56299\,
            ce => \N__47764\,
            sr => \_gnd_net_\
        );

    \ALU.r3_12_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28423\,
            lcout => r3_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56299\,
            ce => \N__47764\,
            sr => \_gnd_net_\
        );

    \ALU.r3_5_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37216\,
            lcout => r3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56299\,
            ce => \N__47764\,
            sr => \_gnd_net_\
        );

    \ALU.r3_13_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26242\,
            lcout => r3_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56299\,
            ce => \N__47764\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_5_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30049\,
            in1 => \N__24079\,
            in2 => \N__24049\,
            in3 => \N__24036\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_6Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_5_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__29669\,
            in1 => \N__23998\,
            in2 => \N__23992\,
            in3 => \N__49925\,
            lcout => \TXbuffer_18_15_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_5_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__30050\,
            in1 => \N__23989\,
            in2 => \N__23965\,
            in3 => \N__23932\,
            lcout => \TXbuffer_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_5_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__26049\,
            in1 => \N__23926\,
            in2 => \N__30080\,
            in3 => \N__25922\,
            lcout => \TXbuffer_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_5_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__37125\,
            in1 => \N__29987\,
            in2 => \N__30394\,
            in3 => \N__25138\,
            lcout => \TXbuffer_18_10_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_4_c_RNO_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__40487\,
            in1 => \N__53212\,
            in2 => \N__53812\,
            in3 => \N__42788\,
            lcout => \ALU.r0_12_prm_6_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_6_s1_c_RNO_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54555\,
            in1 => \N__53590\,
            in2 => \N__53250\,
            in3 => \N__43283\,
            lcout => \ALU.r0_12_prm_4_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_81_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000011000000"
        )
    port map (
            in0 => \N__45500\,
            in1 => \N__24238\,
            in2 => \N__24165\,
            in3 => \N__43929\,
            lcout => \ALU.madd_46_0\,
            ltout => \ALU.madd_46_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_115_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__24216\,
            in1 => \N__24204\,
            in2 => \N__24193\,
            in3 => \N__24190\,
            lcout => \ALU.madd_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_3_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__29078\,
            in1 => \N__29009\,
            in2 => \N__36753\,
            in3 => \N__44308\,
            lcout => \ALU.a5_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2BKQ8_6_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43648\,
            in2 => \_gnd_net_\,
            in3 => \N__43282\,
            lcout => \ALU.un14_log_0_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g2_0_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__44309\,
            in1 => \N__43281\,
            in2 => \N__45513\,
            in3 => \N__40486\,
            lcout => \ALU.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_7_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48760\,
            in2 => \_gnd_net_\,
            in3 => \N__44765\,
            lcout => \ALU.a0_b_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_34_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__48762\,
            in1 => \N__26590\,
            in2 => \N__45257\,
            in3 => \N__26689\,
            lcout => \ALU.madd_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_33_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__24289\,
            in1 => \N__49288\,
            in2 => \N__24148\,
            in3 => \N__43896\,
            lcout => \ALU.madd_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_38_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010000000"
        )
    port map (
            in0 => \N__48763\,
            in1 => \N__26589\,
            in2 => \N__45258\,
            in3 => \N__26688\,
            lcout => \ALU.madd_38\,
            ltout => \ALU.madd_38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_60_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26643\,
            in2 => \N__24280\,
            in3 => \N__26661\,
            lcout => \ALU.madd_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_87_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__27163\,
            in1 => \N__27154\,
            in2 => \_gnd_net_\,
            in3 => \N__27139\,
            lcout => \ALU.madd_87\,
            ltout => \ALU.madd_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_120_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26568\,
            in2 => \N__24277\,
            in3 => \N__26556\,
            lcout => \ALU.madd_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_6_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__48761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43606\,
            lcout => \ALU.a0_b_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_92_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011101000"
        )
    port map (
            in0 => \N__24250\,
            in1 => \N__24265\,
            in2 => \N__27127\,
            in3 => \N__24271\,
            lcout => \ALU.madd_92\,
            ltout => \ALU.madd_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_7_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__24352\,
            in1 => \N__26680\,
            in2 => \N__24274\,
            in3 => \N__26599\,
            lcout => \ALU.madd_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_78_0_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__48793\,
            in1 => \N__44790\,
            in2 => \N__43665\,
            in3 => \N__48510\,
            lcout => \ALU.madd_78_0\,
            ltout => \ALU.madd_78_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_88_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24264\,
            in1 => \N__27123\,
            in2 => \N__24253\,
            in3 => \N__24249\,
            lcout => \ALU.madd_332\,
            ltout => \ALU.madd_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_6_l_ofx_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__26598\,
            in1 => \N__28892\,
            in2 => \N__24241\,
            in3 => \N__28876\,
            lcout => \ALU.madd_axb_6_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNII0MP4_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__24376\,
            in1 => \N__28753\,
            in2 => \N__29208\,
            in3 => \N__27700\,
            lcout => \ALU.aZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI6N1R4_4_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32361\,
            in1 => \N__32453\,
            in2 => \_gnd_net_\,
            in3 => \N__29183\,
            lcout => \ALU.a_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_8_l_fx_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__24358\,
            in2 => \N__27223\,
            in3 => \N__24351\,
            lcout => \ALU.madd_axb_8_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_0_ma_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48792\,
            in2 => \_gnd_net_\,
            in3 => \N__46680\,
            lcout => \ALU.madd_cry_0_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_4_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__32675\,
            in1 => \N__40433\,
            in2 => \N__32173\,
            in3 => \N__32589\,
            lcout => \ALU.a2_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJQGK3_3_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24329\,
            in1 => \N__24706\,
            in2 => \_gnd_net_\,
            in3 => \N__33030\,
            lcout => \ALU.b_3\,
            ltout => \ALU.b_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2THO8_3_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110100101"
        )
    port map (
            in0 => \N__31797\,
            in1 => \N__31902\,
            in2 => \N__24310\,
            in3 => \N__32129\,
            lcout => \ALU.un2_addsub_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI0TRV3_1_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__29374\,
            in1 => \N__26731\,
            in2 => \N__28636\,
            in3 => \N__24705\,
            lcout => \ALU.b_1\,
            ltout => \ALU.b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a4_b_1_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__32102\,
            in1 => \N__32460\,
            in2 => \N__24292\,
            in3 => \N__32362\,
            lcout => \ALU.a4_b_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIS1N55_3_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27752\,
            in1 => \N__31901\,
            in2 => \_gnd_net_\,
            in3 => \N__31796\,
            lcout => \ALU.a_3\,
            ltout => \ALU.a_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g1_1_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24462\,
            in1 => \N__40432\,
            in2 => \N__24433\,
            in3 => \N__45218\,
            lcout => \ALU.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNICA4F3_4_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33438\,
            in1 => \N__24701\,
            in2 => \_gnd_net_\,
            in3 => \N__24862\,
            lcout => \ALU.b_4\,
            ltout => \ALU.b_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_214_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__44248\,
            in1 => \N__45989\,
            in2 => \N__24418\,
            in3 => \N__44446\,
            lcout => \ALU.madd_214_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_373_0_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__40431\,
            in1 => \N__44250\,
            in2 => \N__51839\,
            in3 => \N__40986\,
            lcout => \ALU.madd_373_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIBIGK3_2_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24700\,
            in1 => \N__29360\,
            in2 => \_gnd_net_\,
            in3 => \N__33347\,
            lcout => \ALU.b_2\,
            ltout => \ALU.b_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_11_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__44449\,
            in1 => \N__46182\,
            in2 => \N__24406\,
            in3 => \N__46678\,
            lcout => \ALU.madd_134_0_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2QU6A_6_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__53421\,
            in1 => \N__43408\,
            in2 => \N__54215\,
            in3 => \N__44447\,
            lcout => \ALU.lshift_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIC5NE1_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__27685\,
            in1 => \N__33142\,
            in2 => \N__27637\,
            in3 => \N__33523\,
            lcout => \ALU.r4_RNIC5NE1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_172_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__44249\,
            in1 => \N__40430\,
            in2 => \N__43431\,
            in3 => \N__44448\,
            lcout => \ALU.madd_172_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_368_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__37886\,
            in1 => \N__27341\,
            in2 => \N__24496\,
            in3 => \N__47001\,
            lcout => \ALU.madd_368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a12_b_2_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__41315\,
            in1 => \N__29359\,
            in2 => \N__32841\,
            in3 => \N__33349\,
            lcout => \ALU.a12_b_2\,
            ltout => \ALU.a12_b_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_372_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__37887\,
            in1 => \N__27342\,
            in2 => \N__24487\,
            in3 => \N__47002\,
            lcout => \ALU.madd_372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a13_b_1_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__41548\,
            in1 => \N__46710\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.a13_b_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_368_0_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__41314\,
            in1 => \N__37885\,
            in2 => \N__47041\,
            in3 => \N__43862\,
            lcout => \ALU.madd_368_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g1_2_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29215\,
            in1 => \N__32447\,
            in2 => \_gnd_net_\,
            in3 => \N__32350\,
            lcout => \ALU.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_311_0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__40931\,
            in1 => \N__37884\,
            in2 => \N__41565\,
            in3 => \N__43861\,
            lcout => \ALU.madd_311_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_2_rep2_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__32816\,
            in1 => \N__25097\,
            in2 => \_gnd_net_\,
            in3 => \N__26827\,
            lcout => \b_2_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \b_1_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32815\,
            lcout => \bZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \b_fast_2_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__32817\,
            in1 => \N__25098\,
            in2 => \_gnd_net_\,
            in3 => \N__33295\,
            lcout => \b_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \b_fast_1_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25099\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26874\,
            lcout => \b_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \b_1_rep1_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25096\,
            in2 => \_gnd_net_\,
            in3 => \N__24699\,
            lcout => \b_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \b_1_rep2_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__24581\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b_1_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \params_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53356\,
            in2 => \_gnd_net_\,
            in3 => \N__54129\,
            lcout => \paramsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \params_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__53357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \paramsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => \N__56049\,
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIMQ992_3_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__33056\,
            in1 => \N__30924\,
            in2 => \N__33603\,
            in3 => \N__30583\,
            lcout => \ALU.r4_RNIMQ992Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_3_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56260\,
            ce => \N__47809\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_3_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110101"
        )
    port map (
            in0 => \N__35053\,
            in1 => \N__24547\,
            in2 => \N__30414\,
            in3 => \N__30064\,
            lcout => OPEN,
            ltout => \TXbuffer_18_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30065\,
            in1 => \N__24735\,
            in2 => \N__24850\,
            in3 => \N__33057\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_5Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__29676\,
            in1 => \N__49968\,
            in2 => \N__24847\,
            in3 => \N__24742\,
            lcout => \TXbuffer_18_15_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_3_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__30062\,
            in1 => \N__24823\,
            in2 => \N__30395\,
            in3 => \N__24799\,
            lcout => OPEN,
            ltout => \TXbuffer_18_6_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_3_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__24772\,
            in1 => \N__39139\,
            in2 => \N__24745\,
            in3 => \N__30063\,
            lcout => \TXbuffer_RNO_6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_11_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26183\,
            lcout => r4_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56260\,
            ce => \N__47809\,
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIUF9K8_1_10_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52000\,
            in2 => \_gnd_net_\,
            in3 => \N__51652\,
            lcout => \ALU.r5_RNIUF9K8_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_2_rep1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__32043\,
            in1 => \_gnd_net_\,
            in2 => \N__25692\,
            in3 => \N__30568\,
            lcout => \a_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \a_1_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25682\,
            in2 => \_gnd_net_\,
            in3 => \N__32042\,
            lcout => \aZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \a_fast_2_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__32044\,
            in1 => \_gnd_net_\,
            in2 => \N__25693\,
            in3 => \N__31066\,
            lcout => \a_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \a_fast_1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25684\,
            in2 => \_gnd_net_\,
            in3 => \N__27734\,
            lcout => \a_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \a_1_rep1_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__25691\,
            in1 => \N__29160\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \a_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \a_1_rep2_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25683\,
            in2 => \_gnd_net_\,
            in3 => \N__36563\,
            lcout => \a_1_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \b_2_rep1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__33113\,
            in1 => \N__25102\,
            in2 => \_gnd_net_\,
            in3 => \N__32834\,
            lcout => \b_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56265\,
            ce => \N__56046\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIHDA71_4_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__25011\,
            in1 => \N__30553\,
            in2 => \N__25287\,
            in3 => \N__24953\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI403D2_4_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__39000\,
            in1 => \N__28017\,
            in2 => \N__24961\,
            in3 => \N__30925\,
            lcout => \ALU.r6_RNI403D2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_4_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56269\,
            ce => \N__47664\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIJRKU_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25275\,
            in1 => \N__33111\,
            in2 => \N__24957\,
            in3 => \N__24925\,
            lcout => OPEN,
            ltout => \ALU.b_6_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNI7L2O1_4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__28016\,
            in1 => \N__38999\,
            in2 => \N__24865\,
            in3 => \N__26828\,
            lcout => \ALU.r6_RNI7L2O1Z0Z_4\,
            ltout => \ALU.r6_RNI7L2O1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIE2CL3_4_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32830\,
            in2 => \N__25321\,
            in3 => \N__33439\,
            lcout => \ALU.b_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_8_4_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__30046\,
            in1 => \N__25318\,
            in2 => \N__25288\,
            in3 => \N__30309\,
            lcout => OPEN,
            ltout => \TXbuffer_18_6_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_6_4_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__39001\,
            in1 => \N__30047\,
            in2 => \N__25264\,
            in3 => \N__25261\,
            lcout => \TXbuffer_RNO_6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_10_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28160\,
            lcout => r1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r1_11_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26184\,
            lcout => r1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r1_12_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28447\,
            in3 => \_gnd_net_\,
            lcout => r1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r1_13_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26280\,
            lcout => r1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r1_15_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25989\,
            lcout => r1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r1_8_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39523\,
            lcout => r1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r1_9_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34031\,
            lcout => r1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56273\,
            ce => \N__47560\,
            sr => \_gnd_net_\
        );

    \ALU.r4_0_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35000\,
            lcout => r4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_10_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28159\,
            lcout => r4_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_12_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28442\,
            lcout => r4_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_13_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26278\,
            lcout => r4_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_14_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28308\,
            lcout => r4_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_15_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25988\,
            lcout => r4_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_5_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r4_6_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38872\,
            lcout => r4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56278\,
            ce => \N__47802\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNIJRP81_14_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25706\,
            in1 => \N__25575\,
            in2 => \N__28238\,
            in3 => \N__25662\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI54M52_14_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25576\,
            in1 => \N__26021\,
            in2 => \N__25891\,
            in3 => \N__25880\,
            lcout => \ALU.r5_RNI54M52Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINBI91_14_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__25844\,
            in1 => \N__25578\,
            in2 => \N__25831\,
            in3 => \N__25664\,
            lcout => OPEN,
            ltout => \ALU.a_6_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNID4772_14_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25580\,
            in1 => \N__25797\,
            in2 => \N__25768\,
            in3 => \N__25765\,
            lcout => OPEN,
            ltout => \ALU.r6_RNID4772Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIR0IH4_14_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36664\,
            in2 => \N__25735\,
            in3 => \N__25732\,
            lcout => \ALU.a_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_14_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28295\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56283\,
            ce => \N__49730\,
            sr => \_gnd_net_\
        );

    \ALU.r1_RNILTP81_15_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__30107\,
            in1 => \N__25577\,
            in2 => \N__30479\,
            in3 => \N__25663\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI98M52_15_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__25579\,
            in1 => \N__30434\,
            in2 => \N__25495\,
            in3 => \N__29708\,
            lcout => \ALU.r5_RNI98M52Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35009\,
            lcout => r5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_10_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28176\,
            lcout => r5_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_11_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26185\,
            lcout => r5_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_12_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28427\,
            lcout => r5_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_13_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26261\,
            lcout => r5_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_14_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28294\,
            lcout => r5_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_15_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25986\,
            in3 => \_gnd_net_\,
            lcout => r5_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r5_5_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37208\,
            lcout => r5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56286\,
            ce => \N__45805\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s0_c_RNO_0_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39658\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \ALU.r0_12_prm_8_13_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s0_c_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36160\,
            in2 => \N__35713\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_13_s0_cy\,
            carryout => \ALU.r0_12_prm_8_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_13_s0_c_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31476\,
            in2 => \N__26335\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_13_s0\,
            carryout => \ALU.r0_12_prm_7_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_13_s0_c_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31432\,
            in2 => \N__26350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_13_s0\,
            carryout => \ALU.r0_12_prm_6_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_13_s0_c_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26359\,
            in2 => \N__31398\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_13_s0\,
            carryout => \ALU.r0_12_prm_5_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_13_s0_c_inv_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31359\,
            in2 => \N__26371\,
            in3 => \N__41468\,
            lcout => \ALU.a_i_13\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_13_s0\,
            carryout => \ALU.r0_12_prm_4_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_13_s0_c_inv_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26290\,
            in2 => \_gnd_net_\,
            in3 => \N__55220\,
            lcout => \ALU.r0_12_prm_3_13_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_13_s0\,
            carryout => \ALU.r0_12_prm_3_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_13_s0_c_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34597\,
            in2 => \N__31234\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_13_s0\,
            carryout => \ALU.r0_12_prm_2_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_13_s0_c_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35302\,
            in2 => \N__34624\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_16_0_\,
            carryout => \ALU.r0_12_s0_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_13_s0_c_RNIMPTBGM2_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27412\,
            in1 => \N__31513\,
            in2 => \_gnd_net_\,
            in3 => \N__26284\,
            lcout => \ALU.r0_12_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_13_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26241\,
            lcout => r0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56294\,
            ce => \N__49726\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_13_s1_c_RNO_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__41500\,
            in1 => \N__54592\,
            in2 => \N__54061\,
            in3 => \N__52982\,
            lcout => \ALU.r0_12_prm_4_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIK81F5_13_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54028\,
            in1 => \N__54594\,
            in2 => \N__53163\,
            in3 => \N__41504\,
            lcout => \ALU.r5_RNIK81F5Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_13_s0_c_RNO_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110100101"
        )
    port map (
            in0 => \N__41503\,
            in1 => \N__52985\,
            in2 => \N__35427\,
            in3 => \N__54593\,
            lcout => \ALU.r0_12_prm_5_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_12_s1_c_RNO_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54590\,
            in1 => \N__39859\,
            in2 => \N__53160\,
            in3 => \N__41316\,
            lcout => \ALU.r0_12_prm_5_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_13_s0_c_RNO_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100000101"
        )
    port map (
            in0 => \N__41502\,
            in1 => \N__52983\,
            in2 => \N__35426\,
            in3 => \N__54027\,
            lcout => \ALU.r0_12_prm_6_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_13_s1_c_RNO_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54026\,
            in1 => \N__35410\,
            in2 => \N__53161\,
            in3 => \N__41498\,
            lcout => \ALU.r0_12_prm_6_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_13_s0_c_RNO_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001011111"
        )
    port map (
            in0 => \N__41501\,
            in1 => \_gnd_net_\,
            in2 => \N__35425\,
            in3 => \N__52984\,
            lcout => \ALU.r0_12_prm_7_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_13_s1_c_RNO_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54591\,
            in1 => \N__35411\,
            in2 => \N__53162\,
            in3 => \N__41499\,
            lcout => \ALU.r0_12_prm_5_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_9_l_ofx_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__26545\,
            in1 => \N__26533\,
            in2 => \N__26323\,
            in3 => \N__26305\,
            lcout => \ALU.madd_axb_9_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_9_ma_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26544\,
            in2 => \_gnd_net_\,
            in3 => \N__26532\,
            lcout => \ALU.madd_cry_9_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_124_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26581\,
            in1 => \N__26575\,
            in2 => \_gnd_net_\,
            in3 => \N__26557\,
            lcout => \ALU.madd_124\,
            ltout => \ALU.madd_124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_165_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26536\,
            in3 => \N__26531\,
            lcout => \ALU.madd_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_0_s1_c_RNO_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110001100011"
        )
    port map (
            in0 => \N__53946\,
            in1 => \N__48910\,
            in2 => \N__55955\,
            in3 => \N__38007\,
            lcout => \ALU.r0_12_prm_1_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a6_b_6_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__26514\,
            in1 => \N__43607\,
            in2 => \N__32261\,
            in3 => \N__26447\,
            lcout => \ALU.a6_b_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_0_s0_c_RNO_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110001100011"
        )
    port map (
            in0 => \N__53948\,
            in1 => \N__48912\,
            in2 => \N__55956\,
            in3 => \N__38008\,
            lcout => \ALU.r0_12_prm_1_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIKG5N5_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__48911\,
            in1 => \N__53947\,
            in2 => \N__53257\,
            in3 => \N__54556\,
            lcout => \ALU.r2_RNIKG5N5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_29_0_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__42723\,
            in1 => \N__37967\,
            in2 => \N__45496\,
            in3 => \N__46748\,
            lcout => \ALU.madd_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_14_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__37969\,
            in1 => \N__40731\,
            in2 => \N__26383\,
            in3 => \N__42725\,
            lcout => \ALU.madd_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_1_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__31935\,
            in1 => \N__31828\,
            in2 => \N__36771\,
            in3 => \N__46747\,
            lcout => \ALU.a3_b_1\,
            ltout => \ALU.a3_b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_18_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__37968\,
            in1 => \N__40730\,
            in2 => \N__26374\,
            in3 => \N__42724\,
            lcout => \ALU.madd_18\,
            ltout => \ALU.madd_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_43_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011101000"
        )
    port map (
            in0 => \N__29562\,
            in1 => \N__28593\,
            in2 => \N__26695\,
            in3 => \N__28617\,
            lcout => \ALU.madd_43\,
            ltout => \ALU.madd_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_5_l_fx_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__26725\,
            in1 => \N__26628\,
            in2 => \N__26692\,
            in3 => \N__29266\,
            lcout => \ALU.madd_axb_5_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_3_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32685\,
            in1 => \N__32593\,
            in2 => \N__36770\,
            in3 => \N__44313\,
            lcout => \ALU.a2_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_94_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100000000000"
        )
    port map (
            in0 => \N__26724\,
            in1 => \N__26611\,
            in2 => \N__26632\,
            in3 => \N__26679\,
            lcout => \ALU.madd_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_56_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26662\,
            in1 => \N__26650\,
            in2 => \_gnd_net_\,
            in3 => \N__26644\,
            lcout => \ALU.madd_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_51_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__44276\,
            in1 => \N__26902\,
            in2 => \N__26893\,
            in3 => \N__49254\,
            lcout => \ALU.madd_51\,
            ltout => \ALU.madd_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_65_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26718\,
            in2 => \N__26614\,
            in3 => \N__26610\,
            lcout => \ALU.madd_331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a1_b_4_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__31647\,
            in1 => \N__31738\,
            in2 => \N__36765\,
            in3 => \N__40531\,
            lcout => \ALU.a1_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_73_0_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__40532\,
            in1 => \N__49238\,
            in2 => \N__42787\,
            in3 => \N__44274\,
            lcout => OPEN,
            ltout => \ALU.madd_73_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_73_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__45190\,
            in1 => \_gnd_net_\,
            in2 => \N__26905\,
            in3 => \N__48361\,
            lcout => \ALU.madd_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a1_b_5_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__31739\,
            in1 => \N__45189\,
            in2 => \N__32185\,
            in3 => \N__31648\,
            lcout => \ALU.a1_b_5\,
            ltout => \ALU.a1_b_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_55_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__44275\,
            in1 => \N__26889\,
            in2 => \N__26878\,
            in3 => \N__49253\,
            lcout => \ALU.madd_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_2_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__43818\,
            in1 => \N__36734\,
            in2 => \N__32591\,
            in3 => \N__32677\,
            lcout => \ALU.a2_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIMTDQ_1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34368\,
            in1 => \N__33202\,
            in2 => \_gnd_net_\,
            in3 => \N__33663\,
            lcout => OPEN,
            ltout => \ALU.r4_RNIMTDQZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI73OM1_1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__26875\,
            in1 => \N__26833\,
            in2 => \N__26734\,
            in3 => \N__32935\,
            lcout => \ALU.b_7_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_46_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__42727\,
            in1 => \N__35116\,
            in2 => \N__26707\,
            in3 => \N__43820\,
            lcout => \ALU.madd_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a5_b_1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__29080\,
            in1 => \N__32106\,
            in2 => \N__29014\,
            in3 => \N__46679\,
            lcout => \ALU.a5_b_1\,
            ltout => \ALU.a5_b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_50_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011000000"
        )
    port map (
            in0 => \N__42726\,
            in1 => \N__35115\,
            in2 => \N__27166\,
            in3 => \N__43819\,
            lcout => \ALU.madd_50\,
            ltout => \ALU.madd_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_83_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27153\,
            in2 => \N__27142\,
            in3 => \N__27138\,
            lcout => \ALU.madd_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIHCHO8_2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001010011"
        )
    port map (
            in0 => \N__32676\,
            in1 => \N__32579\,
            in2 => \N__32174\,
            in3 => \N__43817\,
            lcout => \ALU.un2_addsub_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_2_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__27115\,
            in1 => \N__27895\,
            in2 => \N__49978\,
            in3 => \N__27097\,
            lcout => \TXbufferZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56253\,
            ce => \N__56051\,
            sr => \_gnd_net_\
        );

    \clkdiv_RNIQAHO1_0_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27082\,
            in1 => \N__27055\,
            in2 => \N__27031\,
            in3 => \N__26989\,
            lcout => params5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_3_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26937\,
            in1 => \N__28524\,
            in2 => \_gnd_net_\,
            in3 => \N__29331\,
            lcout => \ALU.madd_axb_3\,
            ltout => \ALU.madd_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_3_s_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26941\,
            in3 => \N__38544\,
            lcout => \ALU.mult_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_28_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26938\,
            in1 => \N__28525\,
            in2 => \_gnd_net_\,
            in3 => \N__29332\,
            lcout => \ALU.madd_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_0_0_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26926\,
            in2 => \N__26917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \ALU.madd_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_0_THRU_LUT4_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42898\,
            in2 => \_gnd_net_\,
            in3 => \N__27268\,
            lcout => \ALU.madd_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_0\,
            carryout => \ALU.madd_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_1_THRU_LUT4_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50052\,
            in2 => \_gnd_net_\,
            in3 => \N__27265\,
            lcout => \ALU.madd_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_1\,
            carryout => \ALU.madd_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_2_THRU_LUT4_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38559\,
            in2 => \_gnd_net_\,
            in3 => \N__27262\,
            lcout => \ALU.madd_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_2\,
            carryout => \ALU.madd_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_4_s_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28563\,
            in2 => \N__28552\,
            in3 => \N__27259\,
            lcout => \ALU.mult_5\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_3\,
            carryout => \ALU.madd_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_5_s_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29262\,
            in2 => \N__27256\,
            in3 => \N__27244\,
            lcout => \ALU.mult_6\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_4\,
            carryout => \ALU.madd_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_6_0_s_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27241\,
            in2 => \N__28855\,
            in3 => \N__27229\,
            lcout => \ALU.mult_7\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_5\,
            carryout => \ALU.madd_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_6_THRU_LUT4_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39561\,
            in2 => \_gnd_net_\,
            in3 => \N__27226\,
            lcout => \ALU.madd_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_6\,
            carryout => \ALU.madd_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_8_s_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27219\,
            in2 => \N__27196\,
            in3 => \N__27181\,
            lcout => \ALU.mult_9\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \ALU.madd_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_9_0_s_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27178\,
            in2 => \N__27550\,
            in3 => \N__27538\,
            lcout => \ALU.mult_10\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_8\,
            carryout => \ALU.madd_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_9_THRU_LUT4_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27535\,
            in3 => \N__27490\,
            lcout => \ALU.madd_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_9\,
            carryout => \ALU.madd_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_11_s_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27487\,
            in2 => \N__27460\,
            in3 => \N__27445\,
            lcout => \ALU.mult_12\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_10\,
            carryout => \ALU.madd_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_12_0_s_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27442\,
            in2 => \N__27430\,
            in3 => \N__27397\,
            lcout => \ALU.mult_13\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_11\,
            carryout => \ALU.madd_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_13_0_s_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27394\,
            in2 => \N__27379\,
            in3 => \N__27364\,
            lcout => \ALU.mult_14\,
            ltout => OPEN,
            carryin => \ALU.madd_cry_12\,
            carryout => \ALU.madd_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.madd_cry_13_THRU_LUT4_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27361\,
            lcout => \ALU.madd_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_398_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__27328\,
            in2 => \N__27316\,
            in3 => \N__27307\,
            lcout => \ALU.madd_398_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJJH11_0_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27629\,
            in1 => \N__27680\,
            in2 => \_gnd_net_\,
            in3 => \N__30978\,
            lcout => \ALU.r4_RNIJJH11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIBROO_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30979\,
            in1 => \N__34854\,
            in2 => \_gnd_net_\,
            in3 => \N__34941\,
            lcout => OPEN,
            ltout => \ALU.r0_RNIBROOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIVVDO2_0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__27763\,
            in1 => \N__30928\,
            in2 => \N__27757\,
            in3 => \N__27720\,
            lcout => \ALU.a_7_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__34942\,
            in1 => \N__30067\,
            in2 => \N__30416\,
            in3 => \N__39438\,
            lcout => OPEN,
            ltout => \TXbuffer_18_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__27681\,
            in1 => \N__30079\,
            in2 => \N__27658\,
            in3 => \N__34065\,
            lcout => \TXbuffer_RNO_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__30066\,
            in2 => \N__30415\,
            in3 => \N__30656\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30068\,
            in1 => \N__33717\,
            in2 => \N__27640\,
            in3 => \N__27630\,
            lcout => \TXbuffer_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_1_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30060\,
            in1 => \N__27785\,
            in2 => \N__27559\,
            in3 => \N__29429\,
            lcout => \TXbuffer_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_4_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__27589\,
            in1 => \N__30371\,
            in2 => \N__30081\,
            in3 => \N__28701\,
            lcout => \TXbuffer_18_13_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__30061\,
            in1 => \N__31010\,
            in2 => \N__30397\,
            in3 => \N__32959\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30058\,
            in1 => \N__33691\,
            in2 => \N__28000\,
            in3 => \N__33664\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110010001"
        )
    port map (
            in0 => \N__27997\,
            in1 => \N__49970\,
            in2 => \N__27982\,
            in3 => \N__27979\,
            lcout => \TXbufferZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56261\,
            ce => \N__56048\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__30054\,
            in1 => \N__27972\,
            in2 => \N__30396\,
            in3 => \N__33388\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30059\,
            in1 => \N__27936\,
            in2 => \N__27898\,
            in3 => \N__33634\,
            lcout => \TXbuffer_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r7_6_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38874\,
            lcout => r7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_7_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38740\,
            lcout => r7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_8_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39524\,
            lcout => r7_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_9_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r7_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42147\,
            lcout => r7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40287\,
            lcout => r7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_3_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50188\,
            lcout => r7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r7_4_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39083\,
            lcout => r7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56266\,
            ce => \N__45888\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s0_c_RNO_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33010\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \ALU.r0_12_prm_8_10_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s0_c_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42342\,
            in2 => \N__41998\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_10_s0_cy\,
            carryout => \ALU.r0_12_prm_8_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_10_s0_c_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34513\,
            in2 => \N__51562\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_10_s0\,
            carryout => \ALU.r0_12_prm_7_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_10_s0_c_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34737\,
            in2 => \N__35257\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_10_s0\,
            carryout => \ALU.r0_12_prm_6_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_10_s0_c_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34698\,
            in2 => \N__45565\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_10_s0\,
            carryout => \ALU.r0_12_prm_5_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_10_s0_c_inv_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34665\,
            in2 => \N__34612\,
            in3 => \N__51794\,
            lcout => \ALU.a_i_10\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_10_s0\,
            carryout => \ALU.r0_12_prm_4_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_10_s0_c_inv_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55167\,
            in1 => \N__28213\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_10_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_10_s0\,
            carryout => \ALU.r0_12_prm_3_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_10_s0_c_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35641\,
            in2 => \N__35857\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_10_s0\,
            carryout => \ALU.r0_12_prm_2_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_10_s0_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36109\,
            in2 => \N__34201\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \ALU.r0_12_s0_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_10_s0_c_RNI4UV4363_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28207\,
            in1 => \N__34639\,
            in2 => \_gnd_net_\,
            in3 => \N__28195\,
            lcout => \ALU.r0_12_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_10_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28158\,
            lcout => r0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56274\,
            ce => \N__49719\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s0_c_RNO_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46525\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \ALU.r0_12_prm_8_14_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s0_c_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47980\,
            in2 => \N__39634\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_14_s0_cy\,
            carryout => \ALU.r0_12_prm_8_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_14_s0_c_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47928\,
            in2 => \N__42955\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_14_s0\,
            carryout => \ALU.r0_12_prm_7_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_14_s0_c_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47895\,
            in2 => \N__39646\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_14_s0\,
            carryout => \ALU.r0_12_prm_6_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_14_s0_c_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39667\,
            in2 => \N__47866\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_14_s0\,
            carryout => \ALU.r0_12_prm_5_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_14_s0_c_inv_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47823\,
            in2 => \N__39685\,
            in3 => \N__46959\,
            lcout => \ALU.a_i_14\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_14_s0\,
            carryout => \ALU.r0_12_prm_4_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_14_s0_c_inv_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55168\,
            in1 => \_gnd_net_\,
            in2 => \N__28336\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_14_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_14_s0\,
            carryout => \ALU.r0_12_prm_3_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_14_s0_c_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49140\,
            in2 => \N__36052\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_14_s0\,
            carryout => \ALU.r0_12_prm_2_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_14_s0_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49083\,
            in2 => \N__31216\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \ALU.r0_12_s0_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_14_s0_c_RNI357RUG3_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28327\,
            in1 => \N__49033\,
            in2 => \_gnd_net_\,
            in3 => \N__28315\,
            lcout => \ALU.r0_12_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_14_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28293\,
            lcout => r1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56284\,
            ce => \N__47569\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s0_c_RNO_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35656\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \ALU.r0_12_prm_8_12_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s0_c_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37468\,
            in2 => \N__34480\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_12_s0_cy\,
            carryout => \ALU.r0_12_prm_8_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_12_s0_c_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37437\,
            in2 => \N__31285\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_12_s0\,
            carryout => \ALU.r0_12_prm_7_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_12_s0_c_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37410\,
            in2 => \N__31270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_12_s0\,
            carryout => \ALU.r0_12_prm_6_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_12_s0_c_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37369\,
            in2 => \N__31318\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_12_s0\,
            carryout => \ALU.r0_12_prm_5_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_12_s0_c_inv_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37323\,
            in2 => \N__36175\,
            in3 => \N__41350\,
            lcout => \ALU.a_i_12\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_12_s0\,
            carryout => \ALU.r0_12_prm_4_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_12_s0_c_inv_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55166\,
            in1 => \N__28465\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_12_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_12_s0\,
            carryout => \ALU.r0_12_prm_3_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_12_s0_c_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37654\,
            in2 => \N__35695\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_12_s0\,
            carryout => \ALU.r0_12_prm_2_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_12_s0_c_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37594\,
            in2 => \N__36064\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \ALU.r0_12_s0_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_12_s0_c_RNIS2VGA6_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37552\,
            in1 => \N__28459\,
            in2 => \_gnd_net_\,
            in3 => \N__28450\,
            lcout => \ALU.r0_12_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28402\,
            lcout => r0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56291\,
            ce => \N__49718\,
            sr => \_gnd_net_\
        );

    \TXbuffer_5_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__28510\,
            in1 => \N__28501\,
            in2 => \N__49967\,
            in3 => \N__28492\,
            lcout => \TXbufferZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56295\,
            ce => \N__56039\,
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_1_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__32548\,
            in1 => \N__32692\,
            in2 => \N__32277\,
            in3 => \N__46797\,
            lcout => \ALU.a2_b_1\,
            ltout => \ALU.a2_b_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_8_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__28480\,
            in1 => \N__49353\,
            in2 => \N__28483\,
            in3 => \N__37994\,
            lcout => \ALU.madd_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a1_b_2_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__31666\,
            in1 => \N__31719\,
            in2 => \N__32276\,
            in3 => \N__43931\,
            lcout => \ALU.a1_b_2\,
            ltout => \ALU.a1_b_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_4_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__28474\,
            in1 => \N__49352\,
            in2 => \N__28468\,
            in3 => \N__37993\,
            lcout => \ALU.madd_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_3_c_RNO_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__44359\,
            in1 => \N__53951\,
            in2 => \N__53216\,
            in3 => \N__49360\,
            lcout => \ALU.r0_12_prm_6_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a2_b_0_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__32691\,
            in1 => \N__32549\,
            in2 => \N__32236\,
            in3 => \N__37992\,
            lcout => \ALU.a2_b_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_2_c_RNO_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54553\,
            in1 => \N__48402\,
            in2 => \N__53217\,
            in3 => \N__43932\,
            lcout => \ALU.r0_12_prm_5_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIL9636_2_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__48403\,
            in1 => \N__53090\,
            in2 => \N__54047\,
            in3 => \N__54554\,
            lcout => \ALU.r4_RNIL9636Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_39_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28621\,
            in1 => \N__28606\,
            in2 => \N__29563\,
            in3 => \N__28597\,
            lcout => \ALU.madd_39\,
            ltout => \ALU.madd_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_45_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__31591\,
            in1 => \N__28918\,
            in2 => \N__28582\,
            in3 => \N__28537\,
            lcout => \ALU.madd_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI97EK9_5_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__53949\,
            in1 => \N__45360\,
            in2 => \N__54787\,
            in3 => \N__43365\,
            lcout => \ALU.lshift_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_23_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__31590\,
            in1 => \N__28917\,
            in2 => \_gnd_net_\,
            in3 => \N__28536\,
            lcout => OPEN,
            ltout => \ALU.madd_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_4_l_fx_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28579\,
            in2 => \N__28573\,
            in3 => \N__28570\,
            lcout => \ALU.madd_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_19_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31589\,
            in1 => \N__28916\,
            in2 => \_gnd_net_\,
            in3 => \N__28535\,
            lcout => \ALU.madd_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIM8HG5_5_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__53950\,
            in1 => \N__53159\,
            in2 => \N__54788\,
            in3 => \N__45361\,
            lcout => \ALU.r4_RNIM8HG5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_1_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__41942\,
            in1 => \N__48955\,
            in2 => \N__29319\,
            in3 => \N__43947\,
            lcout => \ALU.madd_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_0_s1_c_RNO_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__48944\,
            in1 => \N__38028\,
            in2 => \_gnd_net_\,
            in3 => \N__55230\,
            lcout => \ALU.r0_12_prm_3_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_66_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28893\,
            in2 => \_gnd_net_\,
            in3 => \N__28868\,
            lcout => \ALU.madd_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKO1J4_5_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29237\,
            in1 => \N__29076\,
            in2 => \_gnd_net_\,
            in3 => \N__29004\,
            lcout => \ALU.a_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_4_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48943\,
            in2 => \_gnd_net_\,
            in3 => \N__40523\,
            lcout => \ALU.a0_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIUM9JC_2_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33936\,
            in2 => \_gnd_net_\,
            in3 => \N__28906\,
            lcout => \ALU.r4_RNIUM9JCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_6_ma_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28894\,
            in2 => \_gnd_net_\,
            in3 => \N__28869\,
            lcout => \ALU.madd_cry_6_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_0_s0_c_RNO_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100010001"
        )
    port map (
            in0 => \N__48945\,
            in1 => \N__38029\,
            in2 => \N__53213\,
            in3 => \N__53804\,
            lcout => \ALU.r0_12_prm_6_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI18BO_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28840\,
            in1 => \N__28724\,
            in2 => \_gnd_net_\,
            in3 => \N__28798\,
            lcout => \ALU.r2_RNI18BOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_0_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34987\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56245\,
            ce => \N__47671\,
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI4H0S_1_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28705\,
            in1 => \N__28663\,
            in2 => \_gnd_net_\,
            in3 => \N__29518\,
            lcout => \ALU.r2_RNI4H0SZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_RNIC9P41_1_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29517\,
            in1 => \N__29440\,
            in2 => \_gnd_net_\,
            in3 => \N__29407\,
            lcout => \ALU.r6_RNIC9P41Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIDAOQ3_2_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__33340\,
            in1 => \N__32862\,
            in2 => \_gnd_net_\,
            in3 => \N__29365\,
            lcout => \ALU.b_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIHU8AD1_15_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37498\,
            in1 => \N__51509\,
            in2 => \_gnd_net_\,
            in3 => \N__31333\,
            lcout => \ALU.rshift_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_3_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__44335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48998\,
            lcout => \ALU.a0_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNID26E8_0_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__48999\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37988\,
            lcout => \ALU.un14_log_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_13_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__29290\,
            in1 => \_gnd_net_\,
            in2 => \N__29299\,
            in3 => \N__29275\,
            lcout => \ALU.madd_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_3_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010100000"
        )
    port map (
            in0 => \N__41951\,
            in1 => \N__48983\,
            in2 => \N__29320\,
            in3 => \N__43916\,
            lcout => \ALU.madd_3\,
            ltout => \ALU.madd_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_axb_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29289\,
            in1 => \_gnd_net_\,
            in2 => \N__29278\,
            in3 => \N__29274\,
            lcout => \ALU.madd_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI7AQC9_15_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40175\,
            in2 => \_gnd_net_\,
            in3 => \N__40009\,
            lcout => \ALU.un14_log_0_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_1_c_RNO_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53098\,
            in2 => \_gnd_net_\,
            in3 => \N__41952\,
            lcout => \ALU.r0_12_prm_7_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_2_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__31934\,
            in1 => \N__31829\,
            in2 => \N__32272\,
            in3 => \N__43915\,
            lcout => \ALU.a3_b_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIRCFPA_0_7_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__53742\,
            in1 => \N__46151\,
            in2 => \N__54697\,
            in3 => \N__44552\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI67NNK_10_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__54520\,
            in1 => \N__52151\,
            in2 => \N__29539\,
            in3 => \N__51805\,
            lcout => \ALU.r5_RNI67NNKZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_2_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40274\,
            lcout => r1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56250\,
            ce => \N__47581\,
            sr => \_gnd_net_\
        );

    \ALU.r1_3_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50171\,
            lcout => r1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56250\,
            ce => \N__47581\,
            sr => \_gnd_net_\
        );

    \ALU.r1_4_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39052\,
            lcout => r1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56250\,
            ce => \N__47581\,
            sr => \_gnd_net_\
        );

    \ALU.r1_1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42129\,
            lcout => r1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56250\,
            ce => \N__47581\,
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIJEMP_7_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__36917\,
            in1 => \N__30740\,
            in2 => \N__33304\,
            in3 => \N__33184\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI82OE1_7_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__33744\,
            in1 => \N__34089\,
            in2 => \N__29536\,
            in3 => \N__33138\,
            lcout => \ALU.r4_RNI82OE1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_7_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38727\,
            lcout => r0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56254\,
            ce => \N__49756\,
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_3_7_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__30084\,
            in1 => \N__30487\,
            in2 => \N__30418\,
            in3 => \N__36918\,
            lcout => OPEN,
            ltout => \TXbuffer_18_10_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_7_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30083\,
            in1 => \N__30451\,
            in2 => \N__30421\,
            in3 => \N__33745\,
            lcout => \TXbuffer_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_7_7_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__30741\,
            in1 => \N__30082\,
            in2 => \N__30417\,
            in3 => \N__30118\,
            lcout => OPEN,
            ltout => \TXbuffer_18_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_5_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__34090\,
            in1 => \N__30085\,
            in2 => \N__29728\,
            in3 => \N__29725\,
            lcout => OPEN,
            ltout => \TXbuffer_RNO_5Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_2_7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__29683\,
            in1 => \N__49940\,
            in2 => \N__29587\,
            in3 => \N__29584\,
            lcout => \TXbuffer_18_15_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI5IT71_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30971\,
            in1 => \N__32955\,
            in2 => \N__31095\,
            in3 => \N__35082\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIDI992_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30571\,
            in1 => \N__33653\,
            in2 => \N__29566\,
            in3 => \N__34361\,
            lcout => \ALU.r4_RNIDI992Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_fast_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \a_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56255\,
            ce => \N__56050\,
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIHUT71_7_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__30751\,
            in1 => \N__31086\,
            in2 => \N__36922\,
            in3 => \N__30973\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI6BA92_7_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__30936\,
            in1 => \N__34083\,
            in2 => \N__30727\,
            in3 => \N__33738\,
            lcout => \ALU.r4_RNI6BA92Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIJ0U71_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__39431\,
            in1 => \N__31088\,
            in2 => \N__30664\,
            in3 => \N__30972\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIAFA92_8_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__30937\,
            in1 => \N__34055\,
            in2 => \N__30625\,
            in3 => \N__33716\,
            lcout => \ALU.r4_RNIAFA92Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI9MT71_3_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__35049\,
            in1 => \N__31087\,
            in2 => \N__33237\,
            in3 => \N__30970\,
            lcout => \ALU.a_3_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI7KT71_2_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__33407\,
            in1 => \N__31068\,
            in2 => \N__33384\,
            in3 => \N__30975\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIHM992_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__33627\,
            in1 => \N__34325\,
            in2 => \N__30574\,
            in3 => \N__30569\,
            lcout => \ALU.r4_RNIHM992Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40288\,
            lcout => r0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56256\,
            ce => \N__49731\,
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIBOT71_4_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__30977\,
            in1 => \N__33467\,
            in2 => \N__31085\,
            in3 => \N__33497\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIQU992_4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__30930\,
            in1 => \N__33561\,
            in2 => \N__31099\,
            in3 => \N__34290\,
            lcout => \ALU.r4_RNIQU992Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_4_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39078\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56256\,
            ce => \N__49731\,
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIL2U71_9_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__31134\,
            in1 => \N__31067\,
            in2 => \N__31012\,
            in3 => \N__30976\,
            lcout => OPEN,
            ltout => \ALU.a_3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIEJA92_9_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__34391\,
            in1 => \N__30929\,
            in2 => \N__30817\,
            in3 => \N__33680\,
            lcout => \ALU.r4_RNIEJA92Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s0_c_RNO_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43033\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \ALU.r0_12_prm_8_9_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s0_c_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42586\,
            in2 => \N__36853\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_9_s0_cy\,
            carryout => \ALU.r0_12_prm_8_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_9_s0_c_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42541\,
            in2 => \N__45910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_9_s0\,
            carryout => \ALU.r0_12_prm_7_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_9_s0_c_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45544\,
            in2 => \N__30769\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_9_s0\,
            carryout => \ALU.r0_12_prm_6_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_9_s0_c_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42507\,
            in2 => \N__42037\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_9_s0\,
            carryout => \ALU.r0_12_prm_5_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_9_s0_c_inv_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__52302\,
            in1 => \N__42468\,
            in2 => \N__48100\,
            in3 => \_gnd_net_\,
            lcout => \ALU.a_i_9\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_9_s0\,
            carryout => \ALU.r0_12_prm_4_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_9_s0_c_inv_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31186\,
            in2 => \_gnd_net_\,
            in3 => \N__55262\,
            lcout => \ALU.r0_12_prm_3_9_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_9_s0\,
            carryout => \ALU.r0_12_prm_3_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_9_s0_c_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42430\,
            in2 => \N__31180\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_9_s0\,
            carryout => \ALU.r0_12_prm_2_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_9_s0_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42399\,
            in2 => \N__35677\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \ALU.r0_12_s0_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_9_s0_c_RNI39QBSO_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31162\,
            in1 => \N__42970\,
            in2 => \_gnd_net_\,
            in3 => \N__31150\,
            lcout => \ALU.r0_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_9_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34015\,
            lcout => r0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56262\,
            ce => \N__49732\,
            sr => \_gnd_net_\
        );

    \ALU.r4_RNISU5D9_1_9_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__52309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47476\,
            lcout => \ALU.r4_RNISU5D9_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s1_c_RNO_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55528\,
            in2 => \_gnd_net_\,
            in3 => \N__34424\,
            lcout => \ALU.r0_12_prm_8_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIA5SI9_12_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__53753\,
            in1 => \N__41293\,
            in2 => \N__54557\,
            in3 => \N__40981\,
            lcout => \ALU.rshift_10_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_5_s0_c_RNO_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100100000011"
        )
    port map (
            in0 => \N__53856\,
            in1 => \N__45453\,
            in2 => \N__45262\,
            in3 => \N__53196\,
            lcout => \ALU.r0_12_prm_6_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_12_s0_c_RNO_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__39861\,
            in1 => \N__53857\,
            in2 => \N__53243\,
            in3 => \N__41294\,
            lcout => \ALU.r0_12_prm_6_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIUF9K8_0_10_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__51827\,
            in1 => \_gnd_net_\,
            in2 => \N__52035\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r5_RNIUF9K8_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_10_s1_c_RNO_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53195\,
            in1 => \N__52024\,
            in2 => \_gnd_net_\,
            in3 => \N__51826\,
            lcout => \ALU.r0_12_prm_7_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_15_s1_c_RNO_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__36248\,
            in1 => \N__55927\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_2_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_13_s0_c_RNO_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55950\,
            in2 => \_gnd_net_\,
            in3 => \N__34589\,
            lcout => \ALU.r0_12_prm_2_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_14_s0_c_RNO_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55951\,
            in1 => \N__53758\,
            in2 => \_gnd_net_\,
            in3 => \N__49073\,
            lcout => \ALU.r0_12_prm_1_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIUF9K8_10_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52028\,
            in2 => \_gnd_net_\,
            in3 => \N__51831\,
            lcout => \ALU.un14_log_0_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s1_c_RNO_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__55529\,
            in1 => \N__36014\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_8_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNISMSV4_15_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__54603\,
            in1 => \N__53757\,
            in2 => \_gnd_net_\,
            in3 => \N__40097\,
            lcout => \ALU.r5_RNISMSV4Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI465TI_13_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__31342\,
            in1 => \N__46988\,
            in2 => \N__54777\,
            in3 => \N__41556\,
            lcout => \ALU.r5_RNI465TIZ0Z_13\,
            ltout => \ALU.r5_RNI465TIZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIOL1S71_10_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51033\,
            in2 => \N__31336\,
            in3 => \N__32917\,
            lcout => \ALU.r5_RNIOL1S71Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNID2JJ9_13_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35428\,
            in2 => \_gnd_net_\,
            in3 => \N__41557\,
            lcout => \ALU.un14_log_0_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_15_s0_c_RNO_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53759\,
            in1 => \N__40160\,
            in2 => \N__53241\,
            in3 => \N__39992\,
            lcout => \ALU.r0_12_prm_6_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_12_s0_c_RNO_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111000011"
        )
    port map (
            in0 => \N__54582\,
            in1 => \N__39874\,
            in2 => \N__41368\,
            in3 => \N__53194\,
            lcout => \ALU.r0_12_prm_5_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_10_s1_c_RNO_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__51832\,
            in1 => \N__54581\,
            in2 => \N__53242\,
            in3 => \N__52002\,
            lcout => \ALU.r0_12_prm_5_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI7AQC9_1_15_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__39994\,
            in1 => \_gnd_net_\,
            in2 => \N__40174\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r2_RNI7AQC9_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s0_c_RNO_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55527\,
            in2 => \_gnd_net_\,
            in3 => \N__34423\,
            lcout => \ALU.r0_12_prm_8_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_12_s0_c_RNO_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__41358\,
            in1 => \N__39873\,
            in2 => \_gnd_net_\,
            in3 => \N__53193\,
            lcout => \ALU.r0_12_prm_7_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_15_s0_c_RNO_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54606\,
            in1 => \N__40159\,
            in2 => \N__53240\,
            in3 => \N__39993\,
            lcout => \ALU.r0_12_prm_5_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s1_c_RNO_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39889\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \ALU.r0_12_prm_8_13_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s1_c_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36118\,
            in2 => \N__36159\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_13_s1_cy\,
            carryout => \ALU.r0_12_prm_8_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_13_s1_c_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31492\,
            in2 => \N__31477\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_13_s1\,
            carryout => \ALU.r0_12_prm_7_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_13_s1_c_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31444\,
            in2 => \N__31428\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_13_s1\,
            carryout => \ALU.r0_12_prm_6_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_13_s1_c_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31411\,
            in2 => \N__31399\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_13_s1\,
            carryout => \ALU.r0_12_prm_5_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_13_s1_c_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31372\,
            in2 => \N__31360\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_13_s1\,
            carryout => \ALU.r0_12_prm_4_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_13_s1_c_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55263\,
            in2 => \N__56476\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_13_s1\,
            carryout => \ALU.r0_12_prm_3_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_13_s1_c_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34555\,
            in2 => \N__34596\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_13_s1\,
            carryout => \ALU.r0_12_prm_2_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_13_s1_c_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35301\,
            in2 => \N__31504\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \ALU.r0_12_s1_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_13_THRU_LUT4_0_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31516\,
            lcout => \ALU.r0_12_s1_13_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_13_s1_c_RNO_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55957\,
            in1 => \N__53985\,
            in2 => \_gnd_net_\,
            in3 => \N__35300\,
            lcout => \ALU.r0_12_prm_1_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_6_s1_c_RNO_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55840\,
            in2 => \_gnd_net_\,
            in3 => \N__38257\,
            lcout => \ALU.r0_12_prm_2_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_0_s0_c_RNO_LC_10_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__55221\,
            in1 => \N__49002\,
            in2 => \_gnd_net_\,
            in3 => \N__38031\,
            lcout => \ALU.r0_12_prm_3_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_6_s1_c_RNO_LC_10_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53080\,
            in2 => \_gnd_net_\,
            in3 => \N__41629\,
            lcout => \ALU.r0_12_prm_7_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_6_s1_c_RNO_LC_10_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__43656\,
            in1 => \N__54894\,
            in2 => \N__53214\,
            in3 => \N__43416\,
            lcout => \ALU.r0_12_prm_5_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_RNO_4_LC_10_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__54032\,
            in1 => \N__48399\,
            in2 => \N__54920\,
            in3 => \N__49398\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_RNO_3_LC_10_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__54552\,
            in1 => \N__45452\,
            in2 => \N__31495\,
            in3 => \N__42849\,
            lcout => \ALU.r0_12_prm_8_2_c_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a3_b_3_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__31936\,
            in1 => \N__44352\,
            in2 => \N__32229\,
            in3 => \N__31839\,
            lcout => \ALU.a3_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a1_b_1_LC_10_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__31664\,
            in1 => \N__31731\,
            in2 => \N__32228\,
            in3 => \N__46798\,
            lcout => \ALU.a1_b_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a1_b_3_LC_10_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__44351\,
            in1 => \N__32178\,
            in2 => \N__31740\,
            in3 => \N__31665\,
            lcout => \ALU.a1_b_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_135_0_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__40504\,
            in1 => \N__44350\,
            in2 => \N__45418\,
            in3 => \N__43308\,
            lcout => \ALU.madd_135_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_6_s1_c_RNO_LC_10_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54056\,
            in1 => \N__43655\,
            in2 => \N__53215\,
            in3 => \N__43309\,
            lcout => \ALU.r0_12_prm_6_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_4_c_RNO_0_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42818\,
            in2 => \_gnd_net_\,
            in3 => \N__40533\,
            lcout => \ALU.un14_log_0_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIO7CSJ_4_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000011"
        )
    port map (
            in0 => \N__42816\,
            in1 => \N__31540\,
            in2 => \N__54790\,
            in3 => \N__49397\,
            lcout => \ALU.r4_RNIO7CSJZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI9H7SJ_5_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__31531\,
            in1 => \N__45383\,
            in2 => \N__54800\,
            in3 => \N__42817\,
            lcout => \ALU.r4_RNI9H7SJZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI8B628_0_5_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45231\,
            lcout => \ALU.r4_RNI8B628_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_0_s0_c_RNO_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100001111"
        )
    port map (
            in0 => \N__38026\,
            in1 => \_gnd_net_\,
            in2 => \N__53218\,
            in3 => \N__48935\,
            lcout => \ALU.r0_12_prm_7_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIMVMDA_0_1_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__48933\,
            in1 => \N__53782\,
            in2 => \N__54791\,
            in3 => \N__48639\,
            lcout => \ALU.N_622_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_0_s0_c_RNO_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__38027\,
            in1 => \N__54658\,
            in2 => \N__53219\,
            in3 => \N__48936\,
            lcout => \ALU.r0_12_prm_5_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_0_s1_c_RNO_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__48934\,
            in1 => \N__53091\,
            in2 => \_gnd_net_\,
            in3 => \N__38025\,
            lcout => \ALU.r0_12_prm_7_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIUU8UD_3_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31963\,
            in2 => \_gnd_net_\,
            in3 => \N__49324\,
            lcout => \ALU.r4_RNIUU8UDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNINNEH9_0_15_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__54062\,
            in1 => \N__40176\,
            in2 => \N__47070\,
            in3 => \N__54617\,
            lcout => \ALU.N_845_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKUMQ8_1_8_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__46192\,
            in1 => \_gnd_net_\,
            in2 => \N__46446\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r4_RNIKUMQ8_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a8_b_8_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46422\,
            in2 => \_gnd_net_\,
            in3 => \N__46191\,
            lcout => \ALU.a8_b_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_490_5_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__35594\,
            in1 => \N__42844\,
            in2 => \N__45451\,
            in3 => \N__52003\,
            lcout => \ALU.madd_490_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_RNO_4_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__49325\,
            in1 => \N__54616\,
            in2 => \N__42862\,
            in3 => \N__54055\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_RNO_3_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__54618\,
            in1 => \N__45391\,
            in2 => \N__32923\,
            in3 => \N__43415\,
            lcout => OPEN,
            ltout => \ALU.r0_12_prm_8_3_c_RNOZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_RNO_2_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__50995\,
            in1 => \N__51442\,
            in2 => \N__32920\,
            in3 => \N__32910\,
            lcout => \ALU.rshift_15_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s1_c_RNO_1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__38050\,
            in1 => \N__38075\,
            in2 => \N__51527\,
            in3 => \N__50992\,
            lcout => \ALU.r0_12_prm_8_10_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKTVI8_0_4_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010011010"
        )
    port map (
            in0 => \N__40511\,
            in1 => \N__32224\,
            in2 => \N__32374\,
            in3 => \N__32469\,
            lcout => \ALU.un9_addsub_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNITPNQ3_0_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__32861\,
            in1 => \N__32752\,
            in2 => \_gnd_net_\,
            in3 => \N__32718\,
            lcout => \ALU.b_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIHCHO8_0_2_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011110111000"
        )
    port map (
            in0 => \N__32684\,
            in1 => \N__32223\,
            in2 => \N__32592\,
            in3 => \N__43897\,
            lcout => \ALU.un9_addsub_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKTVI8_4_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001010011"
        )
    port map (
            in0 => \N__32468\,
            in1 => \N__32360\,
            in2 => \N__32257\,
            in3 => \N__40512\,
            lcout => OPEN,
            ltout => \ALU.un2_addsub_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI20C8C_4_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31966\,
            in3 => \N__33882\,
            lcout => \ALU.r4_RNI20C8CZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s0_c_RNO_1_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__38051\,
            in1 => \N__38076\,
            in2 => \N__51528\,
            in3 => \N__50993\,
            lcout => \ALU.rshift_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_g0_12_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43898\,
            in1 => \N__44529\,
            in2 => \N__46217\,
            in3 => \N__46822\,
            lcout => \ALU.madd_76_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKUMQ8_8_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46161\,
            in2 => \_gnd_net_\,
            in3 => \N__46412\,
            lcout => \ALU.un14_log_0_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI14AH9_11_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__53911\,
            in1 => \N__51804\,
            in2 => \N__40989\,
            in3 => \N__54835\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI1RK3K_9_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__54836\,
            in1 => \N__46160\,
            in2 => \N__32983\,
            in3 => \N__52255\,
            lcout => \ALU.r4_RNI1RK3KZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIQK1ED_4_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32980\,
            in3 => \N__42838\,
            lcout => \ALU.r4_RNIQK1EDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIVLAIA_9_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46162\,
            in1 => \N__53912\,
            in2 => \_gnd_net_\,
            in3 => \N__52256\,
            lcout => \ALU.r4_RNIVLAIAZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2H9PK_6_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__44588\,
            in1 => \N__32971\,
            in2 => \N__43437\,
            in3 => \N__54837\,
            lcout => \ALU.r4_RNI2H9PKZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_7_s0_c_RNO_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__44797\,
            in1 => \N__53913\,
            in2 => \N__53220\,
            in3 => \N__44589\,
            lcout => \ALU.r0_12_prm_6_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIE5LH_1_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32954\,
            in1 => \N__35069\,
            in2 => \_gnd_net_\,
            in3 => \N__33174\,
            lcout => \ALU.r0_RNIE5LHZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI50MP_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__33204\,
            in1 => \N__33296\,
            in2 => \N__34853\,
            in3 => \N__34932\,
            lcout => \ALU.b_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_fast_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33205\,
            lcout => \b_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56248\,
            ce => \N__56052\,
            sr => \_gnd_net_\
        );

    \ALU.r0_RNID8MP_4_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__33507\,
            in1 => \N__33299\,
            in2 => \N__33468\,
            in3 => \N__33183\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNISLNE1_4_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__33137\,
            in1 => \N__34289\,
            in2 => \N__33442\,
            in3 => \N__33560\,
            lcout => \ALU.r4_RNISLNE1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNI94MP_2_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__33411\,
            in1 => \N__33297\,
            in2 => \N__33380\,
            in3 => \N__33181\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKDNE1_2_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__33135\,
            in1 => \N__34329\,
            in2 => \N__33352\,
            in3 => \N__33626\,
            lcout => \ALU.r4_RNIKDNE1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_RNIB6MP_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__35042\,
            in1 => \N__33298\,
            in2 => \N__33233\,
            in3 => \N__33182\,
            lcout => OPEN,
            ltout => \ALU.b_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIOHNE1_3_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__33136\,
            in1 => \N__33064\,
            in2 => \N__33040\,
            in3 => \N__33585\,
            lcout => \ALU.r4_RNIOHNE1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_6_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38855\,
            lcout => r5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_7_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38741\,
            lcout => r5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_8_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39513\,
            lcout => r5_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_9_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34022\,
            lcout => r5_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_1_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42139\,
            lcout => r5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40275\,
            lcout => r5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50175\,
            lcout => r5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.r5_4_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39062\,
            lcout => r5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => \N__45801\,
            sr => \_gnd_net_\
        );

    \ALU.mult_a0_b_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49008\,
            in2 => \N__40647\,
            in3 => \N__38015\,
            lcout => \ALU.mult_0\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \ALU.un2_addsub_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_0_c_RNIJPSHD_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34489\,
            in2 => \N__33544\,
            in3 => \N__33964\,
            lcout => \ALU.un2_addsub_cry_0_c_RNIJPSHDZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_0\,
            carryout => \ALU.un2_addsub_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_1_c_RNI1H7SG_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33961\,
            in2 => \N__33949\,
            in3 => \N__33925\,
            lcout => \ALU.un2_addsub_cry_1_c_RNI1H7SGZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_1\,
            carryout => \ALU.un2_addsub_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_2_c_RNI3K9SG_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33922\,
            in2 => \N__33910\,
            in3 => \N__33895\,
            lcout => \ALU.un2_addsub_cry_2_c_RNI3K9SGZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_2\,
            carryout => \ALU.un2_addsub_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_3_c_RNI8MVBG_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33892\,
            in2 => \N__33883\,
            in3 => \N__33856\,
            lcout => \ALU.un2_addsub_cry_3_c_RNI8MVBGZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_3\,
            carryout => \ALU.un2_addsub_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_4_c_RNILPG3D_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45479\,
            in2 => \N__33853\,
            in3 => \N__33835\,
            lcout => \ALU.un2_addsub_cry_4_c_RNILPG3DZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_4\,
            carryout => \ALU.un2_addsub_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_5_c_RNIO30SD_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43438\,
            in2 => \N__33832\,
            in3 => \N__33808\,
            lcout => \ALU.un2_addsub_cry_5_c_RNIO30SDZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_5\,
            carryout => \ALU.un2_addsub_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_6_c_RNIPJK8E_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44593\,
            in2 => \N__40666\,
            in3 => \N__33805\,
            lcout => \ALU.un2_addsub_cry_6_c_RNIPJK8EZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_6\,
            carryout => \ALU.un2_addsub_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_7_c_RNI5ELEE_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46177\,
            in2 => \N__33802\,
            in3 => \N__33790\,
            lcout => \ALU.un2_addsub_cry_7_c_RNI5ELEEZ0\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \ALU.un2_addsub_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_8_c_RNINO51F_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52301\,
            in2 => \N__47287\,
            in3 => \N__33787\,
            lcout => \ALU.un2_addsub_cry_8_c_RNINO51FZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_8\,
            carryout => \ALU.un2_addsub_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_9_c_RNIS67KD_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51716\,
            in2 => \N__34189\,
            in3 => \N__34171\,
            lcout => \ALU.un2_addsub_cry_9_c_RNIS67KDZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_9\,
            carryout => \ALU.un2_addsub_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_10_c_RNIS4T7D_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40982\,
            in2 => \N__34168\,
            in3 => \N__34147\,
            lcout => \ALU.un2_addsub_cry_10_c_RNIS4T7DZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_10\,
            carryout => \ALU.un2_addsub_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_11_c_RNICP8AE_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41357\,
            in2 => \N__34144\,
            in3 => \N__34132\,
            lcout => \ALU.un2_addsub_cry_11_c_RNICP8AEZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_11\,
            carryout => \ALU.un2_addsub_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_12_c_RNI74A7E_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41561\,
            in2 => \N__34129\,
            in3 => \N__34111\,
            lcout => \ALU.un2_addsub_cry_12_c_RNI74A7EZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_12\,
            carryout => \ALU.un2_addsub_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_13_c_RNIR5I0E_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47040\,
            in2 => \N__34108\,
            in3 => \N__34096\,
            lcout => \ALU.un2_addsub_cry_13_c_RNIR5I0EZ0\,
            ltout => OPEN,
            carryin => \ALU.un2_addsub_cry_13\,
            carryout => \ALU.un2_addsub_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un2_addsub_cry_14_c_RNIHN1F9_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__40154\,
            in1 => \N__39988\,
            in2 => \_gnd_net_\,
            in3 => \N__34093\,
            lcout => \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_7_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => \N__47787\,
            sr => \_gnd_net_\
        );

    \ALU.r4_8_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39493\,
            lcout => r4_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => \N__47787\,
            sr => \_gnd_net_\
        );

    \ALU.r4_9_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34014\,
            lcout => r4_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => \N__47787\,
            sr => \_gnd_net_\
        );

    \ALU.r4_1_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__42143\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => r4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => \N__47787\,
            sr => \_gnd_net_\
        );

    \ALU.r4_2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40289\,
            lcout => r4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => \N__47787\,
            sr => \_gnd_net_\
        );

    \ALU.r4_4_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39082\,
            lcout => r4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => \N__47787\,
            sr => \_gnd_net_\
        );

    \ALU.r5_RNITS6F71_13_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__51105\,
            in1 => \N__34258\,
            in2 => \N__51531\,
            in3 => \N__34462\,
            lcout => OPEN,
            ltout => \ALU.lshift_15_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI7QTIG2_5_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51507\,
            in1 => \N__50752\,
            in2 => \N__34237\,
            in3 => \N__43011\,
            lcout => \ALU.lshift_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s1_c_RNO_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__51106\,
            in1 => \N__44889\,
            in2 => \N__51532\,
            in3 => \N__44844\,
            lcout => \ALU.r0_12_prm_8_11_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNISP2L9_12_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39860\,
            in2 => \_gnd_net_\,
            in3 => \N__41349\,
            lcout => \ALU.un14_log_0_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_11_s0_c_RNO_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55942\,
            in2 => \_gnd_net_\,
            in3 => \N__35833\,
            lcout => \ALU.r0_12_prm_2_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_10_s0_c_RNO_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010101111"
        )
    port map (
            in0 => \N__53999\,
            in1 => \_gnd_net_\,
            in2 => \N__55961\,
            in3 => \N__36101\,
            lcout => \ALU.r0_12_prm_1_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_N_884_i_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.N_884_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIAP7U9_10_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53998\,
            in1 => \N__51825\,
            in2 => \_gnd_net_\,
            in3 => \N__52300\,
            lcout => \ALU.r5_RNIAP7U9Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s0_c_RNO_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101001011"
        )
    port map (
            in0 => \N__51473\,
            in1 => \N__37486\,
            in2 => \N__55536\,
            in3 => \N__41029\,
            lcout => \ALU.r0_12_prm_8_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI89OPA_2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__53973\,
            in1 => \N__48408\,
            in2 => \N__54781\,
            in3 => \N__49419\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNII2A0L_1_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__54580\,
            in1 => \N__49017\,
            in2 => \N__34465\,
            in3 => \N__48655\,
            lcout => \ALU.r4_RNII2A0LZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIOK1781_9_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51100\,
            in1 => \N__34461\,
            in2 => \_gnd_net_\,
            in3 => \N__43010\,
            lcout => OPEN,
            ltout => \ALU.r4_RNIOK1781Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI79MLT1_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__51472\,
            in1 => \N__51101\,
            in2 => \N__34447\,
            in3 => \N__50740\,
            lcout => \ALU.lshift_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s0_c_RNO_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55523\,
            in2 => \_gnd_net_\,
            in3 => \N__36013\,
            lcout => \ALU.r0_12_prm_8_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_10_s1_c_RNO_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__51829\,
            in1 => \N__54583\,
            in2 => \N__54048\,
            in3 => \N__52992\,
            lcout => \ALU.r0_12_prm_4_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI27VE5_10_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__53976\,
            in1 => \N__54605\,
            in2 => \N__53165\,
            in3 => \N__51830\,
            lcout => \ALU.r5_RNI27VE5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_13_s1_c_RNO_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55920\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34579\,
            lcout => \ALU.r0_12_prm_2_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_10_s1_c_RNO_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55919\,
            in2 => \_gnd_net_\,
            in3 => \N__35636\,
            lcout => \ALU.r0_12_prm_2_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_10_s1_c_RNO_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53975\,
            in1 => \N__52001\,
            in2 => \N__53164\,
            in3 => \N__51828\,
            lcout => \ALU.r0_12_prm_6_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s0_c_RNO_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__54604\,
            in1 => \N__53974\,
            in2 => \N__50707\,
            in3 => \N__40155\,
            lcout => \ALU.rshift_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_11_s0_c_RNO_1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__51104\,
            in1 => \N__44888\,
            in2 => \N__51541\,
            in3 => \N__44843\,
            lcout => \ALU.rshift_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s1_c_RNO_0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34534\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \ALU.r0_12_prm_8_10_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s1_c_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42256\,
            in2 => \N__42346\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_10_s1_cy\,
            carryout => \ALU.r0_12_prm_8_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_10_s1_c_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34522\,
            in2 => \N__34512\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_10_s1\,
            carryout => \ALU.r0_12_prm_7_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_10_s1_c_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34744\,
            in2 => \N__34738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_10_s1\,
            carryout => \ALU.r0_12_prm_6_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_10_s1_c_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34711\,
            in2 => \N__34705\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_10_s1\,
            carryout => \ALU.r0_12_prm_5_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_10_s1_c_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34681\,
            in2 => \N__34675\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_10_s1\,
            carryout => \ALU.r0_12_prm_4_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_10_s1_c_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55264\,
            in2 => \N__56477\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_10_s1\,
            carryout => \ALU.r0_12_prm_3_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_10_s1_c_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35637\,
            in2 => \N__34651\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_10_s1\,
            carryout => \ALU.r0_12_prm_2_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_10_s1_c_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36108\,
            in2 => \N__36073\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \ALU.r0_12_s1_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_10_THRU_LUT4_0_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34642\,
            lcout => \ALU.r0_12_s1_10_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_13_s0_c_RNO_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55958\,
            in1 => \N__53986\,
            in2 => \_gnd_net_\,
            in3 => \N__35296\,
            lcout => \ALU.r0_12_prm_1_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_6_s1_c_THRU_CRY_0_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37726\,
            in2 => \N__37734\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_1_0_\,
            carryout => \ALU.r0_12_prm_8_6_s1_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_6_s1_c_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34819\,
            in2 => \N__37689\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_6_s1_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_6_s1_c_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41642\,
            in2 => \N__34789\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_6_s1\,
            carryout => \ALU.r0_12_prm_7_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_6_s1_c_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34780\,
            in2 => \N__38361\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_6_s1\,
            carryout => \ALU.r0_12_prm_6_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_6_s1_c_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34774\,
            in2 => \N__38340\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_6_s1\,
            carryout => \ALU.r0_12_prm_5_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_6_s1_c_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34765\,
            in2 => \N__38296\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_6_s1\,
            carryout => \ALU.r0_12_prm_4_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_6_s1_c_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55222\,
            in2 => \N__56512\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_6_s1\,
            carryout => \ALU.r0_12_prm_3_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_6_s1_c_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38266\,
            in2 => \N__34753\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_6_s1\,
            carryout => \ALU.r0_12_prm_2_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_6_s1_c_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38204\,
            in2 => \N__36358\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \ALU.r0_12_s1_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_6_THRU_LUT4_0_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34825\,
            lcout => \ALU.r0_12_s1_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIAP9541_4_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__50994\,
            in1 => \N__42222\,
            in2 => \N__51483\,
            in3 => \N__42205\,
            lcout => \ALU.lshift_6\,
            ltout => \ALU.lshift_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_6_s1_c_RNO_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34822\,
            in3 => \N__55458\,
            lcout => \ALU.r0_12_prm_8_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2BKQ8_0_6_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43657\,
            in2 => \_gnd_net_\,
            in3 => \N__43403\,
            lcout => \ALU.r4_RNI2BKQ8_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIUGHG5_6_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__43404\,
            in1 => \N__54783\,
            in2 => \N__53152\,
            in3 => \N__54036\,
            lcout => \ALU.r4_RNIUGHG5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI5OTIG2_2_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__36376\,
            in1 => \N__41098\,
            in2 => \N__51484\,
            in3 => \N__41707\,
            lcout => \ALU.rshift_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNID26E8_1_0_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49001\,
            in2 => \_gnd_net_\,
            in3 => \N__38016\,
            lcout => \ALU.un9_addsub_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_0_s0_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40704\,
            in2 => \N__40198\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \ALU.r0_12_prm_8_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_0_s0_c_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36439\,
            in2 => \N__34813\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_0_s0\,
            carryout => \ALU.r0_12_prm_7_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_0_s0_c_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36312\,
            in2 => \N__34801\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_0_s0\,
            carryout => \ALU.r0_12_prm_6_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_0_s0_c_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37756\,
            in2 => \N__34921\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_0_s0\,
            carryout => \ALU.r0_12_prm_5_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_0_s0_c_inv_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36279\,
            in2 => \N__34912\,
            in3 => \N__48909\,
            lcout => \ALU.N_883_i\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_0_s0\,
            carryout => \ALU.r0_12_prm_4_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_0_s0_c_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36440\,
            in2 => \N__34894\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_0_s0\,
            carryout => \ALU.r0_12_prm_3_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_0_s0_c_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40617\,
            in2 => \N__36367\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_0_s0\,
            carryout => \ALU.r0_12_prm_2_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_0_s0_c_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36399\,
            in2 => \N__34882\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_2_0_s0\,
            carryout => \ALU.r0_12_s0_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_0_s0_c_RNIGKQLG2_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36382\,
            in1 => \N__34867\,
            in2 => \_gnd_net_\,
            in3 => \N__34858\,
            lcout => \ALU.r0_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_0_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34970\,
            lcout => r1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56234\,
            ce => \N__47576\,
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIRCFPA_7_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__53872\,
            in1 => \N__46199\,
            in2 => \N__54888\,
            in3 => \N__44530\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIODO6K_5_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__43379\,
            in1 => \N__54821\,
            in2 => \N__35101\,
            in3 => \N__45484\,
            lcout => \ALU.r4_RNIODO6KZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNILIPV9_6_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53873\,
            in1 => \N__43380\,
            in2 => \_gnd_net_\,
            in3 => \N__44531\,
            lcout => OPEN,
            ltout => \ALU.r4_RNILIPV9Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI1G9PK_6_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54822\,
            in2 => \N__35098\,
            in3 => \N__38631\,
            lcout => \ALU.r4_RNI1G9PKZ0Z_6\,
            ltout => \ALU.r4_RNI1G9PKZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNICUATH1_15_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__36835\,
            in1 => \N__51423\,
            in2 => \N__35095\,
            in3 => \N__38052\,
            lcout => \ALU.rshift_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJTDS9_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__53871\,
            in1 => \N__45483\,
            in2 => \N__54887\,
            in3 => \N__42837\,
            lcout => \ALU.lshift_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_5_s0_c_RNO_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55941\,
            in2 => \_gnd_net_\,
            in3 => \N__45686\,
            lcout => \ALU.r0_12_prm_2_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI8R2TI_11_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54817\,
            in1 => \N__38649\,
            in2 => \_gnd_net_\,
            in3 => \N__41728\,
            lcout => \ALU.r5_RNI8R2TIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42154\,
            lcout => r0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56240\,
            ce => \N__49685\,
            sr => \_gnd_net_\
        );

    \ALU.r0_3_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50136\,
            lcout => r0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56240\,
            ce => \N__49685\,
            sr => \_gnd_net_\
        );

    \ALU.r0_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34986\,
            lcout => r0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56240\,
            ce => \N__49685\,
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI9S2TI_11_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__35665\,
            in1 => \N__51815\,
            in2 => \N__54638\,
            in3 => \N__40991\,
            lcout => OPEN,
            ltout => \ALU.r5_RNI9S2TIZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI8VM481_11_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__51474\,
            in1 => \N__51047\,
            in2 => \N__35164\,
            in3 => \N__36867\,
            lcout => OPEN,
            ltout => \ALU.lshift_15_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIS8K872_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51475\,
            in1 => \N__46493\,
            in2 => \N__35161\,
            in3 => \N__44827\,
            lcout => \ALU.lshift_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIKS4A9_11_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40990\,
            in1 => \_gnd_net_\,
            in2 => \N__51838\,
            in3 => \N__53644\,
            lcout => \ALU.r5_RNIKS4A9Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI468UD_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35158\,
            in2 => \_gnd_net_\,
            in3 => \N__48395\,
            lcout => \ALU.r4_RNI468UDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_7_s0_c_RNO_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55808\,
            in1 => \N__53646\,
            in2 => \_gnd_net_\,
            in3 => \N__45001\,
            lcout => \ALU.r0_12_prm_1_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_6_s0_c_RNO_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__53645\,
            in1 => \N__55807\,
            in2 => \_gnd_net_\,
            in3 => \N__38185\,
            lcout => \ALU.r0_12_prm_1_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIE0AK8_11_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__40992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35605\,
            lcout => \ALU.un14_log_0_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a6_b_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37960\,
            in2 => \N__49018\,
            in3 => \N__43377\,
            lcout => \ALU.a6_b_0\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \ALU.un9_addsub_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_0_c_RNIG8GLJ_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48638\,
            in2 => \N__35239\,
            in3 => \N__35221\,
            lcout => \ALU.un9_addsub_cry_0_c_RNIG8GLJZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_0\,
            carryout => \ALU.un9_addsub_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_1_c_RNIKO6AJ_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35218\,
            in2 => \N__48409\,
            in3 => \N__35212\,
            lcout => \ALU.un9_addsub_cry_1_c_RNIKO6AJZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_1\,
            carryout => \ALU.un9_addsub_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_2_c_RNIOR8AJ_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49424\,
            in2 => \N__35209\,
            in3 => \N__35194\,
            lcout => \ALU.un9_addsub_cry_2_c_RNIOR8AJZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_2\,
            carryout => \ALU.un9_addsub_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_3_c_RNIV8DFI_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35191\,
            in2 => \N__42868\,
            in3 => \N__35182\,
            lcout => \ALU.un9_addsub_cry_3_c_RNIV8DFIZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_3\,
            carryout => \ALU.un9_addsub_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_4_c_RNI8AH88_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45250\,
            in2 => \N__45514\,
            in3 => \N__35179\,
            lcout => \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_4\,
            carryout => \ALU.un9_addsub_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_5_c_RNI3C019_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43378\,
            in2 => \N__43667\,
            in3 => \N__35176\,
            lcout => \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_5\,
            carryout => \ALU.un9_addsub_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_6_c_RNIJH4R8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44594\,
            in2 => \N__44806\,
            in3 => \N__35173\,
            lcout => \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_6\,
            carryout => \ALU.un9_addsub_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_7_c_RNIN3519_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46200\,
            in2 => \N__46461\,
            in3 => \N__35170\,
            lcout => \ALU.un9_addsub_cry_7_c_RNINZ0Z3519\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \ALU.un9_addsub_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_8_c_RNI06LJ9_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52293\,
            in2 => \N__47475\,
            in3 => \N__35167\,
            lcout => \ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_8\,
            carryout => \ALU.un9_addsub_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_9_c_RNI3PPQ8_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51795\,
            in2 => \N__52029\,
            in3 => \N__35608\,
            lcout => \ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_9\,
            carryout => \ALU.un9_addsub_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_10_c_RNIRLO09_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40911\,
            in2 => \N__35604\,
            in3 => \N__35434\,
            lcout => \ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_10\,
            carryout => \ALU.un9_addsub_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_11_c_RNIAHI1A_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41356\,
            in2 => \N__39875\,
            in3 => \N__35431\,
            lcout => \ALU.un9_addsub_cry_11_c_RNIAHI1AZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_11\,
            carryout => \ALU.un9_addsub_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_12_c_RNISR30A_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41571\,
            in2 => \N__35424\,
            in3 => \N__35266\,
            lcout => \ALU.un9_addsub_cry_12_c_RNISR30AZ0\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_12\,
            carryout => \ALU.un9_addsub_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_13_c_RNI7LBP9_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47056\,
            in2 => \N__47182\,
            in3 => \N__35263\,
            lcout => \ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9\,
            ltout => OPEN,
            carryin => \ALU.un9_addsub_cry_13\,
            carryout => \ALU.un9_addsub_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un9_addsub_cry_14_c_RNIO7DP9_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40173\,
            in1 => \N__39981\,
            in2 => \_gnd_net_\,
            in3 => \N__35260\,
            lcout => \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_10_s0_c_RNO_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__52034\,
            in1 => \N__53895\,
            in2 => \N__53236\,
            in3 => \N__51796\,
            lcout => \ALU.r0_12_prm_6_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_15_s0_c_RNO_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55861\,
            in1 => \N__53894\,
            in2 => \_gnd_net_\,
            in3 => \N__37273\,
            lcout => \ALU.r0_12_prm_1_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_14_s1_c_RNO_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010101111"
        )
    port map (
            in0 => \N__53893\,
            in1 => \_gnd_net_\,
            in2 => \N__55847\,
            in3 => \N__49054\,
            lcout => \ALU.r0_12_prm_1_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_8_s1_c_RNO_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55776\,
            in2 => \_gnd_net_\,
            in3 => \N__39391\,
            lcout => \ALU.r0_12_prm_2_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_12_s1_c_RNO_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55772\,
            in2 => \_gnd_net_\,
            in3 => \N__37636\,
            lcout => \ALU.r0_12_prm_2_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_3_c_RNO_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49423\,
            in2 => \_gnd_net_\,
            in3 => \N__44365\,
            lcout => \ALU.un14_log_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s0_c_RNO_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55521\,
            in2 => \_gnd_net_\,
            in3 => \N__36141\,
            lcout => \ALU.r0_12_prm_8_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_12_s0_c_RNO_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55930\,
            in2 => \_gnd_net_\,
            in3 => \N__37637\,
            lcout => \ALU.r0_12_prm_2_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_9_s0_c_RNO_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55931\,
            in1 => \N__53780\,
            in2 => \_gnd_net_\,
            in3 => \N__42391\,
            lcout => \ALU.r0_12_prm_1_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIKUTI9_13_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__53778\,
            in1 => \N__41555\,
            in2 => \N__54607\,
            in3 => \N__41301\,
            lcout => \ALU.lshift_3_ns_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_15_s0_c_RNO_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36235\,
            lcout => \ALU.r0_12_prm_2_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s0_c_RNO_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__51103\,
            in1 => \_gnd_net_\,
            in2 => \N__51537\,
            in3 => \N__41706\,
            lcout => \ALU.rshift_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_10_s0_c_RNO_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35632\,
            lcout => \ALU.r0_12_prm_2_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_12_s1_c_RNO_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__53779\,
            in1 => \N__54447\,
            in2 => \N__53104\,
            in3 => \N__41302\,
            lcout => \ALU.r0_12_prm_4_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_11_s1_c_RNO_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55933\,
            in2 => \_gnd_net_\,
            in3 => \N__35834\,
            lcout => \ALU.r0_12_prm_2_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_1_c_RNO_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54860\,
            in1 => \N__48652\,
            in2 => \N__53221\,
            in3 => \N__46831\,
            lcout => \ALU.r0_12_prm_5_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_12_s1_c_RNO_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__54001\,
            in1 => \N__55932\,
            in2 => \_gnd_net_\,
            in3 => \N__37576\,
            lcout => \ALU.r0_12_prm_1_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIKU3HJ_10_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54859\,
            in1 => \N__39358\,
            in2 => \_gnd_net_\,
            in3 => \N__35785\,
            lcout => OPEN,
            ltout => \ALU.r5_RNIKU3HJZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIQK1V71_5_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51089\,
            in2 => \N__35779\,
            in3 => \N__38943\,
            lcout => \ALU.r4_RNIQK1V71Z0Z_5\,
            ltout => \ALU.r4_RNIQK1V71Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI8E2N22_2_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51523\,
            in2 => \N__35776\,
            in3 => \N__41025\,
            lcout => \ALU.lshift_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_11_s0_c_RNO_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__35748\,
            in1 => \N__55946\,
            in2 => \_gnd_net_\,
            in3 => \N__54000\,
            lcout => \ALU.r0_12_prm_1_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINPPC9_14_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47194\,
            in2 => \_gnd_net_\,
            in3 => \N__47032\,
            lcout => \ALU.un14_log_0_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI5P1F5_15_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54611\,
            in1 => \N__54024\,
            in2 => \N__53222\,
            in3 => \N__40106\,
            lcout => \ALU.r5_RNI5P1F5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_14_s0_c_RNO_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55939\,
            in2 => \_gnd_net_\,
            in3 => \N__49132\,
            lcout => \ALU.r0_12_prm_2_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s0_c_RNO_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36037\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \ALU.r0_12_prm_8_15_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s0_c_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36027\,
            in2 => \N__35995\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_15_s0_cy\,
            carryout => \ALU.r0_12_prm_8_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_15_s0_c_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39898\,
            in2 => \N__35982\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_15_s0\,
            carryout => \ALU.r0_12_prm_7_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_15_s0_c_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35962\,
            in2 => \N__35953\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_15_s0\,
            carryout => \ALU.r0_12_prm_6_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_15_s0_c_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35920\,
            in2 => \N__35910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_15_s0\,
            carryout => \ALU.r0_12_prm_5_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_15_s0_c_inv_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35887\,
            in2 => \N__35874\,
            in3 => \N__40156\,
            lcout => \ALU.a_i_15\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_15_s0\,
            carryout => \ALU.r0_12_prm_4_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_15_s0_c_inv_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36265\,
            in2 => \_gnd_net_\,
            in3 => \N__55234\,
            lcout => \ALU.r0_12_prm_3_15_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_15_s0\,
            carryout => \ALU.r0_12_prm_3_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_15_s0_c_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36252\,
            in2 => \N__36214\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_15_s0\,
            carryout => \ALU.r0_12_prm_2_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_15_s0_c_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36202\,
            in2 => \N__37290\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \ALU.r0_12_s0_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s0_15_THRU_LUT4_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36193\,
            lcout => \ALU.r0_12_s0_15_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIB8HG5_12_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54615\,
            in1 => \N__54025\,
            in2 => \N__53223\,
            in3 => \N__41351\,
            lcout => \ALU.r5_RNIB8HG5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s1_c_RNO_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55535\,
            in2 => \_gnd_net_\,
            in3 => \N__36140\,
            lcout => \ALU.r0_12_prm_8_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_10_s1_c_RNO_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55959\,
            in1 => \N__54049\,
            in2 => \_gnd_net_\,
            in3 => \N__36100\,
            lcout => \ALU.r0_12_prm_1_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_12_s0_c_RNO_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__54050\,
            in1 => \N__55960\,
            in2 => \_gnd_net_\,
            in3 => \N__37586\,
            lcout => \ALU.r0_12_prm_1_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_0_s1_c_RNO_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__53968\,
            in1 => \N__54806\,
            in2 => \N__53154\,
            in3 => \N__49015\,
            lcout => \ALU.r0_12_prm_4_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_0_s1_c_RNO_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54810\,
            in1 => \N__49014\,
            in2 => \N__53153\,
            in3 => \N__38030\,
            lcout => \ALU.r0_12_prm_5_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_6_s1_c_RNO_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55841\,
            in1 => \N__53969\,
            in2 => \_gnd_net_\,
            in3 => \N__38206\,
            lcout => \ALU.r0_12_prm_1_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJTDS9_0_5_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__53967\,
            in1 => \N__45494\,
            in2 => \N__54886\,
            in3 => \N__42848\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI9H7SJ_6_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__54805\,
            in1 => \N__43429\,
            in2 => \N__36349\,
            in3 => \N__44603\,
            lcout => \ALU.r4_RNI9H7SJZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_0_s1_c_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37504\,
            in2 => \N__40705\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_2_0_\,
            carryout => \ALU.r0_12_prm_8_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_0_s1_c_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36346\,
            in2 => \N__36447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_0_s1\,
            carryout => \ALU.r0_12_prm_7_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_0_s1_c_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36334\,
            in2 => \N__36316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_0_s1\,
            carryout => \ALU.r0_12_prm_6_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_0_s1_c_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36292\,
            in2 => \N__37752\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_0_s1\,
            carryout => \ALU.r0_12_prm_5_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_0_s1_c_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36286\,
            in2 => \N__36280\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_0_s1\,
            carryout => \ALU.r0_12_prm_4_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_0_s1_c_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36463\,
            in2 => \N__36448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_0_s1\,
            carryout => \ALU.r0_12_prm_3_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_0_s1_c_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38116\,
            in2 => \N__40618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_0_s1\,
            carryout => \ALU.r0_12_prm_2_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_0_s1_c_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36415\,
            in2 => \N__36400\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_2_0_s1\,
            carryout => \ALU.r0_12_s1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_0_THRU_LUT4_0_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36385\,
            lcout => \ALU.r0_12_s1_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_5_s0_c_RNO_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__45405\,
            in1 => \N__54651\,
            in2 => \N__53228\,
            in3 => \N__45260\,
            lcout => \ALU.r0_12_prm_5_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIO5SA91_2_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__51080\,
            in1 => \N__48166\,
            in2 => \N__51491\,
            in3 => \N__41118\,
            lcout => \ALU.rshift_15_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_4_c_RNO_0_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42825\,
            in2 => \_gnd_net_\,
            in3 => \N__40534\,
            lcout => \ALU.r0_12_prm_5_4_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI97EK9_0_5_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__53781\,
            in1 => \N__45404\,
            in2 => \N__54789\,
            in3 => \N__43420\,
            lcout => \ALU.rshift_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_0_s0_c_RNO_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40607\,
            in2 => \_gnd_net_\,
            in3 => \N__55736\,
            lcout => \ALU.r0_12_prm_2_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_1_c_RNO_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53807\,
            in1 => \N__48617\,
            in2 => \N__53158\,
            in3 => \N__46749\,
            lcout => \ALU.r0_12_prm_6_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIK9PV9_15_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000011"
        )
    port map (
            in0 => \N__54702\,
            in1 => \N__51003\,
            in2 => \N__51482\,
            in3 => \N__50621\,
            lcout => \ALU.rshift_15_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_3_c_RNO_0_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49341\,
            in2 => \_gnd_net_\,
            in3 => \N__44360\,
            lcout => \ALU.r0_12_prm_5_3_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIODO6K_7_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__36826\,
            in1 => \N__46190\,
            in2 => \N__54813\,
            in3 => \N__44595\,
            lcout => \ALU.r4_RNIODO6KZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI9OH6A_1_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53806\,
            in1 => \N__48989\,
            in2 => \_gnd_net_\,
            in3 => \N__48616\,
            lcout => OPEN,
            ltout => \ALU.r4_RNI9OH6AZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJH1SA_1_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__54701\,
            in1 => \N__51268\,
            in2 => \N__36820\,
            in3 => \N__51002\,
            lcout => \ALU.lshift_15_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_6_s0_c_RNO_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55517\,
            in2 => \_gnd_net_\,
            in3 => \N__37688\,
            lcout => \ALU.r0_12_prm_8_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_a10_b_4_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__36817\,
            in1 => \N__36805\,
            in2 => \N__36768\,
            in3 => \N__40488\,
            lcout => \ALU.a10_b_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIHENK8_0_7_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44805\,
            in2 => \_gnd_net_\,
            in3 => \N__44537\,
            lcout => \ALU.r4_RNIHENK8_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIFR136_7_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__44538\,
            in1 => \N__52719\,
            in2 => \N__54885\,
            in3 => \N__53874\,
            lcout => \ALU.r4_RNIFR136Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIF01FK_2_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__49412\,
            in1 => \N__54796\,
            in2 => \N__36895\,
            in3 => \N__48400\,
            lcout => \ALU.r4_RNIF01FKZ0Z_2\,
            ltout => \ALU.r4_RNIF01FKZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIJCHBK1_6_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__51414\,
            in1 => \N__36886\,
            in2 => \N__36877\,
            in3 => \N__36874\,
            lcout => \ALU.lshift_9\,
            ltout => \ALU.lshift_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s1_c_RNO_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36856\,
            in3 => \N__55513\,
            lcout => \ALU.r0_12_prm_8_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s0_c_RNO_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__42561\,
            in1 => \_gnd_net_\,
            in2 => \N__55534\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_8_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_4_c_RNO_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52718\,
            in2 => \_gnd_net_\,
            in3 => \N__38463\,
            lcout => \ALU.r0_12_prm_7_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_7_s0_c_THRU_CRY_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44169\,
            in2 => \N__44173\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \ALU.r0_12_prm_8_7_s0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_7_s0_c_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42985\,
            in2 => \N__44125\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_7_s0_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_7_s0_c_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48079\,
            in2 => \N__48004\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_7_s0\,
            carryout => \ALU.r0_12_prm_7_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_7_s0_c_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44095\,
            in2 => \N__36976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_7_s0\,
            carryout => \ALU.r0_12_prm_6_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_7_s0_c_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44055\,
            in2 => \N__43159\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_7_s0\,
            carryout => \ALU.r0_12_prm_5_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_7_s0_c_inv_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44028\,
            in2 => \N__36964\,
            in3 => \N__44596\,
            lcout => \ALU.a_i_7\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_7_s0\,
            carryout => \ALU.r0_12_prm_4_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_7_s0_c_inv_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55282\,
            in1 => \N__36955\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_7_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_7_s0\,
            carryout => \ALU.r0_12_prm_3_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_7_s0_c_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44013\,
            in2 => \N__38953\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_7_s0\,
            carryout => \ALU.r0_12_prm_2_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_7_s0_c_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45005\,
            in2 => \N__36949\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \ALU.r0_12_s0_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_7_s0_c_RNIJOSTUN1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44914\,
            in1 => \N__36940\,
            in2 => \_gnd_net_\,
            in3 => \N__36925\,
            lcout => \ALU.r0_12_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_7_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38711\,
            lcout => r1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56241\,
            ce => \N__47559\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s0_c_RNO_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38884\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \ALU.r0_12_prm_8_5_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s0_c_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48151\,
            in2 => \N__48118\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_5_s0_cy\,
            carryout => \ALU.r0_12_prm_8_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_5_s0_c_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47267\,
            in2 => \N__37060\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_5_s0\,
            carryout => \ALU.r0_12_prm_7_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_5_s0_c_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44944\,
            in2 => \N__37042\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_5_s0\,
            carryout => \ALU.r0_12_prm_6_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_5_s0_c_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45766\,
            in2 => \N__37024\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_5_s0\,
            carryout => \ALU.r0_12_prm_5_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_5_s0_c_inv_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45714\,
            in2 => \N__37012\,
            in3 => \N__45510\,
            lcout => \ALU.a_i_5\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_5_s0\,
            carryout => \ALU.r0_12_prm_4_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_5_s0_c_inv_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55272\,
            in1 => \N__36994\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_5_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_5_s0\,
            carryout => \ALU.r0_12_prm_3_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_5_s0_c_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45687\,
            in2 => \N__36988\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_5_s0\,
            carryout => \ALU.r0_12_prm_2_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_5_s0_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45625\,
            in2 => \N__44188\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \ALU.r0_12_s0_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_5_s0_c_RNITPI7KJ_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45592\,
            in1 => \N__37234\,
            in2 => \_gnd_net_\,
            in3 => \N__37219\,
            lcout => \ALU.r0_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_5_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37150\,
            lcout => r1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56249\,
            ce => \N__47543\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s0_c_RNO_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38614\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \ALU.r0_12_prm_8_8_s0_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s0_c_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38917\,
            in2 => \N__39331\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_8_s0_cy\,
            carryout => \ALU.r0_12_prm_8_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_8_s0_c_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38893\,
            in2 => \N__39292\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_8_s0\,
            carryout => \ALU.r0_12_prm_7_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_8_s0_c_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37084\,
            in2 => \N__39264\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_8_s0\,
            carryout => \ALU.r0_12_prm_6_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_8_s0_c_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40774\,
            in2 => \N__42025\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_8_s0\,
            carryout => \ALU.r0_12_prm_5_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_8_s0_c_inv_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38980\,
            in2 => \N__39234\,
            in3 => \N__46180\,
            lcout => \ALU.a_i_8\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_8_s0\,
            carryout => \ALU.r0_12_prm_4_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_8_s0_c_inv_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55268\,
            in1 => \N__37066\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_3_8_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_8_s0\,
            carryout => \ALU.r0_12_prm_3_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_8_s0_c_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39401\,
            in2 => \N__39370\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_8_s0\,
            carryout => \ALU.r0_12_prm_2_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_8_s0_c_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39618\,
            in2 => \N__37306\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \ALU.r0_12_s0_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s0_8_THRU_LUT4_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37309\,
            lcout => \ALU.r0_12_s0_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_8_s1_c_RNO_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__39617\,
            in1 => \N__55903\,
            in2 => \_gnd_net_\,
            in3 => \N__53897\,
            lcout => \ALU.r0_12_prm_1_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_8_s0_c_RNO_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55902\,
            in1 => \N__53896\,
            in2 => \_gnd_net_\,
            in3 => \N__39616\,
            lcout => \ALU.r0_12_prm_1_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_15_s1_c_RNO_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55940\,
            in1 => \N__54002\,
            in2 => \_gnd_net_\,
            in3 => \N__37283\,
            lcout => \ALU.r0_12_prm_1_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNISU5D9_0_9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47478\,
            lcout => \ALU.r4_RNISU5D9_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNISP2L9_1_12_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41354\,
            lcout => \ALU.r5_RNISP2L9_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_12_s1_c_RNO_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__41353\,
            in1 => \N__53064\,
            in2 => \_gnd_net_\,
            in3 => \N__39876\,
            lcout => \ALU.r0_12_prm_7_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_9_s1_c_RNO_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53175\,
            in1 => \N__47477\,
            in2 => \_gnd_net_\,
            in3 => \N__52321\,
            lcout => \ALU.r0_12_prm_7_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s1_c_RNO_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101001011"
        )
    port map (
            in0 => \N__51441\,
            in1 => \N__37485\,
            in2 => \N__55537\,
            in3 => \N__41024\,
            lcout => \ALU.r0_12_prm_8_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s1_c_RNO_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38905\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \ALU.r0_12_prm_8_12_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s1_c_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37474\,
            in2 => \N__37464\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_12_s1_cy\,
            carryout => \ALU.r0_12_prm_8_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_12_s1_c_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37447\,
            in2 => \N__37441\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_12_s1\,
            carryout => \ALU.r0_12_prm_7_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_12_s1_c_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37414\,
            in2 => \N__39718\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_12_s1\,
            carryout => \ALU.r0_12_prm_6_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_12_s1_c_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37384\,
            in2 => \N__37362\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_12_s1\,
            carryout => \ALU.r0_12_prm_5_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_12_s1_c_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37345\,
            in2 => \N__37333\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_12_s1\,
            carryout => \ALU.r0_12_prm_4_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_12_s1_c_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55280\,
            in2 => \N__56508\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_12_s1\,
            carryout => \ALU.r0_12_prm_3_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_12_s1_c_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37650\,
            in2 => \N__37615\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_12_s1\,
            carryout => \ALU.r0_12_prm_2_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_12_s1_c_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37603\,
            in2 => \N__37593\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \ALU.r0_12_s1_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_12_THRU_LUT4_0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37555\,
            lcout => \ALU.r0_12_s1_12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_15_s1_c_RNO_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54782\,
            in1 => \N__40158\,
            in2 => \N__52963\,
            in3 => \N__40007\,
            lcout => \ALU.r0_12_prm_5_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_15_s1_c_RNO_1_LC_13_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__54802\,
            in1 => \N__53964\,
            in2 => \N__50679\,
            in3 => \N__40183\,
            lcout => \ALU.r0_12_prm_8_15_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \params_3_LC_13_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__54803\,
            in1 => \N__51224\,
            in2 => \N__50932\,
            in3 => \N__53966\,
            lcout => \paramsZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56227\,
            ce => \N__56057\,
            sr => \_gnd_net_\
        );

    \params_2_LC_13_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__53965\,
            in1 => \N__50856\,
            in2 => \_gnd_net_\,
            in3 => \N__54804\,
            lcout => \paramsZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56227\,
            ce => \N__56057\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_0_s1_c_RNO_LC_13_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55489\,
            in2 => \_gnd_net_\,
            in3 => \N__40694\,
            lcout => \ALU.r0_12_prm_8_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIAV175_15_LC_13_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__54801\,
            in1 => \N__53963\,
            in2 => \N__50931\,
            in3 => \N__40182\,
            lcout => \ALU.r5_RNIAV175Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.lshift63_2_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51212\,
            in2 => \_gnd_net_\,
            in3 => \N__50873\,
            lcout => \ALU.lshift63Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_0_s1_c_RNO_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55722\,
            in2 => \_gnd_net_\,
            in3 => \N__40606\,
            lcout => \ALU.r0_12_prm_2_0_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIHENK8_7_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44784\,
            in2 => \_gnd_net_\,
            in3 => \N__44600\,
            lcout => \ALU.un14_log_0_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_RNO_2_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__50874\,
            in1 => \N__38110\,
            in2 => \N__51296\,
            in3 => \N__38098\,
            lcout => OPEN,
            ltout => \ALU.rshift_15_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_RNO_1_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__38083\,
            in1 => \N__51221\,
            in2 => \N__38062\,
            in3 => \N__38059\,
            lcout => \ALU.rshift_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_6_s0_c_RNO_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55723\,
            in2 => \_gnd_net_\,
            in3 => \N__38265\,
            lcout => \ALU.r0_12_prm_2_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNID26E8_0_0_LC_13_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49000\,
            in2 => \_gnd_net_\,
            in3 => \N__38032\,
            lcout => \ALU.r4_RNID26E8_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_6_s0_c_THRU_CRY_0_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37730\,
            in2 => \N__37735\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_3_0_\,
            carryout => \ALU.r0_12_prm_8_6_s0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_6_s0_c_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37693\,
            in2 => \N__37663\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_6_s0_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_6_s0_c_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41649\,
            in2 => \N__41602\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_6_s0\,
            carryout => \ALU.r0_12_prm_7_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_6_s0_c_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38365\,
            in2 => \N__41587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_6_s0\,
            carryout => \ALU.r0_12_prm_6_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_6_s0_c_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38341\,
            in2 => \N__43174\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_6_s0\,
            carryout => \ALU.r0_12_prm_5_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_6_s0_c_inv_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38289\,
            in2 => \N__38317\,
            in3 => \N__43436\,
            lcout => \ALU.a_i_6\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_6_s0\,
            carryout => \ALU.r0_12_prm_4_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_6_s0_c_inv_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38275\,
            in3 => \N__55172\,
            lcout => \ALU.r0_12_prm_3_6_s0_sf\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_6_s0\,
            carryout => \ALU.r0_12_prm_3_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_6_s0_c_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38258\,
            in2 => \N__38215\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_6_s0\,
            carryout => \ALU.r0_12_prm_2_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_6_s0_c_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38205\,
            in2 => \N__38161\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_4_0_\,
            carryout => \ALU.r0_12_s0_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_6_s0_c_RNINEODV21_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38146\,
            in1 => \N__38134\,
            in2 => \_gnd_net_\,
            in3 => \N__38119\,
            lcout => \ALU.r0_12_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r1_6_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38815\,
            lcout => r1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56230\,
            ce => \N__47577\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_THRU_CRY_0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41067\,
            in2 => \N__41071\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_5_0_\,
            carryout => \ALU.r0_12_prm_8_4_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41803\,
            in2 => \N__40756\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_4_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_4_c_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38467\,
            in2 => \N__38434\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_4\,
            carryout => \ALU.r0_12_prm_7_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_4_c_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38425\,
            in2 => \N__38410\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_4\,
            carryout => \ALU.r0_12_prm_6_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_4_c_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40342\,
            in2 => \N__38395\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_4\,
            carryout => \ALU.r0_12_prm_5_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_4_c_inv_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38383\,
            in2 => \N__42616\,
            in3 => \N__42851\,
            lcout => \ALU.a_i_4\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_4\,
            carryout => \ALU.r0_12_prm_4_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_4_c_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38530\,
            in2 => \N__38377\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_4\,
            carryout => \ALU.r0_12_prm_3_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_4_c_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38602\,
            in2 => \N__38578\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_4\,
            carryout => \ALU.r0_12_prm_2_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_4_c_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41761\,
            in2 => \N__41737\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \ALU.r0_12_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_4_THRU_LUT4_0_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38659\,
            lcout => \ALU.r0_12_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI0QK3K_11_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38656\,
            in1 => \N__54795\,
            in2 => \_gnd_net_\,
            in3 => \N__38632\,
            lcout => \ALU.r5_RNI0QK3KZ0Z_11\,
            ltout => \ALU.r5_RNI0QK3KZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s0_c_RNO_1_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__50984\,
            in1 => \N__51359\,
            in2 => \N__38617\,
            in3 => \N__41686\,
            lcout => \ALU.rshift_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s1_c_RNO_1_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__41687\,
            in1 => \N__50985\,
            in2 => \N__51446\,
            in3 => \N__41091\,
            lcout => \ALU.r0_12_prm_8_8_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_4_c_RNO_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55729\,
            in2 => \_gnd_net_\,
            in3 => \N__38598\,
            lcout => \ALU.r0_12_prm_2_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_4_c_RNO_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__55261\,
            in1 => \N__38569\,
            in2 => \_gnd_net_\,
            in3 => \N__38548\,
            lcout => \ALU.r0_12_prm_3_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIR63FA_4_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__53805\,
            in1 => \N__42850\,
            in2 => \N__54884\,
            in3 => \N__49408\,
            lcout => \ALU.lshift_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s1_c_RNO_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55400\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39317\,
            lcout => \ALU.r0_12_prm_8_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_7_s0_c_RNO_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55730\,
            in2 => \_gnd_net_\,
            in3 => \N__44014\,
            lcout => \ALU.r0_12_prm_2_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNILGU5F1_5_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__41056\,
            in1 => \N__38944\,
            in2 => \N__51301\,
            in3 => \N__41043\,
            lcout => \ALU.lshift_8\,
            ltout => \ALU.lshift_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s0_c_RNO_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38920\,
            in3 => \N__55399\,
            lcout => \ALU.r0_12_prm_8_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_12_s1_c_RNO_1_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51231\,
            in1 => \N__51032\,
            in2 => \_gnd_net_\,
            in3 => \N__41685\,
            lcout => \ALU.r0_12_prm_8_12_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_8_s0_c_RNO_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__52544\,
            in1 => \N__46382\,
            in2 => \_gnd_net_\,
            in3 => \N__46220\,
            lcout => \ALU.r0_12_prm_7_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s0_c_RNO_1_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__51102\,
            in1 => \N__43144\,
            in2 => \N__51302\,
            in3 => \N__41662\,
            lcout => \ALU.rshift_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r6_6_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38827\,
            lcout => r6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => \N__45846\,
            sr => \_gnd_net_\
        );

    \ALU.r6_7_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38712\,
            lcout => r6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => \N__45846\,
            sr => \_gnd_net_\
        );

    \ALU.r6_8_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39494\,
            lcout => r6_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => \N__45846\,
            sr => \_gnd_net_\
        );

    \ALU.r6_2_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40243\,
            lcout => r6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => \N__45846\,
            sr => \_gnd_net_\
        );

    \ALU.r6_3_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50159\,
            lcout => r6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => \N__45846\,
            sr => \_gnd_net_\
        );

    \ALU.r6_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39043\,
            lcout => r6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => \N__45846\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_RNO_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000001111"
        )
    port map (
            in0 => \N__51039\,
            in1 => \N__51244\,
            in2 => \N__55522\,
            in3 => \N__50765\,
            lcout => \ALU.r0_12_prm_8_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIN3236_8_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__52819\,
            in1 => \N__54057\,
            in2 => \N__46227\,
            in3 => \N__54914\,
            lcout => \ALU.r4_RNIN3236Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_8_s1_c_RNO_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__52820\,
            in1 => \N__54058\,
            in2 => \N__46228\,
            in3 => \N__54915\,
            lcout => \ALU.r0_12_prm_4_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_RNO_3_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010101000101"
        )
    port map (
            in0 => \N__38974\,
            in1 => \N__42861\,
            in2 => \N__54924\,
            in3 => \N__49425\,
            lcout => OPEN,
            ltout => \ALU.r0_12_prm_8_1_c_RNOZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_RNO_2_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__51245\,
            in1 => \N__51040\,
            in2 => \N__38956\,
            in3 => \N__41796\,
            lcout => OPEN,
            ltout => \ALU.rshift_15_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_RNO_1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51246\,
            in1 => \N__43140\,
            in2 => \N__39346\,
            in3 => \N__43065\,
            lcout => \ALU.rshift_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s1_c_RNO_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39343\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \ALU.r0_12_prm_8_8_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_8_s1_c_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39327\,
            in2 => \N__39304\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_8_s1_cy\,
            carryout => \ALU.r0_12_prm_8_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_8_s1_c_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39291\,
            in2 => \N__45922\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_8_s1\,
            carryout => \ALU.r0_12_prm_7_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_8_s1_c_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39265\,
            in2 => \N__42007\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_8_s1\,
            carryout => \ALU.r0_12_prm_6_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_8_s1_c_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42021\,
            in2 => \N__45580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_8_s1\,
            carryout => \ALU.r0_12_prm_5_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_8_s1_c_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39241\,
            in2 => \N__39235\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_8_s1\,
            carryout => \ALU.r0_12_prm_4_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_8_s1_c_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55192\,
            in2 => \N__56475\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_8_s1\,
            carryout => \ALU.r0_12_prm_3_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_8_s1_c_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39402\,
            in2 => \N__39217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_8_s1\,
            carryout => \ALU.r0_12_prm_2_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_8_s1_c_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39622\,
            in2 => \N__39589\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \ALU.r0_12_s1_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_8_s0_c_RNIO9TN7H2_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__39580\,
            in1 => \N__39562\,
            in2 => \N__39538\,
            in3 => \N__39529\,
            lcout => \ALU.r0_12_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_8_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39472\,
            lcout => r0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56252\,
            ce => \N__49716\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_9_s1_c_RNO_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42440\,
            lcout => \ALU.r0_12_prm_2_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_8_s0_c_RNO_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55899\,
            in2 => \_gnd_net_\,
            in3 => \N__39403\,
            lcout => \ALU.r0_12_prm_2_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNITTMB9_12_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53996\,
            in1 => \N__41352\,
            in2 => \_gnd_net_\,
            in3 => \N__40962\,
            lcout => \ALU.r5_RNITTMB9Z0Z_12\,
            ltout => \ALU.r5_RNITTMB9Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI355TI_13_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54858\,
            in1 => \_gnd_net_\,
            in2 => \N__39349\,
            in3 => \N__39709\,
            lcout => \ALU.r5_RNI355TIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_9_s1_c_RNO_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54584\,
            in1 => \N__47482\,
            in2 => \N__53205\,
            in3 => \N__52221\,
            lcout => \ALU.r0_12_prm_5_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_9_s1_c_RNO_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55901\,
            in1 => \N__53997\,
            in2 => \_gnd_net_\,
            in3 => \N__42395\,
            lcout => \ALU.r0_12_prm_1_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s1_c_RNO_1_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__51037\,
            in1 => \N__43139\,
            in2 => \N__51304\,
            in3 => \N__43066\,
            lcout => \ALU.r0_12_prm_8_9_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_14_s1_c_RNO_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54906\,
            in1 => \N__53960\,
            in2 => \N__53206\,
            in3 => \N__47008\,
            lcout => \ALU.r0_12_prm_4_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNITG1F5_14_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__53961\,
            in1 => \N__54907\,
            in2 => \N__53239\,
            in3 => \N__47031\,
            lcout => \ALU.r5_RNITG1F5Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_14_s0_c_RNO_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__47185\,
            in1 => \N__53180\,
            in2 => \N__54923\,
            in3 => \N__47010\,
            lcout => \ALU.r0_12_prm_5_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s0_c_RNO_1_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51300\,
            in1 => \N__51038\,
            in2 => \_gnd_net_\,
            in3 => \N__43128\,
            lcout => \ALU.rshift_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_14_s0_c_RNO_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__47184\,
            in1 => \N__53962\,
            in2 => \N__53207\,
            in3 => \N__47009\,
            lcout => \ALU.r0_12_prm_6_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s0_c_RNO_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__47969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55533\,
            lcout => \ALU.r0_12_prm_8_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_14_s1_c_RNO_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53176\,
            in1 => \N__47183\,
            in2 => \_gnd_net_\,
            in3 => \N__47030\,
            lcout => \ALU.r0_12_prm_7_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIUH636_3_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54905\,
            in1 => \N__53958\,
            in2 => \N__53182\,
            in3 => \N__49426\,
            lcout => \ALU.r4_RNIUH636Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_15_s0_c_RNO_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53014\,
            in1 => \N__40157\,
            in2 => \_gnd_net_\,
            in3 => \N__40008\,
            lcout => \ALU.r0_12_prm_7_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_14_s1_c_RNO_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53957\,
            in1 => \N__47197\,
            in2 => \N__53181\,
            in3 => \N__47052\,
            lcout => \ALU.r0_12_prm_6_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_13_s1_c_RNO_1_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43127\,
            in1 => \N__51303\,
            in2 => \_gnd_net_\,
            in3 => \N__51099\,
            lcout => \ALU.r0_12_prm_8_13_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_12_s1_c_RNO_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010010101"
        )
    port map (
            in0 => \N__39872\,
            in1 => \N__53959\,
            in2 => \N__53183\,
            in3 => \N__41355\,
            lcout => \ALU.r0_12_prm_6_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIPV8A9_0_13_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53956\,
            in1 => \N__41478\,
            in2 => \_gnd_net_\,
            in3 => \N__47050\,
            lcout => \ALU.r5_RNIPV8A9_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_THRU_CRY_0_LC_14_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39696\,
            in2 => \N__39700\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_1_0_\,
            carryout => \ALU.r0_12_prm_8_2_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_LC_14_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40204\,
            in2 => \N__40213\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_2_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_2_c_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40746\,
            in2 => \N__40714\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_2\,
            carryout => \ALU.r0_12_prm_7_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_2_c_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40543\,
            in2 => \N__42937\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_2\,
            carryout => \ALU.r0_12_prm_6_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_2_c_LC_14_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40336\,
            in2 => \N__43723\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_2\,
            carryout => \ALU.r0_12_prm_5_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_2_c_inv_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40324\,
            in2 => \N__40312\,
            in3 => \N__48405\,
            lcout => \ALU.a_i_2\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_2\,
            carryout => \ALU.r0_12_prm_4_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_2_c_LC_14_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42874\,
            in2 => \N__42925\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_2\,
            carryout => \ALU.r0_12_prm_3_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_2_c_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40552\,
            in2 => \N__40579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_2\,
            carryout => \ALU.r0_12_prm_2_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_2_c_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43708\,
            in2 => \N__43678\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_2_0_\,
            carryout => \ALU.r0_12_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_2_THRU_LUT4_0_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40303\,
            lcout => \ALU.r0_12_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_RNO_0_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51223\,
            in1 => \N__50878\,
            in2 => \_gnd_net_\,
            in3 => \N__42204\,
            lcout => \ALU.lshift_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_2_c_RNO_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000110011"
        )
    port map (
            in0 => \N__51222\,
            in1 => \N__55491\,
            in2 => \N__50961\,
            in3 => \N__42203\,
            lcout => \ALU.r0_12_prm_8_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_0_s0_c_RNO_LC_14_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55490\,
            in2 => \_gnd_net_\,
            in3 => \N__40687\,
            lcout => \ALU.r0_12_prm_8_0_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_2_c_RNO_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53139\,
            in2 => \_gnd_net_\,
            in3 => \N__40747\,
            lcout => \ALU.r0_12_prm_7_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI80BM5_0_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__54811\,
            in1 => \N__53970\,
            in2 => \N__50669\,
            in3 => \N__48907\,
            lcout => \ALU.lshift_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIHENK8_1_7_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__44601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44789\,
            lcout => \ALU.r4_RNIHENK8_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIFQDK8_0_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56488\,
            in1 => \N__40648\,
            in2 => \_gnd_net_\,
            in3 => \N__48908\,
            lcout => \ALU.un2_addsub_axb_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_2_c_RNO_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55659\,
            in2 => \_gnd_net_\,
            in3 => \N__40572\,
            lcout => \ALU.r0_12_prm_2_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_2_c_RNO_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53971\,
            in1 => \N__48404\,
            in2 => \N__53231\,
            in3 => \N__43963\,
            lcout => \ALU.r0_12_prm_6_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_7_s1_c_RNO_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__44008\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55737\,
            lcout => \ALU.r0_12_prm_2_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIAHIIA_2_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54037\,
            in1 => \N__48323\,
            in2 => \_gnd_net_\,
            in3 => \N__48614\,
            lcout => \ALU.r4_RNIAHIIAZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_4_c_RNO_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54631\,
            in1 => \N__42867\,
            in2 => \N__52971\,
            in3 => \N__40522\,
            lcout => \ALU.r0_12_prm_5_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIN0D5A_0_10_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__54038\,
            in1 => \N__51840\,
            in2 => \N__52308\,
            in3 => \N__54626\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNILV3HJ_12_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__54627\,
            in1 => \N__41367\,
            in2 => \N__40999\,
            in3 => \N__40996\,
            lcout => \ALU.r5_RNILV3HJZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNID1636_1_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54040\,
            in1 => \N__54630\,
            in2 => \N__53103\,
            in3 => \N__48615\,
            lcout => \ALU.r4_RNID1636Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_8_s0_c_RNO_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54629\,
            in1 => \N__46465\,
            in2 => \N__52970\,
            in3 => \N__46216\,
            lcout => \ALU.r0_12_prm_5_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_5_s1_c_RNO_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54039\,
            in1 => \N__54628\,
            in2 => \N__53102\,
            in3 => \N__45506\,
            lcout => \ALU.r0_12_prm_4_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNIU6R05_0_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__53925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49012\,
            lcout => \ALU.N_610_1\,
            ltout => \ALU.N_610_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNILVIQF_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54718\,
            in2 => \N__40762\,
            in3 => \N__42294\,
            lcout => \ALU.r4_RNILVIQFZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIVFRGQ_0_2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__54719\,
            in1 => \N__42321\,
            in2 => \N__51087\,
            in3 => \N__41044\,
            lcout => \ALU.r4_RNIVFRGQ_0Z0Z_2\,
            ltout => \ALU.r4_RNIVFRGQ_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_RNO_0_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40759\,
            in3 => \N__51498\,
            lcout => \ALU.lshift_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIN0D5A_10_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__53923\,
            in1 => \N__51837\,
            in2 => \N__54823\,
            in3 => \N__52277\,
            lcout => \ALU.lshift_3_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_6_s0_c_RNO_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54041\,
            in1 => \N__43668\,
            in2 => \N__53144\,
            in3 => \N__43435\,
            lcout => \ALU.r0_12_prm_6_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNI7NOB9_13_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53924\,
            in1 => \N__41572\,
            in2 => \_gnd_net_\,
            in3 => \N__41366\,
            lcout => \ALU.r5_RNI7NOB9Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_7_s1_c_RNO_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54632\,
            in1 => \N__53926\,
            in2 => \N__53143\,
            in3 => \N__44543\,
            lcout => \ALU.r0_12_prm_4_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_RNO_2_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51026\,
            in1 => \N__41119\,
            in2 => \_gnd_net_\,
            in3 => \N__41090\,
            lcout => OPEN,
            ltout => \ALU.r0_12_prm_8_4_c_RNOZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_RNO_1_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51465\,
            in2 => \N__41074\,
            in3 => \N__41770\,
            lcout => \ALU.rshift_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNI80BM5_0_0_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000101"
        )
    port map (
            in0 => \N__51025\,
            in1 => \N__54899\,
            in2 => \N__51520\,
            in3 => \N__42316\,
            lcout => \ALU.lshift_15_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI6PL1L_2_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__41050\,
            in1 => \N__48401\,
            in2 => \N__54921\,
            in3 => \N__48640\,
            lcout => \ALU.r4_RNI6PL1LZ0Z_2\,
            ltout => \ALU.r4_RNI6PL1LZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIVFRGQ_2_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__51024\,
            in1 => \N__54898\,
            in2 => \N__41032\,
            in3 => \N__42317\,
            lcout => \ALU.r4_RNIVFRGQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_RNO_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011110101"
        )
    port map (
            in0 => \N__41809\,
            in1 => \_gnd_net_\,
            in2 => \N__51521\,
            in3 => \N__55476\,
            lcout => \ALU.r0_12_prm_8_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIRL1V71_7_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51027\,
            in1 => \N__43055\,
            in2 => \_gnd_net_\,
            in3 => \N__41797\,
            lcout => \ALU.r4_RNIRL1V71Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_4_c_RNO_3_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__54901\,
            in1 => \N__50611\,
            in2 => \N__51074\,
            in3 => \N__41727\,
            lcout => \ALU.r0_12_prm_8_4_c_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_4_c_RNO_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__53886\,
            in1 => \N__55806\,
            in2 => \_gnd_net_\,
            in3 => \N__41760\,
            lcout => \ALU.r0_12_prm_1_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r5_RNIUE7TI_13_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54900\,
            in1 => \N__50610\,
            in2 => \_gnd_net_\,
            in3 => \N__41726\,
            lcout => \ALU.r5_RNIUE7TIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s1_c_RNO_1_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__51028\,
            in1 => \N__43123\,
            in2 => \N__51522\,
            in3 => \N__41661\,
            lcout => \ALU.r0_12_prm_8_5_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI8B628_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45511\,
            in2 => \_gnd_net_\,
            in3 => \N__45179\,
            lcout => \ALU.un14_log_0_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_6_s0_c_RNO_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__52537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41650\,
            lcout => \ALU.r0_12_prm_7_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_5_s1_c_RNO_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55805\,
            in1 => \N__53885\,
            in2 => \_gnd_net_\,
            in3 => \N__45635\,
            lcout => \ALU.r0_12_prm_1_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_RNO_0_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46510\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50705\,
            lcout => \ALU.lshift_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_THRU_CRY_0_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41979\,
            in2 => \N__41983\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \ALU.r0_12_prm_8_1_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46471\,
            in2 => \N__41968\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_1_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_1_c_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41956\,
            in2 => \N__41923\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_1\,
            carryout => \ALU.r0_12_prm_7_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_1_c_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41905\,
            in2 => \N__46549\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_1\,
            carryout => \ALU.r0_12_prm_6_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_1_c_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41893\,
            in2 => \N__46534\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_1\,
            carryout => \ALU.r0_12_prm_5_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_1_c_inv_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41881\,
            in2 => \N__41869\,
            in3 => \N__48647\,
            lcout => \ALU.a_i_1\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_1\,
            carryout => \ALU.r0_12_prm_4_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_1_c_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41860\,
            in2 => \N__41842\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_1\,
            carryout => \ALU.r0_12_prm_3_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_1_c_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50547\,
            in2 => \N__50524\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_1\,
            carryout => \ALU.r0_12_prm_2_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_1_c_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42043\,
            in2 => \N__42061\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \ALU.r0_12_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_1_THRU_LUT4_0_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42166\,
            lcout => \ALU.r0_12_1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_5_s1_c_RNO_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55817\,
            in2 => \_gnd_net_\,
            in3 => \N__45673\,
            lcout => \ALU.r0_12_prm_2_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_1_c_RNO_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55818\,
            in1 => \N__54059\,
            in2 => \_gnd_net_\,
            in3 => \N__42057\,
            lcout => \ALU.r0_12_prm_1_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_9_s0_c_RNO_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010010101"
        )
    port map (
            in0 => \N__52324\,
            in1 => \N__54919\,
            in2 => \N__52938\,
            in3 => \N__47473\,
            lcout => \ALU.r0_12_prm_5_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIKUMQ8_0_8_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46178\,
            lcout => \ALU.r4_RNIKUMQ8_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_9_s1_c_RNO_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__53945\,
            in1 => \N__47471\,
            in2 => \N__53224\,
            in3 => \N__52323\,
            lcout => \ALU.r0_12_prm_6_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_8_s1_c_RNO_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54060\,
            in1 => \N__46460\,
            in2 => \N__52939\,
            in3 => \N__46179\,
            lcout => \ALU.r0_12_prm_6_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s0_c_RNO_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110011001"
        )
    port map (
            in0 => \N__42268\,
            in1 => \N__55481\,
            in2 => \N__42283\,
            in3 => \N__51519\,
            lcout => \ALU.r0_12_prm_8_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI67NNK_7_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000101"
        )
    port map (
            in0 => \N__42361\,
            in1 => \N__46219\,
            in2 => \N__54784\,
            in3 => \N__44610\,
            lcout => \ALU.r4_RNI67NNKZ0Z_7\,
            ltout => \ALU.r4_RNI67NNKZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNICN8R81_7_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51054\,
            in1 => \_gnd_net_\,
            in2 => \N__42349\,
            in3 => \N__42231\,
            lcout => \ALU.r4_RNICN8R81Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIU864P1_2_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51518\,
            in1 => \N__42279\,
            in2 => \_gnd_net_\,
            in3 => \N__42267\,
            lcout => \ALU.lshift_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI38O1G_2_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__42322\,
            in1 => \N__54625\,
            in2 => \N__51088\,
            in3 => \N__42298\,
            lcout => \ALU.r4_RNI38O1GZ0Z_2\,
            ltout => \ALU.r4_RNI38O1GZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_10_s1_c_RNO_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010010101"
        )
    port map (
            in0 => \N__55480\,
            in1 => \N__51514\,
            in2 => \N__42271\,
            in3 => \N__42266\,
            lcout => \ALU.r0_12_prm_8_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI6U6381_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__51058\,
            in1 => \N__42244\,
            in2 => \N__51533\,
            in3 => \N__42238\,
            lcout => OPEN,
            ltout => \ALU.lshift_15_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2FB1C2_4_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__42232\,
            in1 => \N__51513\,
            in2 => \N__42208\,
            in3 => \N__42199\,
            lcout => \ALU.lshift_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s1_c_RNO_0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42172\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \ALU.r0_12_prm_8_9_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s1_c_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42601\,
            in2 => \N__42585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_9_s1_cy\,
            carryout => \ALU.r0_12_prm_8_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_9_s1_c_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42550\,
            in2 => \N__42540\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_9_s1\,
            carryout => \ALU.r0_12_prm_7_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_9_s1_c_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42517\,
            in2 => \N__45543\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_9_s1\,
            carryout => \ALU.r0_12_prm_6_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_9_s1_c_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42508\,
            in2 => \N__42487\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_9_s1\,
            carryout => \ALU.r0_12_prm_5_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_9_s1_c_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52048\,
            in2 => \N__42478\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_9_s1\,
            carryout => \ALU.r0_12_prm_4_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_9_s1_c_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55223\,
            in2 => \N__56506\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_9_s1\,
            carryout => \ALU.r0_12_prm_3_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_9_s1_c_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42454\,
            in2 => \N__42447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_9_s1\,
            carryout => \ALU.r0_12_prm_2_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_9_s1_c_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42406\,
            in2 => \N__42400\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \ALU.r0_12_s1_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_9_THRU_LUT4_0_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42973\,
            lcout => \ALU.r0_12_s1_9_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINPPC9_1_14_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47196\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47011\,
            lcout => \ALU.r2_RNINPPC9_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r2_RNINPPC9_0_14_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47007\,
            in2 => \_gnd_net_\,
            in3 => \N__47195\,
            lcout => \ALU.r2_RNINPPC9_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_14_s1_c_RNO_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55904\,
            in2 => \_gnd_net_\,
            in3 => \N__49136\,
            lcout => \ALU.r0_12_prm_2_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_14_s0_c_RNO_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__47149\,
            in1 => \N__52937\,
            in2 => \_gnd_net_\,
            in3 => \N__47051\,
            lcout => \ALU.r0_12_prm_7_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_2_c_RNO_0_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48407\,
            in2 => \_gnd_net_\,
            in3 => \N__43961\,
            lcout => \ALU.un14_log_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_1_s_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42916\,
            in2 => \_gnd_net_\,
            in3 => \N__42897\,
            lcout => \ALU.mult_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_2_c_RNO_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__55138\,
            in1 => \N__42915\,
            in2 => \_gnd_net_\,
            in3 => \N__42896\,
            lcout => \ALU.r0_12_prm_3_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI87HO5_4_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54786\,
            in1 => \N__53134\,
            in2 => \N__54069\,
            in3 => \N__42866\,
            lcout => \ALU.r4_RNI87HO5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_2_c_RNO_0_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48406\,
            in2 => \_gnd_net_\,
            in3 => \N__43962\,
            lcout => \ALU.r0_12_prm_5_2_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_2_c_RNO_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011110101"
        )
    port map (
            in0 => \N__55640\,
            in1 => \_gnd_net_\,
            in2 => \N__54070\,
            in3 => \N__43707\,
            lcout => \ALU.r0_12_prm_1_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_6_s0_c_RNO_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54829\,
            in1 => \N__43669\,
            in2 => \N__53229\,
            in3 => \N__43430\,
            lcout => \ALU.r0_12_prm_5_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_7_s0_c_RNO_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111000011"
        )
    port map (
            in0 => \N__54785\,
            in1 => \N__44788\,
            in2 => \N__44611\,
            in3 => \N__53135\,
            lcout => \ALU.r0_12_prm_5_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_9_s0_c_RNO_1_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__51001\,
            in1 => \N__43138\,
            in2 => \N__51500\,
            in3 => \N__43054\,
            lcout => \ALU.rshift_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIO5SA91_5_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__51000\,
            in1 => \N__50773\,
            in2 => \N__51499\,
            in3 => \N__43012\,
            lcout => \ALU.lshift_7\,
            ltout => \ALU.lshift_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_7_s1_c_RNO_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__55446\,
            in1 => \_gnd_net_\,
            in2 => \N__42988\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_8_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_7_s1_c_RNO_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54812\,
            in1 => \N__44764\,
            in2 => \N__53230\,
            in3 => \N__44602\,
            lcout => \ALU.r0_12_prm_5_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_7_s0_c_RNO_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44111\,
            lcout => \ALU.r0_12_prm_8_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_7_s1_c_THRU_CRY_0_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44158\,
            in2 => \N__44168\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \ALU.r0_12_prm_8_7_s1_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_7_s1_c_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44131\,
            in2 => \N__44118\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_7_s1_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_7_s1_c_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48078\,
            in2 => \N__46852\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_7_s1\,
            carryout => \ALU.r0_12_prm_7_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_7_s1_c_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44371\,
            in2 => \N__44094\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_7_s1\,
            carryout => \ALU.r0_12_prm_6_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_7_s1_c_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44068\,
            in2 => \N__44062\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_7_s1\,
            carryout => \ALU.r0_12_prm_5_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_7_s1_c_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44041\,
            in2 => \N__44035\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_7_s1\,
            carryout => \ALU.r0_12_prm_4_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_7_s1_c_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55185\,
            in2 => \N__56504\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_7_s1\,
            carryout => \ALU.r0_12_prm_3_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_7_s1_c_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44009\,
            in2 => \N__43972\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_7_s1\,
            carryout => \ALU.r0_12_prm_2_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_7_s1_c_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45013\,
            in2 => \N__44977\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => \ALU.r0_12_s1_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_7_THRU_LUT4_0_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44917\,
            lcout => \ALU.r0_12_s1_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_5_s1_c_RNO_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54022\,
            in1 => \N__45462\,
            in2 => \N__53120\,
            in3 => \N__45261\,
            lcout => \ALU.r0_12_prm_6_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_RNO_1_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__44902\,
            in1 => \N__44872\,
            in2 => \N__51530\,
            in3 => \N__44857\,
            lcout => \ALU.rshift_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_3_c_RNO_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__49512\,
            in1 => \_gnd_net_\,
            in2 => \N__53122\,
            in3 => \_gnd_net_\,
            lcout => \ALU.r0_12_prm_7_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI2I2BV_2_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__50999\,
            in1 => \N__46502\,
            in2 => \N__51529\,
            in3 => \N__44823\,
            lcout => \ALU.lshift_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_7_s1_c_RNO_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010010011"
        )
    port map (
            in0 => \N__54023\,
            in1 => \N__44801\,
            in2 => \N__53121\,
            in3 => \N__44542\,
            lcout => \ALU.r0_12_prm_6_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_3_c_RNO_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54834\,
            in1 => \N__49417\,
            in2 => \N__53130\,
            in3 => \N__44346\,
            lcout => \ALU.r0_12_prm_5_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_5_s0_c_RNO_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55800\,
            in1 => \N__53928\,
            in2 => \_gnd_net_\,
            in3 => \N__45636\,
            lcout => \ALU.r0_12_prm_1_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNISU5D9_9_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47474\,
            in2 => \_gnd_net_\,
            in3 => \N__52310\,
            lcout => \ALU.un14_log_0_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_5_s1_c_RNO_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54833\,
            in1 => \N__45463\,
            in2 => \N__53129\,
            in3 => \N__45259\,
            lcout => \ALU.r0_12_prm_5_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s1_c_RNO_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55448\,
            in2 => \_gnd_net_\,
            in3 => \N__48136\,
            lcout => \ALU.r0_12_prm_8_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_3_c_RNO_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__55799\,
            in1 => \N__53929\,
            in2 => \_gnd_net_\,
            in3 => \N__50232\,
            lcout => \ALU.r0_12_prm_1_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_7_s1_c_RNO_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__53927\,
            in1 => \N__55798\,
            in2 => \_gnd_net_\,
            in3 => \N__45012\,
            lcout => \ALU.r0_12_prm_1_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s1_c_RNO_0_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44965\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \ALU.r0_12_prm_8_5_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s1_c_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44959\,
            in2 => \N__48150\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_5_s1_cy\,
            carryout => \ALU.r0_12_prm_8_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_5_s1_c_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47266\,
            in2 => \N__47209\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_5_s1\,
            carryout => \ALU.r0_12_prm_7_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_5_s1_c_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44953\,
            in2 => \N__44940\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_5_s1\,
            carryout => \ALU.r0_12_prm_6_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_5_s1_c_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45765\,
            in2 => \N__45742\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_5_s1\,
            carryout => \ALU.r0_12_prm_5_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_5_s1_c_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45733\,
            in2 => \N__45721\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_5_s1\,
            carryout => \ALU.r0_12_prm_4_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_5_s1_c_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55281\,
            in2 => \N__56481\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_5_s1\,
            carryout => \ALU.r0_12_prm_3_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_5_s1_c_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45700\,
            in2 => \N__45691\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_5_s1\,
            carryout => \ALU.r0_12_prm_2_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_5_s1_c_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45643\,
            in2 => \N__45637\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \ALU.r0_12_s1_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_5_THRU_LUT4_0_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45595\,
            lcout => \ALU.r0_12_s1_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_8_s1_c_RNO_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54641\,
            in1 => \N__46463\,
            in2 => \N__52941\,
            in3 => \N__46218\,
            lcout => \ALU.r0_12_prm_5_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_10_s0_c_RNO_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54640\,
            in1 => \N__52033\,
            in2 => \N__52940\,
            in3 => \N__51841\,
            lcout => \ALU.r0_12_prm_5_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_1_c_RNO_0_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48654\,
            in2 => \_gnd_net_\,
            in3 => \N__46837\,
            lcout => \ALU.r0_12_prm_5_1_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s0_c_RNO_1_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__50700\,
            in1 => \N__54639\,
            in2 => \_gnd_net_\,
            in3 => \N__50623\,
            lcout => \ALU.rshift_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_1_c_RNO_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__50701\,
            in1 => \N__55488\,
            in2 => \_gnd_net_\,
            in3 => \N__46509\,
            lcout => \ALU.r0_12_prm_8_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_8_s1_c_RNO_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53119\,
            in1 => \N__46464\,
            in2 => \_gnd_net_\,
            in3 => \N__46181\,
            lcout => \ALU.r0_12_prm_7_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_9_s0_c_RNO_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__53118\,
            in1 => \N__47472\,
            in2 => \_gnd_net_\,
            in3 => \N__52326\,
            lcout => \ALU.r0_12_prm_7_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_1_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__50436\,
            in1 => \N__50484\,
            in2 => \N__49800\,
            in3 => \N__54955\,
            lcout => \ALU.un1_yindexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_2_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__50497\,
            in1 => \N__49796\,
            in2 => \_gnd_net_\,
            in3 => \N__50443\,
            lcout => \yZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56246\,
            ce => \N__56053\,
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_2_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__50437\,
            in1 => \N__50485\,
            in2 => \N__49801\,
            in3 => \N__54956\,
            lcout => \ALU.un1_yindexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_3_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__54957\,
            in1 => \N__49787\,
            in2 => \N__50498\,
            in3 => \N__50438\,
            lcout => \ALU.un1_yindexZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_4_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__50439\,
            in1 => \N__50489\,
            in2 => \N__49802\,
            in3 => \N__54958\,
            lcout => \ALU.un1_yindexZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_5_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__54959\,
            in1 => \N__49791\,
            in2 => \N__50499\,
            in3 => \N__50440\,
            lcout => \ALU.un1_yindexZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_6_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__50441\,
            in1 => \N__50493\,
            in2 => \N__49803\,
            in3 => \N__54960\,
            lcout => \ALU.un1_yindexZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_7_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__54961\,
            in1 => \N__49795\,
            in2 => \N__50500\,
            in3 => \N__50442\,
            lcout => \ALU.un1_yindexZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNISU5D9_2_9_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52327\,
            in2 => \_gnd_net_\,
            in3 => \N__47470\,
            lcout => \ALU.r4_RNISU5D9_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_5_s1_c_RNO_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52879\,
            in2 => \_gnd_net_\,
            in3 => \N__47265\,
            lcout => \ALU.r0_12_prm_7_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_14_s1_c_RNO_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__54925\,
            in1 => \N__47148\,
            in2 => \N__53114\,
            in3 => \N__47066\,
            lcout => \ALU.r0_12_prm_5_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_7_s1_c_RNO_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52880\,
            in2 => \_gnd_net_\,
            in3 => \N__48076\,
            lcout => \ALU.r0_12_prm_7_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_1_c_RNO_0_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48653\,
            in2 => \_gnd_net_\,
            in3 => \N__46833\,
            lcout => \ALU.un14_log_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s1_c_RNO_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55506\,
            in2 => \_gnd_net_\,
            in3 => \N__47959\,
            lcout => \ALU.r0_12_prm_8_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_7_s0_c_RNO_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__48077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52893\,
            lcout => \ALU.r0_12_prm_7_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s1_c_RNO_0_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50560\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \ALU.r0_12_prm_8_14_s1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s1_c_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47986\,
            in2 => \N__47976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_14_s1_cy\,
            carryout => \ALU.r0_12_prm_8_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_14_s1_c_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47938\,
            in2 => \N__47929\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_14_s1\,
            carryout => \ALU.r0_12_prm_7_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_14_s1_c_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47908\,
            in2 => \N__47896\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_14_s1\,
            carryout => \ALU.r0_12_prm_6_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_14_s1_c_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47872\,
            in2 => \N__47859\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_14_s1\,
            carryout => \ALU.r0_12_prm_5_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_14_s1_c_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47842\,
            in2 => \N__47833\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_14_s1\,
            carryout => \ALU.r0_12_prm_4_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_14_s1_c_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55260\,
            in2 => \N__56507\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_14_s1\,
            carryout => \ALU.r0_12_prm_3_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_14_s1_c_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49141\,
            in2 => \N__49105\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_14_s1\,
            carryout => \ALU.r0_12_prm_2_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_14_s1_c_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49096\,
            in2 => \N__49084\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \ALU.r0_12_s1_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_s1_14_THRU_LUT4_0_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49036\,
            lcout => \ALU.r0_12_s1_14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \op_0_LC_16_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55641\,
            lcout => \opZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56226\,
            ce => \N__56059\,
            sr => \_gnd_net_\
        );

    \ALU.r4_RNIMVMDA_1_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__49016\,
            in1 => \N__54020\,
            in2 => \N__54889\,
            in3 => \N__48648\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNII2A0L_2_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__54828\,
            in1 => \N__48335\,
            in2 => \N__48169\,
            in3 => \N__49416\,
            lcout => \ALU.r4_RNII2A0LZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_5_s0_c_RNO_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__55434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48137\,
            lcout => \ALU.r0_12_prm_8_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r4_RNI0C236_9_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54021\,
            in1 => \N__54827\,
            in2 => \N__52972\,
            in3 => \N__52320\,
            lcout => \ALU.r4_RNI0C236Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \op_RNI705F_0_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__55585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => op_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_THRU_CRY_0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49545\,
            in2 => \N__49549\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_5_0_\,
            carryout => \ALU.r0_12_prm_8_3_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49534\,
            in2 => \N__50719\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_3_c_THRU_CO\,
            carryout => \ALU.r0_12_prm_8_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_3_c_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49522\,
            in2 => \N__49516\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_8_3\,
            carryout => \ALU.r0_12_prm_7_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_6_3_c_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49492\,
            in2 => \N__49480\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_7_3\,
            carryout => \ALU.r0_12_prm_6_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_5_3_c_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49465\,
            in2 => \N__49459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_6_3\,
            carryout => \ALU.r0_12_prm_5_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_3_c_inv_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49444\,
            in2 => \N__49153\,
            in3 => \N__49393\,
            lcout => \ALU.a_i_3\,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_5_3\,
            carryout => \ALU.r0_12_prm_4_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_3_c_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50068\,
            in2 => \N__50011\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_4_3\,
            carryout => \ALU.r0_12_prm_3_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_3_c_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50074\,
            in2 => \N__50110\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.r0_12_prm_3_3\,
            carryout => \ALU.r0_12_prm_2_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_1_3_c_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50242\,
            in2 => \N__50236\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_6_0_\,
            carryout => \ALU.r0_12_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_3_THRU_LUT4_0_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50203\,
            lcout => \ALU.r0_12_3_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_3_c_RNO_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55801\,
            in2 => \_gnd_net_\,
            in3 => \N__50103\,
            lcout => \ALU.r0_12_prm_2_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_3_3_c_RNO_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__55071\,
            in1 => \N__50031\,
            in2 => \_gnd_net_\,
            in3 => \N__50061\,
            lcout => \ALU.r0_12_prm_3_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_madd_cry_2_s_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__50062\,
            in1 => \_gnd_net_\,
            in2 => \N__50035\,
            in3 => \_gnd_net_\,
            lcout => \ALU.mult_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_0_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50466\,
            lcout => \yZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56229\,
            ce => \N__56055\,
            sr => \_gnd_net_\
        );

    \TXbuffer_7_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__50002\,
            in1 => \N__49987\,
            in2 => \N__49974\,
            in3 => \N__49816\,
            lcout => \TXbufferZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56229\,
            ce => \N__56055\,
            sr => \_gnd_net_\
        );

    \ALU.un1_yindex_8_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50411\,
            in1 => \N__50461\,
            in2 => \N__49807\,
            in3 => \N__54936\,
            lcout => \ALU.un1_yindexZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \y_1_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__50462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50412\,
            lcout => \yZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56231\,
            ce => \N__56054\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_7_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50398\,
            in2 => \_gnd_net_\,
            in3 => \N__56831\,
            lcout => \FTDI.TXshiftZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_7C_net\,
            ce => \N__56578\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_1_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50350\,
            in1 => \N__50389\,
            in2 => \_gnd_net_\,
            in3 => \N__56838\,
            lcout => \FTDI.TXshiftZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__56593\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_2_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50302\,
            in1 => \N__50371\,
            in2 => \_gnd_net_\,
            in3 => \N__56839\,
            lcout => \FTDI.TXshiftZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__56593\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_4_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50248\,
            in1 => \N__50344\,
            in2 => \_gnd_net_\,
            in3 => \N__56836\,
            lcout => \FTDI.TXshiftZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_4C_net\,
            ce => \N__56579\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_3_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56834\,
            in1 => \N__50326\,
            in2 => \_gnd_net_\,
            in3 => \N__50320\,
            lcout => \FTDI.TXshiftZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_4C_net\,
            ce => \N__56579\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_6_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50296\,
            in1 => \N__50287\,
            in2 => \_gnd_net_\,
            in3 => \N__56837\,
            lcout => \FTDI.TXshiftZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_4C_net\,
            ce => \N__56579\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_5_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56835\,
            in1 => \N__50272\,
            in2 => \_gnd_net_\,
            in3 => \N__50266\,
            lcout => \FTDI.TXshiftZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_4C_net\,
            ce => \N__56579\,
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_7_10_s0_c_RNO_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__52741\,
            in1 => \N__52036\,
            in2 => \_gnd_net_\,
            in3 => \N__51797\,
            lcout => \ALU.r0_12_prm_7_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_3_c_RNO_0_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51508\,
            in1 => \N__51098\,
            in2 => \_gnd_net_\,
            in3 => \N__50772\,
            lcout => \ALU.lshift_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_8_14_s1_c_RNO_1_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__50706\,
            in1 => \N__54890\,
            in2 => \_gnd_net_\,
            in3 => \N__50622\,
            lcout => \ALU.r0_12_prm_8_14_s1_c_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_2_1_c_RNO_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50554\,
            in2 => \_gnd_net_\,
            in3 => \N__50548\,
            lcout => \ALU.r0_12_prm_2_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \op_1_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55693\,
            in2 => \_gnd_net_\,
            in3 => \N__55072\,
            lcout => \opZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56228\,
            ce => \N__56058\,
            sr => \_gnd_net_\
        );

    \op_1_cry_1_c_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55142\,
            in2 => \N__55839\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => op_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \op_2_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52448\,
            in2 => \_gnd_net_\,
            in3 => \N__50509\,
            lcout => \opZ0Z_2\,
            ltout => OPEN,
            carryin => op_1_cry_1,
            carryout => op_1_cry_2,
            clk => \N__56232\,
            ce => \N__56056\,
            sr => \_gnd_net_\
        );

    \op_3_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55382\,
            in2 => \_gnd_net_\,
            in3 => \N__50506\,
            lcout => \opZ0Z_3\,
            ltout => OPEN,
            carryin => op_1_cry_2,
            carryout => op_1_cry_3,
            clk => \N__56232\,
            ce => \N__56056\,
            sr => \_gnd_net_\
        );

    \op_4_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54973\,
            in2 => \_gnd_net_\,
            in3 => \N__50503\,
            lcout => \opZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56232\,
            ce => \N__56056\,
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_1_1_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56896\,
            in2 => \_gnd_net_\,
            in3 => \N__56861\,
            lcout => OPEN,
            ltout => \FTDI.N_208_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_1_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__56799\,
            in1 => \N__56741\,
            in2 => \N__55981\,
            in3 => \N__56948\,
            lcout => \FTDI.N_207_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNICVLM_0_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56740\,
            lcout => \FTDI.N_185_0\,
            ltout => \FTDI.N_185_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_1_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001001000"
        )
    port map (
            in0 => \N__56949\,
            in1 => \N__56800\,
            in2 => \N__55978\,
            in3 => \N__55975\,
            lcout => \FTDI.TXstateZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_op_1_1_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55759\,
            in2 => \_gnd_net_\,
            in3 => \N__55381\,
            lcout => OPEN,
            ltout => \ALU.un1_op_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_op_1_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__55098\,
            in1 => \N__52447\,
            in2 => \N__54976\,
            in3 => \N__54972\,
            lcout => \ALU.un1_op_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.r0_12_prm_4_9_s1_c_RNO_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__54922\,
            in1 => \N__53972\,
            in2 => \N__52598\,
            in3 => \N__52325\,
            lcout => \ALU.r0_12_prm_4_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_2_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001110101111"
        )
    port map (
            in0 => \N__56742\,
            in1 => \N__56920\,
            in2 => \N__56904\,
            in3 => \N__56796\,
            lcout => OPEN,
            ltout => \FTDI.TXstate_cnst_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_2_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111100001111"
        )
    port map (
            in0 => \N__56641\,
            in1 => \_gnd_net_\,
            in2 => \N__56644\,
            in3 => \N__56695\,
            lcout => \FTDI.un3_TX_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_RNINKH42_2_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__56743\,
            in1 => \N__56795\,
            in2 => \N__56702\,
            in3 => \N__56640\,
            lcout => \FTDI.un1_TXstate_0_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_0_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__56617\,
            in1 => \N__56611\,
            in2 => \_gnd_net_\,
            in3 => \N__56810\,
            lcout => \FTDI.TXshiftZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_0C_net\,
            ce => \N__56586\,
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_2_c_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56323\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_6_0_\,
            carryout => \FTDI.un3_TX_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_3_c_inv_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__56833\,
            in1 => \N__56545\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \FTDI.un3_TX_axb_3\,
            ltout => OPEN,
            carryin => \FTDI.un3_TX_cry_2\,
            carryout => \FTDI.un3_TX_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__56539\,
            in1 => \N__56832\,
            in2 => \_gnd_net_\,
            in3 => \N__56527\,
            lcout => \FTDI_TX_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_2_c_inv_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__56322\,
            in1 => \N__56505\,
            in2 => \_gnd_net_\,
            in3 => \N__56905\,
            lcout => \FTDI.un3_TX_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_0_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000011"
        )
    port map (
            in0 => \N__56895\,
            in1 => \N__56311\,
            in2 => \N__56713\,
            in3 => \N__56947\,
            lcout => \FTDI.TXstateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNIEFF51_0_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__56946\,
            in1 => \N__56894\,
            in2 => \N__56816\,
            in3 => \N__56866\,
            lcout => \FTDI.TXready\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_3_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__56865\,
            in1 => \N__56739\,
            in2 => \_gnd_net_\,
            in3 => \N__56950\,
            lcout => \FTDI.TXstate_e_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNINQ101_0_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__56737\,
            in1 => \N__56945\,
            in2 => \_gnd_net_\,
            in3 => \N__56863\,
            lcout => \FTDI.N_186_0\,
            ltout => \FTDI.N_186_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_3_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111011001100"
        )
    port map (
            in0 => \N__56914\,
            in1 => \N__56798\,
            in2 => \N__56908\,
            in3 => \N__56900\,
            lcout => \FTDI.TXstateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_2_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__56656\,
            in1 => \N__56673\,
            in2 => \_gnd_net_\,
            in3 => \N__56701\,
            lcout => \FTDI.baudAccZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_0_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__56864\,
            in1 => \N__56797\,
            in2 => \_gnd_net_\,
            in3 => \N__56738\,
            lcout => \FTDI.TXstate_e_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_0_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__56704\,
            in1 => \N__56669\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \FTDI.baudAccZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_1_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56703\,
            in2 => \N__56674\,
            in3 => \N__56655\,
            lcout => \FTDI.baudAccZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
