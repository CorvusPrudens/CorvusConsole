-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Aug 14 2020 14:01:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    RX : in std_logic;
    GPIO3 : out std_logic;
    TX : out std_logic;
    GPIO2 : out std_logic;
    GPIO11 : out std_logic;
    GPIO0 : out std_logic;
    CLK : in std_logic;
    GPIO9 : out std_logic;
    GPIO1 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__16292\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \clkdivZ0Z_0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \clkdivZ0Z_1\ : std_logic;
signal clkdiv_cry_0 : std_logic;
signal \clkdivZ0Z_2\ : std_logic;
signal clkdiv_cry_1 : std_logic;
signal \clkdivZ0Z_3\ : std_logic;
signal clkdiv_cry_2 : std_logic;
signal \clkdivZ0Z_4\ : std_logic;
signal clkdiv_cry_3 : std_logic;
signal \clkdivZ0Z_5\ : std_logic;
signal clkdiv_cry_4 : std_logic;
signal \clkdivZ0Z_6\ : std_logic;
signal clkdiv_cry_5 : std_logic;
signal \clkdivZ0Z_7\ : std_logic;
signal clkdiv_cry_6 : std_logic;
signal clkdiv_cry_7 : std_logic;
signal \clkdivZ0Z_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \clkdivZ0Z_9\ : std_logic;
signal clkdiv_cry_8 : std_logic;
signal \clkdivZ0Z_10\ : std_logic;
signal clkdiv_cry_9 : std_logic;
signal \clkdivZ0Z_11\ : std_logic;
signal clkdiv_cry_10 : std_logic;
signal \clkdivZ0Z_12\ : std_logic;
signal clkdiv_cry_11 : std_logic;
signal \clkdivZ0Z_13\ : std_logic;
signal clkdiv_cry_12 : std_logic;
signal \clkdivZ0Z_14\ : std_logic;
signal clkdiv_cry_13 : std_logic;
signal \clkdivZ0Z_15\ : std_logic;
signal clkdiv_cry_14 : std_logic;
signal clkdiv_cry_15 : std_logic;
signal \clkdivZ0Z_16\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \clkdivZ0Z_17\ : std_logic;
signal clkdiv_cry_16 : std_logic;
signal \clkdivZ0Z_18\ : std_logic;
signal clkdiv_cry_17 : std_logic;
signal \clkdivZ0Z_19\ : std_logic;
signal clkdiv_cry_18 : std_logic;
signal \clkdivZ0Z_20\ : std_logic;
signal clkdiv_cry_19 : std_logic;
signal \clkdivZ0Z_21\ : std_logic;
signal clkdiv_cry_20 : std_logic;
signal \clkdivZ0Z_22\ : std_logic;
signal clkdiv_cry_21 : std_logic;
signal clkdiv_cry_22 : std_logic;
signal \GPIO3_c\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_2\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \ALU.regsA_result_cry_1\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \ALU.regsA_result_cry_4\ : std_logic;
signal \ALU.regsA_result_cry_5\ : std_logic;
signal \ALU.regsA_result_cry_6\ : std_logic;
signal \ALU.regsA_result_cry_7\ : std_logic;
signal \ALU.regsA_result_cry_4_c_RNO\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNIKGQO9\ : std_logic;
signal \FTDI.i2_mux_cascade_\ : std_logic;
signal \FTDI.TXstate_RNIE1MMZ0Z_2\ : std_logic;
signal \FTDI.TXstate_RNIE1MMZ0Z_2_cascade_\ : std_logic;
signal \INVFTDI.TXstate_0C_net\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_1\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \ALU.regsA_result_cry_2_ma_1\ : std_logic;
signal \ALU.regsA_result_cry_1_5\ : std_logic;
signal \ALU.regsA_result_cry_3_ma_1\ : std_logic;
signal \ALU.regsA_result_cry_2_7\ : std_logic;
signal \ALU.regsA_result_cry_4_ma_0\ : std_logic;
signal \ALU.regsA_result_cry_3_7\ : std_logic;
signal \ALU.regsA_result_cry_4_6\ : std_logic;
signal \ALU.regsA_result_cry_5_0\ : std_logic;
signal \ALU.regsA_result_axb_4_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_5_ma_0\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_704\ : std_logic;
signal \ALU.regsA_result_cry_2_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_705\ : std_logic;
signal \ALU.regsA_result_cry_3_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_706\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_871\ : std_logic;
signal \ALU.regsA_result_cry_4_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_707\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_872\ : std_logic;
signal \ALU.regsA_result_cry_5_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_708\ : std_logic;
signal \ALU.regsA_result_cry_6_3\ : std_logic;
signal \ALU.regsA_result_cry_7_1\ : std_logic;
signal \ALU.regsA_result_cry_2_c_RNO\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_873\ : std_logic;
signal \ALU.regsA_result_cry_2_c_RNIC59KA\ : std_logic;
signal \ALU.regsA_result_cry_2\ : std_logic;
signal \ALU.regsA_result_cry_3_0\ : std_logic;
signal \ALU.regsA_result_cry_3_0_THRU_CO\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_739\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_774\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_3\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_740\ : std_logic;
signal \ALU.regsA_result_cry_1_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_741\ : std_logic;
signal \ALU.regsA_result_cry_2_6\ : std_logic;
signal \ALU.regsA_result_axb_2\ : std_logic;
signal \ALU.regsA_result_cry_1_THRU_CO\ : std_logic;
signal \ALU.regsA_result_cry_3\ : std_logic;
signal \ALU.regsA_result_axb_4_0\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_axb_4\ : std_logic;
signal \FTDI.baudAccZ0Z_0\ : std_logic;
signal \FTDI.baudAccZ0Z_1\ : std_logic;
signal \INVFTDI.baudAcc_0C_net\ : std_logic;
signal \FTDI.N_170_0_cascade_\ : std_logic;
signal \FTDI.TXstate_cnst_0_0_2_cascade_\ : std_logic;
signal \INVFTDI.TXstate_2C_net\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_870\ : std_logic;
signal \FTDI.TXstateZ0Z_1\ : std_logic;
signal \FTDI.TXstate_fastZ0Z_3\ : std_logic;
signal \FTDI.TXstateZ0Z_0\ : std_logic;
signal \FTDI_TXready_cascade_\ : std_logic;
signal \un1_testState31_0_cascade_\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_669\ : std_logic;
signal \ALU.regsA_result_cry_0_0\ : std_logic;
signal \ALU.regsA_result_cry_5_c_RNI073QE\ : std_logic;
signal \ALU.regsA_result_cry_1_1\ : std_logic;
signal \ALU.regsA_result_cry_2_c_RNIHNOEF\ : std_logic;
signal \ALU.regsA_result_cry_2_2\ : std_logic;
signal \ALU.regsA_result_cry_7_c_RNI8EG3H\ : std_logic;
signal \ALU.regsA_result_cry_3_2\ : std_logic;
signal \ALU.regsA_result_cry_4_c_RNIA939H\ : std_logic;
signal \ALU.regsA_result_cry_4_1\ : std_logic;
signal \ALU.regsA_result_cry_5_c_RNIKCNNP\ : std_logic;
signal \ALU.regsA_result_cry_5_2\ : std_logic;
signal \ALU.regsA_result_cry_6_c_RNICICNO\ : std_logic;
signal \ALU.regsA_result_cry_6_1\ : std_logic;
signal \ALU.regsA_result_cry_7_9\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \a_fastZ0Z_10\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx_1\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx_1\ : std_logic;
signal \ALU.regsA_result_axb_5_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_1\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx_2\ : std_logic;
signal \ALU.regsA_result_cry_1_6\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx_2\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_671\ : std_logic;
signal \ALU.regsA_result_cry_2_8\ : std_logic;
signal \ALU.regsA_result_axb_4_l_ofx_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_672\ : std_logic;
signal \ALU.regsA_result_cry_3_8\ : std_logic;
signal \ALU.regsA_result_axb_5_l_ofx_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_673\ : std_logic;
signal \ALU.regsA_result_cry_4_7\ : std_logic;
signal \ALU.regsA_result_axb_6_l_ofx_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_674\ : std_logic;
signal \ALU.regsA_result_cry_5_7\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_675\ : std_logic;
signal \ALU.regsA_result_cry_6_6\ : std_logic;
signal \ALU.regsA_result_cry_5_0_THRU_CO\ : std_logic;
signal \ALU.regsA_result_cry_7_0\ : std_logic;
signal \ALU.regsA_result_axb_8_2\ : std_logic;
signal \ALU.regsA_result_cry_6_ma_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_670\ : std_logic;
signal \ALU.regsA_result_cry_2_c_RNO_0\ : std_logic;
signal \ALU.regsA_result_cry_3_ma_0\ : std_logic;
signal \ALU.regsA_result_axb_6\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_0\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \ALU.addsub_cry_0_c_THRU_CO\ : std_logic;
signal \ALU.addsub_cry_0\ : std_logic;
signal \ALU.addsub_axb_2_l_ofxZ0\ : std_logic;
signal \ALU.addsub_cry_1\ : std_logic;
signal \ALU.addsub_cry_2\ : std_logic;
signal \ALU.addsub_cry_3\ : std_logic;
signal \ALU.addsub_cry_4\ : std_logic;
signal \ALU.addsub_cry_5\ : std_logic;
signal \ALU.addsub_cry_6\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \ALU.addsub_cry_7\ : std_logic;
signal \ALU.addsub_cry_8\ : std_logic;
signal \aZ0Z_10\ : std_logic;
signal \ALU.addsub_axb_10_l_ofxZ0\ : std_logic;
signal \ALU.addsub_cry_9\ : std_logic;
signal \ALU.addsub_cry_10\ : std_logic;
signal \aZ0Z_12\ : std_logic;
signal \ALU.addsub_axb_12_l_ofxZ0\ : std_logic;
signal \ALU.addsub_cry_11\ : std_logic;
signal \ALU.addsub_cry_12\ : std_logic;
signal \ALU.addsub_cry_13\ : std_logic;
signal \ALU.addsub_cry_14\ : std_logic;
signal \aZ0Z_15\ : std_logic;
signal \ALU.addsub_axb_15_l_ofxZ0\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \ALU.mult_16\ : std_logic;
signal \ALU.addsub_cry_15\ : std_logic;
signal \ALU.addsub_14\ : std_logic;
signal \ALU.mult_14\ : std_logic;
signal \ALU.mult_ab_128\ : std_logic;
signal \ALU.addsub_8\ : std_logic;
signal res_8 : std_logic;
signal \ALU.addsub_11\ : std_logic;
signal \ALU.mult_11\ : std_logic;
signal \ALU.addsub_0\ : std_logic;
signal \GPIO0_c\ : std_logic;
signal \ALU.addsub_13\ : std_logic;
signal \ALU.mult_13\ : std_logic;
signal \ALU.addsub_12\ : std_logic;
signal \ALU.mult_12\ : std_logic;
signal \ALU.mult_1\ : std_logic;
signal \ALU.addsub_1\ : std_logic;
signal \ALU.addsub_9\ : std_logic;
signal \ALU.mult_9\ : std_logic;
signal \ALU.addsub_10\ : std_logic;
signal \ALU.mult_10\ : std_logic;
signal \ALU.addsub_15\ : std_logic;
signal \ALU.mult_15\ : std_logic;
signal \ALU.addsub_6\ : std_logic;
signal \ALU.mult_2_cascade_\ : std_logic;
signal \ALU.addsub_2\ : std_logic;
signal \ALU.regsA_result_cry_7_ma_0\ : std_logic;
signal \ALU.regsA_result_axb_7_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_axb_8_1\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_2\ : std_logic;
signal \ALU.regsA_result_cry_2_ma_2\ : std_logic;
signal \ALU.regsA_result_cry_3_ma_2\ : std_logic;
signal \ALU.regsA_result_cry_4_ma_1\ : std_logic;
signal \aZ0Z_14\ : std_logic;
signal \ALU.addsub_axb_14_l_ofxZ0\ : std_logic;
signal \aZ0Z_8\ : std_logic;
signal \ALU.addsub_axb_8_l_ofxZ0\ : std_logic;
signal \ALU.addsub_axb_9_l_ofxZ0\ : std_logic;
signal \aZ0Z_9\ : std_logic;
signal \ALU.regsA_result_cry_5_ma_1\ : std_logic;
signal \ALU.regsA_result_cry_0_0_c_RNO\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \ALU.regsA_result_axb_1_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_0_2\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_1_3\ : std_logic;
signal \ALU.regsA_result_cry_3_ma\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_2_5\ : std_logic;
signal \ALU.regsA_result_axb_4_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_3_6\ : std_logic;
signal \ALU.regsA_result_axb_5_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_4_5\ : std_logic;
signal \ALU.regsA_result_cry_5_6\ : std_logic;
signal \ALU.regsA_result_axb_7_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_6_5\ : std_logic;
signal \ALU.regsA_result_cry_7_5\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \ALU.regsA_result_cry_8_2\ : std_logic;
signal \ALU.regsA_result_cry_9_3\ : std_logic;
signal \ALU.regsA_result_cry_10_2\ : std_logic;
signal \ALU.regsA_result_cry_11_3\ : std_logic;
signal \ALU.regsA_result_cry_12_0\ : std_logic;
signal \ALU.regsA_result_cry_13_1\ : std_logic;
signal \ALU.regsA_result_cry_14\ : std_logic;
signal \ALU.regsA_result_axb_14_l_ofx\ : std_logic;
signal \ALU.addsub_axb_7_l_ofxZ0\ : std_logic;
signal \ALU.regsA_result_cry_8_ma\ : std_logic;
signal \ALU.regsA_result_axb_14_0\ : std_logic;
signal \ALU.regsA_result_cry_14_ma\ : std_logic;
signal \ALU.addsub_axb_1_l_ofxZ0\ : std_logic;
signal \bZ0Z_15\ : std_logic;
signal \ALU.overflow_RNOZ0Z_15\ : std_logic;
signal \ALU.addsub_axb_0_l_ofxZ0\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \ALU.regsA_result_cry_0\ : std_logic;
signal \ALU.mult_6\ : std_logic;
signal \ALU.regsA_result_cry_1_0\ : std_logic;
signal \ALU.regsA_result_cry_2_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_932\ : std_logic;
signal \ALU.regsA_result_cry_3_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_933\ : std_logic;
signal \ALU.regsA_result_cry_4_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_934\ : std_logic;
signal \ALU.regsA_result_cry_5_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_935\ : std_logic;
signal \ALU.regsA_result_cry_6_0\ : std_logic;
signal \ALU.regsA_result_cry_7_2\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_936\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_937\ : std_logic;
signal \ALU.regsA_result_cry_8\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_938\ : std_logic;
signal \ALU.regsA_result_cry_9_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_939\ : std_logic;
signal \ALU.regsA_result_cry_10\ : std_logic;
signal \ALU.regsA_result_axb_8\ : std_logic;
signal \ALU.regsA_result_cry_7_THRU_CO\ : std_logic;
signal \ALU.regsA_result_cry_11_0\ : std_logic;
signal \ALU.regsA_result_axb_8_0\ : std_logic;
signal \ALU.mult_5\ : std_logic;
signal \ALU.addsub_5\ : std_logic;
signal \ALU.addsub_7\ : std_logic;
signal \ALU.mult_7\ : std_logic;
signal overflow : std_logic;
signal \N_91\ : std_logic;
signal res_13 : std_logic;
signal res_5 : std_logic;
signal \GPIO2_c\ : std_logic;
signal res_10 : std_logic;
signal res_6 : std_logic;
signal res_14 : std_logic;
signal res_15 : std_logic;
signal res_7 : std_logic;
signal \aZ0Z_11\ : std_logic;
signal \ALU.addsub_axb_11_l_ofxZ0\ : std_logic;
signal \ALU.regsA_result_axb_12_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_11_ma\ : std_logic;
signal \ALU.regsA_result_cry_12_ma\ : std_logic;
signal \ALU.regsA_result_axb_13_l_ofx\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \ALU.regsA_result_cry_1_8\ : std_logic;
signal \ALU.regsA_result_cry_2_10\ : std_logic;
signal \ALU.regsA_result_cry_3_10\ : std_logic;
signal \ALU.regsA_result_cry_5_ma_3\ : std_logic;
signal \ALU.regsA_result_cry_4_9\ : std_logic;
signal \ALU.regsA_result_cry_5_9\ : std_logic;
signal \ALU.regsA_result_cry_6_8\ : std_logic;
signal \ALU.regsA_result_cry_7_7\ : std_logic;
signal \ALU.regsA_result_cry_8_4\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \ALU.regsA_result_cry_9_5\ : std_logic;
signal \ALU.regsA_result_cry_10_4\ : std_logic;
signal \ALU.regsA_result_cry_11_4\ : std_logic;
signal \ALU.regsA_result_cry_13_ma_0\ : std_logic;
signal \ALU.regsA_result_axb_13_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_12_1\ : std_logic;
signal \ALU.regsA_result_cry_13_0\ : std_logic;
signal \ALU.regsA_result_cry_13_0_THRU_CO\ : std_logic;
signal \ALU.regsA_result_cry_12_ma_0\ : std_logic;
signal \ALU.regsA_result_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_531\ : std_logic;
signal \ALU.regsA_result_cry_0_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_532\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_565\ : std_logic;
signal \ALU.regsA_result_cry_1_2\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_533\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_566\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_797\ : std_logic;
signal \ALU.regsA_result_cry_2_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_534\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_567\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_798\ : std_logic;
signal \ALU.regsA_result_cry_3_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_535\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_568\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_799\ : std_logic;
signal \ALU.regsA_result_cry_4_2\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_536\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_569\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_800\ : std_logic;
signal \ALU.regsA_result_cry_5_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_537\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_570\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_801\ : std_logic;
signal \ALU.regsA_result_cry_6_2\ : std_logic;
signal \ALU.regsA_result_cry_7_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_538\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_571\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_802\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_539\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_572\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_803\ : std_logic;
signal \ALU.regsA_result_cry_8_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_540\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_573\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_804\ : std_logic;
signal \ALU.regsA_result_cry_9_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_541\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_574\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_805\ : std_logic;
signal \ALU.regsA_result_cry_10_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_542\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_575\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_806\ : std_logic;
signal \ALU.regsA_result_cry_11_2\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_543\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_576\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_807\ : std_logic;
signal \ALU.regsA_result_cry_12\ : std_logic;
signal \ALU.regsA_result_axb_14\ : std_logic;
signal \ALU.regsA_result_cry_13\ : std_logic;
signal \ALU.regsA_result_axb_12_0\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_832\ : std_logic;
signal \ALU.regsA_result_cry_2_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_833\ : std_logic;
signal \ALU.regsA_result_cry_3_5\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_834\ : std_logic;
signal \ALU.regsA_result_cry_4_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_835\ : std_logic;
signal \ALU.regsA_result_cry_5_5\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_836\ : std_logic;
signal \ALU.regsA_result_cry_6_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_837\ : std_logic;
signal \ALU.regsA_result_cry_7_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_838\ : std_logic;
signal \ALU.regsA_result_cry_8_1\ : std_logic;
signal \ALU.regsA_result_cry_9_2\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_839\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_840\ : std_logic;
signal \ALU.regsA_result_cry_10_1\ : std_logic;
signal \ALU.regsA_result_cry_11\ : std_logic;
signal \ALU.regsA_result_cry_11_THRU_CO\ : std_logic;
signal \ALU.regsA_result_axb_10_l_ofx\ : std_logic;
signal \ALU.addsub_3\ : std_logic;
signal \ALU.mult_3\ : std_logic;
signal res_11 : std_logic;
signal res_3 : std_logic;
signal \GPIO1_c\ : std_logic;
signal res_9 : std_logic;
signal res_12 : std_logic;
signal \TXstate_fast_RNIP6NA1_3\ : std_logic;
signal \ALU.regsA_result_axb_11_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_10_ma\ : std_logic;
signal \ALU.regsA_result_axb_11_l_ofx_1\ : std_logic;
signal \bZ0Z_12\ : std_logic;
signal \ALU.regsA_result_axb_12_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_axb_10_l_ofx_1\ : std_logic;
signal \ALU.regsA_result_cry_11_ma_1\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx_4\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx_4\ : std_logic;
signal \ALU.regsA_result_axb_4_l_ofx_3\ : std_logic;
signal \ALU.regsA_result_axb_5_l_ofx_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_564\ : std_logic;
signal \a_fastZ0Z_2\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_4\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_5\ : std_logic;
signal \ALU.regsA_result_cry_2_ma_4\ : std_logic;
signal \ALU.regsA_result_cry_3_ma_4\ : std_logic;
signal \ALU.regsA_result_cry_4_ma_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_831\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_530\ : std_logic;
signal \a_2_repZ0Z1\ : std_logic;
signal \ALU.regsA_result_cry_0_c_RNO_0\ : std_logic;
signal \ALU.regsA_result_cry_4_ma\ : std_logic;
signal \ALU.regsA_result_cry_6_ma_2\ : std_logic;
signal \ALU.regsA_result_axb_6_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_5_ma\ : std_logic;
signal \ALU.regsA_result_axb_6_l_ofx_2\ : std_logic;
signal \ALU.regsA_result_cry_7_ma_2\ : std_logic;
signal \ALU.regsA_result_axb_7_l_ofx_2\ : std_logic;
signal \ALU.regsA_result_cry_6_ma\ : std_logic;
signal \ALU.regsA_result_cry_8_ma_1\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \ALU.regsA_result_cry_1_7\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_601\ : std_logic;
signal \ALU.regsA_result_cry_2_9\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_602\ : std_logic;
signal \ALU.regsA_result_cry_3_9\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_603\ : std_logic;
signal \ALU.regsA_result_cry_4_8\ : std_logic;
signal \ALU.regsA_result_axb_6_l_ofx_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_604\ : std_logic;
signal \ALU.regsA_result_cry_5_8\ : std_logic;
signal \ALU.regsA_result_axb_7_l_ofx_1\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_605\ : std_logic;
signal \ALU.regsA_result_cry_6_7\ : std_logic;
signal \ALU.regsA_result_axb_8_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_8_ma_0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_606\ : std_logic;
signal \ALU.regsA_result_cry_7_6\ : std_logic;
signal \ALU.regsA_result_cry_8_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_607\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_608\ : std_logic;
signal \ALU.regsA_result_cry_9_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_609\ : std_logic;
signal \ALU.regsA_result_cry_10_3\ : std_logic;
signal \ALU.regsA_result_axb_12_1\ : std_logic;
signal \ALU.regsA_result_cry_11_1\ : std_logic;
signal \ALU.regsA_result_axb_12\ : std_logic;
signal \ALU.regsA_result_axb_10_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_11_ma_0\ : std_logic;
signal \bZ0Z_11\ : std_logic;
signal \ALU.regsA_result_axb_11_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_10_ma_0\ : std_logic;
signal \TXbufferZ0Z_1\ : std_logic;
signal \TXbufferZ0Z_2\ : std_logic;
signal \FTDI.TXshiftZ0Z_2\ : std_logic;
signal \TXbufferZ0Z_6\ : std_logic;
signal \TXbufferZ0Z_4\ : std_logic;
signal \FTDI.TXshiftZ0Z_1\ : std_logic;
signal \TXbufferZ0Z_0\ : std_logic;
signal \FTDI.TXshiftZ0Z_4\ : std_logic;
signal \TXbufferZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_6\ : std_logic;
signal \TXbufferZ0Z_5\ : std_logic;
signal \FTDI.TXshiftZ0Z_5\ : std_logic;
signal \INVFTDI.TXshift_1C_net\ : std_logic;
signal \INVFTDI.RXbuffer_2C_net\ : std_logic;
signal \INVFTDI.RXbuffer_5C_net\ : std_logic;
signal \RXbuffer_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_599\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_3\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx_3\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx_3\ : std_logic;
signal \ALU.regsA_result_cry_0_c_RNO\ : std_logic;
signal \a_fastZ0Z_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_796\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_634\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_5\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \ALU.regsA_result_axb_2_l_ofx_5\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_635\ : std_logic;
signal \ALU.regsA_result_cry_1_9\ : std_logic;
signal \ALU.regsA_result_axb_3_l_ofx_5\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_636\ : std_logic;
signal \ALU.regsA_result_cry_2_11\ : std_logic;
signal \ALU.regsA_result_axb_4_l_ofx_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_637\ : std_logic;
signal \ALU.regsA_result_cry_3_11\ : std_logic;
signal \ALU.regsA_result_axb_5_l_ofx_4\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_638\ : std_logic;
signal \ALU.regsA_result_cry_4_10\ : std_logic;
signal \ALU.regsA_result_axb_6_l_ofx_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_639\ : std_logic;
signal \ALU.regsA_result_cry_5_10\ : std_logic;
signal \ALU.regsA_result_axb_7_l_ofx_3\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_640\ : std_logic;
signal \ALU.regsA_result_cry_6_9\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_641\ : std_logic;
signal \ALU.regsA_result_cry_7_8\ : std_logic;
signal \ALU.regsA_result_cry_8_5\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_642\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \ALU.regsA_result_cry_9\ : std_logic;
signal \ALU.regsA_result_cry_9_THRU_CO\ : std_logic;
signal \ALU.regsA_result_cry_9_ma_0\ : std_logic;
signal \ALU.regsA_result_cry_2_ma_3\ : std_logic;
signal \ALU.regsA_result_cry_7_ma_1\ : std_logic;
signal \ALU.regsA_result_axb_10\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_4\ : std_logic;
signal \ALU.regsA_result_cry_1_0_c_RNO_0_6\ : std_logic;
signal \ALU.regsA_result_axb_4_l_ofx_2\ : std_logic;
signal \RXbuffer_4\ : std_logic;
signal \ALU.regsA_result_axb_5_l_ofx_2\ : std_logic;
signal \ALU.addsub_axb_4_l_ofxZ0\ : std_logic;
signal \ALU.regsA_result_cry_4_ma_2\ : std_logic;
signal \ALU.regsA_result_cry_5_ma_2\ : std_logic;
signal \ALU.regsA_result_cry_6_ma_1\ : std_logic;
signal \ALU.regsA_result_axb_9_l_ofx\ : std_logic;
signal \aZ0Z_4\ : std_logic;
signal \ALU.regsA_result_axb_9_l_ofx_0\ : std_logic;
signal \ALU.regsA_result_cry_10_ma_1\ : std_logic;
signal \RXbuffer_2\ : std_logic;
signal \TXbufferZ0Z_7\ : std_logic;
signal \FTDI.TXshiftZ0Z_7\ : std_logic;
signal \INVFTDI.TXshift_7C_net\ : std_logic;
signal \RX_c\ : std_logic;
signal \FTDI.m13_ns_1_cascade_\ : std_logic;
signal \FTDI.N_201_2\ : std_logic;
signal \FTDI.N_23_cascade_\ : std_logic;
signal \FTDI.RXstateZ0Z_0\ : std_logic;
signal \INVFTDI.RXstate_3C_net\ : std_logic;
signal \FTDI.RXstateZ0Z_3\ : std_logic;
signal \FTDI.RXstateZ0Z_2\ : std_logic;
signal \FTDI.N_28\ : std_logic;
signal \FTDI.RXstateZ0Z_1\ : std_logic;
signal \INVFTDI.RXstate_2C_net\ : std_logic;
signal \RXready_RNIICV7_0\ : std_logic;
signal \RXbuffer_1\ : std_logic;
signal \opZ0Z_1\ : std_logic;
signal \ALU.addsub_4\ : std_logic;
signal \ALU.mult_4\ : std_logic;
signal res_4 : std_logic;
signal \ALU.regsA_result_cry_2_ma_0\ : std_logic;
signal \RXbuffer_5\ : std_logic;
signal \RXready_RNIICV7_1\ : std_logic;
signal \ALU.regsA_result_cry_1_ma\ : std_logic;
signal \ALU.regsA_result_cry_3_ma_3\ : std_logic;
signal \ALU.regsA_result_cry_2_ma\ : std_logic;
signal \RXbuffer_7\ : std_logic;
signal \bZ0Z_1\ : std_logic;
signal \ALU.regsA_result_cry_2_ma_5\ : std_logic;
signal \bZ0Z_2\ : std_logic;
signal \ALU.regsA_result_cry_3_ma_5\ : std_logic;
signal \ALU.regsA_result_cry_4_ma_4\ : std_logic;
signal \bZ0Z_4\ : std_logic;
signal \ALU.regsA_result_cry_5_ma_4\ : std_logic;
signal \ALU.regsA_result_cry_6_ma_3\ : std_logic;
signal \aZ0Z_1\ : std_logic;
signal \ALU.regsA_result_axb_8_l_ofx\ : std_logic;
signal \ALU.regsA_result_cry_7_ma\ : std_logic;
signal \ALU.regsA_result_axb_8_l_ofx_1\ : std_logic;
signal \ALU.regsA_result_cry_9_ma_1\ : std_logic;
signal \aZ0Z_2\ : std_logic;
signal \ALU.regsA_result_axb_9_l_ofx_1\ : std_logic;
signal \ALU.regsA_result_axb_8_l_ofx_2\ : std_logic;
signal \bZ0Z_9\ : std_logic;
signal \ALU.regsA_result_axb_9_l_ofx_2\ : std_logic;
signal \ALU.addsub_axb_6_l_ofxZ0\ : std_logic;
signal \ALU.mult_AdderTree2_bigtree_600\ : std_logic;
signal \aZ0Z_6\ : std_logic;
signal \bZ0Z_0\ : std_logic;
signal \ALU.regsA_result_cry_2_c_RNO_1\ : std_logic;
signal \aZ0Z_3\ : std_logic;
signal \bZ0Z_3\ : std_logic;
signal \ALU.addsub_axb_3_l_ofxZ0\ : std_logic;
signal \bZ0Z_8\ : std_logic;
signal \ALU.regsA_result_cry_9_ma_2\ : std_logic;
signal \bZ0Z_6\ : std_logic;
signal \ALU.regsA_result_cry_7_ma_3\ : std_logic;
signal \aZ0Z_7\ : std_logic;
signal \bZ0Z_7\ : std_logic;
signal \ALU.regsA_result_cry_8_ma_2\ : std_logic;
signal \FTDI.baudAccZ0Z_2\ : std_logic;
signal \FTDI.un1_TXstate_0_sqmuxa_0_i\ : std_logic;
signal \TXstartZ0\ : std_logic;
signal \un1_testState31_0_0\ : std_logic;
signal \bZ0Z_10\ : std_logic;
signal \ALU.regsA_result_cry_9_ma\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \FTDI.un3_TX_0\ : std_logic;
signal \FTDI.gap8\ : std_logic;
signal \FTDI.gapZ0Z_1\ : std_logic;
signal \FTDI.gapZ0Z_0\ : std_logic;
signal \FTDI.gapZ0Z_2\ : std_logic;
signal \INVFTDI.gap_1C_net\ : std_logic;
signal m7_x1 : std_logic;
signal \m7_x0_cascade_\ : std_logic;
signal \RXready_RNIICV7_2\ : std_logic;
signal \testState30_testState30_1_cascade_\ : std_logic;
signal \aZ0Z_5\ : std_logic;
signal \bZ0Z_5\ : std_logic;
signal \ALU.addsub_axb_5_l_ofxZ0\ : std_logic;
signal \aZ0Z_0\ : std_logic;
signal \ALU.regsA_result_cry_13_ma\ : std_logic;
signal \aZ0Z_13\ : std_logic;
signal \bZ0Z_13\ : std_logic;
signal \ALU.addsub_axb_13_l_ofxZ0\ : std_logic;
signal \RXbuffer_0\ : std_logic;
signal \opZ0Z_0\ : std_logic;
signal \RXbuffer_6\ : std_logic;
signal \bZ0Z_14\ : std_logic;
signal \RXready_RNIICV7\ : std_logic;
signal \i3_mux_i_x0_cascade_\ : std_logic;
signal \FTDI_TXready\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \testState27\ : std_logic;
signal \testStateZ0Z_0\ : std_logic;
signal \testStateZ0Z_2\ : std_logic;
signal \testStateZ0Z_1\ : std_logic;
signal \RXready\ : std_logic;
signal i3_mux_i_x1 : std_logic;
signal \FTDI.un3_TX_0_i\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \FTDI.un3_TX_axb_3\ : std_logic;
signal \FTDI.un3_TX_cry_2\ : std_logic;
signal \FTDI.TXstateZ0Z_3\ : std_logic;
signal \FTDI.TXshiftZ0Z_0\ : std_logic;
signal \FTDI.un3_TX_cry_3\ : std_logic;
signal \FTDI_TX_0_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \GPIO1_wire\ : std_logic;
signal \GPIO3_wire\ : std_logic;
signal \GPIO0_wire\ : std_logic;
signal \GPIO2_wire\ : std_logic;
signal \RX_wire\ : std_logic;
signal \GPIO11_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \GPIO9_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    GPIO1 <= \GPIO1_wire\;
    GPIO3 <= \GPIO3_wire\;
    GPIO0 <= \GPIO0_wire\;
    GPIO2 <= \GPIO2_wire\;
    \RX_wire\ <= RX;
    GPIO11 <= \GPIO11_wire\;
    TX <= \TX_wire\;
    GPIO9 <= \GPIO9_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__16290\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16292\,
            DIN => \N__16291\,
            DOUT => \N__16290\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__16292\,
            PADOUT => \N__16291\,
            PADIN => \N__16290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16281\,
            DIN => \N__16280\,
            DOUT => \N__16279\,
            PACKAGEPIN => \GPIO1_wire\
        );

    \GPIO1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16281\,
            PADOUT => \N__16280\,
            PADIN => \N__16279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9440\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16272\,
            DIN => \N__16271\,
            DOUT => \N__16270\,
            PACKAGEPIN => \GPIO3_wire\
        );

    \GPIO3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16272\,
            PADOUT => \N__16271\,
            PADIN => \N__16270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6281\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16263\,
            DIN => \N__16262\,
            DOUT => \N__16261\,
            PACKAGEPIN => \GPIO0_wire\
        );

    \GPIO0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16263\,
            PADOUT => \N__16262\,
            PADIN => \N__16261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7550\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16254\,
            DIN => \N__16253\,
            DOUT => \N__16252\,
            PACKAGEPIN => \GPIO2_wire\
        );

    \GPIO2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16254\,
            PADOUT => \N__16253\,
            PADIN => \N__16252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8456\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RX_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16245\,
            DIN => \N__16244\,
            DOUT => \N__16243\,
            PACKAGEPIN => \RX_wire\
        );

    \RX_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__16245\,
            PADOUT => \N__16244\,
            PADIN => \N__16243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO11_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16236\,
            DIN => \N__16235\,
            DOUT => \N__16234\,
            PACKAGEPIN => \GPIO11_wire\
        );

    \GPIO11_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16236\,
            PADOUT => \N__16235\,
            PADIN => \N__16234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TX_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16227\,
            DIN => \N__16226\,
            DOUT => \N__16225\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16227\,
            PADOUT => \N__16226\,
            PADIN => \N__16225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15326\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO9_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16218\,
            DIN => \N__16217\,
            DOUT => \N__16216\,
            PACKAGEPIN => \GPIO9_wire\
        );

    \GPIO9_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16218\,
            PADOUT => \N__16217\,
            PADIN => \N__16216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14056\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__16199\,
            I => \i3_mux_i_x0_cascade_\
        );

    \I__3891\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16192\
        );

    \I__3890\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16189\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__16192\,
            I => \N__16182\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__16189\,
            I => \N__16179\
        );

    \I__3887\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16176\
        );

    \I__3886\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16169\
        );

    \I__3885\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16164\
        );

    \I__3884\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16164\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__16182\,
            I => \N__16161\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__16179\,
            I => \N__16158\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__16176\,
            I => \N__16155\
        );

    \I__3880\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16148\
        );

    \I__3879\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16148\
        );

    \I__3878\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16148\
        );

    \I__3877\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16145\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__16169\,
            I => \N__16140\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__16164\,
            I => \N__16140\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__16161\,
            I => \N__16133\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__16158\,
            I => \N__16133\
        );

    \I__3872\ : Span4Mux_v
    port map (
            O => \N__16155\,
            I => \N__16133\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__16148\,
            I => \FTDI_TXready\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__16145\,
            I => \FTDI_TXready\
        );

    \I__3869\ : Odrv12
    port map (
            O => \N__16140\,
            I => \FTDI_TXready\
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__16133\,
            I => \FTDI_TXready\
        );

    \I__3867\ : ClkMux
    port map (
            O => \N__16124\,
            I => \N__15968\
        );

    \I__3866\ : ClkMux
    port map (
            O => \N__16123\,
            I => \N__15968\
        );

    \I__3865\ : ClkMux
    port map (
            O => \N__16122\,
            I => \N__15968\
        );

    \I__3864\ : ClkMux
    port map (
            O => \N__16121\,
            I => \N__15968\
        );

    \I__3863\ : ClkMux
    port map (
            O => \N__16120\,
            I => \N__15968\
        );

    \I__3862\ : ClkMux
    port map (
            O => \N__16119\,
            I => \N__15968\
        );

    \I__3861\ : ClkMux
    port map (
            O => \N__16118\,
            I => \N__15968\
        );

    \I__3860\ : ClkMux
    port map (
            O => \N__16117\,
            I => \N__15968\
        );

    \I__3859\ : ClkMux
    port map (
            O => \N__16116\,
            I => \N__15968\
        );

    \I__3858\ : ClkMux
    port map (
            O => \N__16115\,
            I => \N__15968\
        );

    \I__3857\ : ClkMux
    port map (
            O => \N__16114\,
            I => \N__15968\
        );

    \I__3856\ : ClkMux
    port map (
            O => \N__16113\,
            I => \N__15968\
        );

    \I__3855\ : ClkMux
    port map (
            O => \N__16112\,
            I => \N__15968\
        );

    \I__3854\ : ClkMux
    port map (
            O => \N__16111\,
            I => \N__15968\
        );

    \I__3853\ : ClkMux
    port map (
            O => \N__16110\,
            I => \N__15968\
        );

    \I__3852\ : ClkMux
    port map (
            O => \N__16109\,
            I => \N__15968\
        );

    \I__3851\ : ClkMux
    port map (
            O => \N__16108\,
            I => \N__15968\
        );

    \I__3850\ : ClkMux
    port map (
            O => \N__16107\,
            I => \N__15968\
        );

    \I__3849\ : ClkMux
    port map (
            O => \N__16106\,
            I => \N__15968\
        );

    \I__3848\ : ClkMux
    port map (
            O => \N__16105\,
            I => \N__15968\
        );

    \I__3847\ : ClkMux
    port map (
            O => \N__16104\,
            I => \N__15968\
        );

    \I__3846\ : ClkMux
    port map (
            O => \N__16103\,
            I => \N__15968\
        );

    \I__3845\ : ClkMux
    port map (
            O => \N__16102\,
            I => \N__15968\
        );

    \I__3844\ : ClkMux
    port map (
            O => \N__16101\,
            I => \N__15968\
        );

    \I__3843\ : ClkMux
    port map (
            O => \N__16100\,
            I => \N__15968\
        );

    \I__3842\ : ClkMux
    port map (
            O => \N__16099\,
            I => \N__15968\
        );

    \I__3841\ : ClkMux
    port map (
            O => \N__16098\,
            I => \N__15968\
        );

    \I__3840\ : ClkMux
    port map (
            O => \N__16097\,
            I => \N__15968\
        );

    \I__3839\ : ClkMux
    port map (
            O => \N__16096\,
            I => \N__15968\
        );

    \I__3838\ : ClkMux
    port map (
            O => \N__16095\,
            I => \N__15968\
        );

    \I__3837\ : ClkMux
    port map (
            O => \N__16094\,
            I => \N__15968\
        );

    \I__3836\ : ClkMux
    port map (
            O => \N__16093\,
            I => \N__15968\
        );

    \I__3835\ : ClkMux
    port map (
            O => \N__16092\,
            I => \N__15968\
        );

    \I__3834\ : ClkMux
    port map (
            O => \N__16091\,
            I => \N__15968\
        );

    \I__3833\ : ClkMux
    port map (
            O => \N__16090\,
            I => \N__15968\
        );

    \I__3832\ : ClkMux
    port map (
            O => \N__16089\,
            I => \N__15968\
        );

    \I__3831\ : ClkMux
    port map (
            O => \N__16088\,
            I => \N__15968\
        );

    \I__3830\ : ClkMux
    port map (
            O => \N__16087\,
            I => \N__15968\
        );

    \I__3829\ : ClkMux
    port map (
            O => \N__16086\,
            I => \N__15968\
        );

    \I__3828\ : ClkMux
    port map (
            O => \N__16085\,
            I => \N__15968\
        );

    \I__3827\ : ClkMux
    port map (
            O => \N__16084\,
            I => \N__15968\
        );

    \I__3826\ : ClkMux
    port map (
            O => \N__16083\,
            I => \N__15968\
        );

    \I__3825\ : ClkMux
    port map (
            O => \N__16082\,
            I => \N__15968\
        );

    \I__3824\ : ClkMux
    port map (
            O => \N__16081\,
            I => \N__15968\
        );

    \I__3823\ : ClkMux
    port map (
            O => \N__16080\,
            I => \N__15968\
        );

    \I__3822\ : ClkMux
    port map (
            O => \N__16079\,
            I => \N__15968\
        );

    \I__3821\ : ClkMux
    port map (
            O => \N__16078\,
            I => \N__15968\
        );

    \I__3820\ : ClkMux
    port map (
            O => \N__16077\,
            I => \N__15968\
        );

    \I__3819\ : ClkMux
    port map (
            O => \N__16076\,
            I => \N__15968\
        );

    \I__3818\ : ClkMux
    port map (
            O => \N__16075\,
            I => \N__15968\
        );

    \I__3817\ : ClkMux
    port map (
            O => \N__16074\,
            I => \N__15968\
        );

    \I__3816\ : ClkMux
    port map (
            O => \N__16073\,
            I => \N__15968\
        );

    \I__3815\ : GlobalMux
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__3814\ : gio2CtrlBuf
    port map (
            O => \N__15965\,
            I => \CLK_c_g\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__15962\,
            I => \N__15958\
        );

    \I__3812\ : SRMux
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__3811\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15951\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15948\
        );

    \I__3809\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15944\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__15951\,
            I => \N__15941\
        );

    \I__3807\ : Span4Mux_h
    port map (
            O => \N__15948\,
            I => \N__15938\
        );

    \I__3806\ : InMux
    port map (
            O => \N__15947\,
            I => \N__15935\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__15944\,
            I => \N__15932\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__15941\,
            I => \N__15929\
        );

    \I__3803\ : Span4Mux_h
    port map (
            O => \N__15938\,
            I => \N__15926\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__15935\,
            I => \N__15923\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__15932\,
            I => \testState27\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__15929\,
            I => \testState27\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__15926\,
            I => \testState27\
        );

    \I__3798\ : Odrv12
    port map (
            O => \N__15923\,
            I => \testState27\
        );

    \I__3797\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15903\
        );

    \I__3796\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15895\
        );

    \I__3795\ : InMux
    port map (
            O => \N__15912\,
            I => \N__15895\
        );

    \I__3794\ : InMux
    port map (
            O => \N__15911\,
            I => \N__15895\
        );

    \I__3793\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15884\
        );

    \I__3792\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15884\
        );

    \I__3791\ : InMux
    port map (
            O => \N__15908\,
            I => \N__15884\
        );

    \I__3790\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15884\
        );

    \I__3789\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15884\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__15903\,
            I => \N__15876\
        );

    \I__3787\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15873\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__15895\,
            I => \N__15867\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15867\
        );

    \I__3784\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15864\
        );

    \I__3783\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15861\
        );

    \I__3782\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15858\
        );

    \I__3781\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15855\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__15879\,
            I => \N__15850\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__15876\,
            I => \N__15844\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__15873\,
            I => \N__15844\
        );

    \I__3777\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15841\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__15867\,
            I => \N__15836\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__15864\,
            I => \N__15836\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__15861\,
            I => \N__15829\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__15858\,
            I => \N__15829\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__15855\,
            I => \N__15829\
        );

    \I__3771\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15819\
        );

    \I__3770\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15819\
        );

    \I__3769\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15819\
        );

    \I__3768\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15816\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__15844\,
            I => \N__15813\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__15841\,
            I => \N__15806\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__15836\,
            I => \N__15806\
        );

    \I__3764\ : Span4Mux_v
    port map (
            O => \N__15829\,
            I => \N__15806\
        );

    \I__3763\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15799\
        );

    \I__3762\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15799\
        );

    \I__3761\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15799\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__15819\,
            I => \N__15796\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__15816\,
            I => \testStateZ0Z_0\
        );

    \I__3758\ : Odrv4
    port map (
            O => \N__15813\,
            I => \testStateZ0Z_0\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__15806\,
            I => \testStateZ0Z_0\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__15799\,
            I => \testStateZ0Z_0\
        );

    \I__3755\ : Odrv12
    port map (
            O => \N__15796\,
            I => \testStateZ0Z_0\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__15785\,
            I => \N__15779\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__15784\,
            I => \N__15775\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__15783\,
            I => \N__15772\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__15782\,
            I => \N__15769\
        );

    \I__3750\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15765\
        );

    \I__3749\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15762\
        );

    \I__3748\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15757\
        );

    \I__3747\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15754\
        );

    \I__3746\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15751\
        );

    \I__3745\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15748\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__15765\,
            I => \N__15745\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__15762\,
            I => \N__15742\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__15761\,
            I => \N__15739\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__15760\,
            I => \N__15736\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__15757\,
            I => \N__15724\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15724\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15724\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15717\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__15745\,
            I => \N__15717\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__15742\,
            I => \N__15717\
        );

    \I__3734\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15710\
        );

    \I__3733\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15710\
        );

    \I__3732\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15710\
        );

    \I__3731\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15703\
        );

    \I__3730\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15703\
        );

    \I__3729\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15703\
        );

    \I__3728\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15700\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__15724\,
            I => \N__15695\
        );

    \I__3726\ : Span4Mux_h
    port map (
            O => \N__15717\,
            I => \N__15695\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__15710\,
            I => \N__15692\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__15703\,
            I => \N__15689\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__15700\,
            I => \testStateZ0Z_2\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__15695\,
            I => \testStateZ0Z_2\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__15692\,
            I => \testStateZ0Z_2\
        );

    \I__3720\ : Odrv12
    port map (
            O => \N__15689\,
            I => \testStateZ0Z_2\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__15680\,
            I => \N__15671\
        );

    \I__3718\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15666\
        );

    \I__3717\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15666\
        );

    \I__3716\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15663\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__15676\,
            I => \N__15658\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__15675\,
            I => \N__15655\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__15674\,
            I => \N__15652\
        );

    \I__3712\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15647\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__15666\,
            I => \N__15640\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__15663\,
            I => \N__15640\
        );

    \I__3709\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15637\
        );

    \I__3708\ : InMux
    port map (
            O => \N__15661\,
            I => \N__15634\
        );

    \I__3707\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15625\
        );

    \I__3706\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15625\
        );

    \I__3705\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15625\
        );

    \I__3704\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15625\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__15650\,
            I => \N__15622\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15619\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__15646\,
            I => \N__15616\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__15645\,
            I => \N__15613\
        );

    \I__3699\ : Span4Mux_v
    port map (
            O => \N__15640\,
            I => \N__15607\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__15637\,
            I => \N__15607\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15602\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__15625\,
            I => \N__15598\
        );

    \I__3695\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15595\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__15619\,
            I => \N__15592\
        );

    \I__3693\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15585\
        );

    \I__3692\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15585\
        );

    \I__3691\ : InMux
    port map (
            O => \N__15612\,
            I => \N__15585\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__15607\,
            I => \N__15581\
        );

    \I__3689\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15578\
        );

    \I__3688\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15575\
        );

    \I__3687\ : Span4Mux_v
    port map (
            O => \N__15602\,
            I => \N__15569\
        );

    \I__3686\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15566\
        );

    \I__3685\ : Span4Mux_v
    port map (
            O => \N__15598\,
            I => \N__15563\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15556\
        );

    \I__3683\ : Span4Mux_h
    port map (
            O => \N__15592\,
            I => \N__15556\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__15585\,
            I => \N__15556\
        );

    \I__3681\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15553\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__15581\,
            I => \N__15546\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__15578\,
            I => \N__15546\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__15575\,
            I => \N__15546\
        );

    \I__3677\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15539\
        );

    \I__3676\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15539\
        );

    \I__3675\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15539\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__15569\,
            I => \N__15536\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__15566\,
            I => \N__15529\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__15563\,
            I => \N__15529\
        );

    \I__3671\ : Span4Mux_v
    port map (
            O => \N__15556\,
            I => \N__15529\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__15553\,
            I => \testStateZ0Z_1\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__15546\,
            I => \testStateZ0Z_1\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__15539\,
            I => \testStateZ0Z_1\
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__15536\,
            I => \testStateZ0Z_1\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__15529\,
            I => \testStateZ0Z_1\
        );

    \I__3665\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15510\
        );

    \I__3664\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15510\
        );

    \I__3663\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15505\
        );

    \I__3662\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15505\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__15510\,
            I => \N__15493\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__15505\,
            I => \N__15493\
        );

    \I__3659\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15486\
        );

    \I__3658\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15486\
        );

    \I__3657\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15486\
        );

    \I__3656\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15483\
        );

    \I__3655\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15478\
        );

    \I__3654\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15478\
        );

    \I__3653\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15475\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__15493\,
            I => \N__15470\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__15486\,
            I => \N__15470\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__15483\,
            I => \RXready\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__15478\,
            I => \RXready\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__15475\,
            I => \RXready\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__15470\,
            I => \RXready\
        );

    \I__3646\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__15458\,
            I => i3_mux_i_x1
        );

    \I__3644\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15451\
        );

    \I__3643\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15448\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__15451\,
            I => \FTDI.un3_TX_0_i\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__15448\,
            I => \FTDI.un3_TX_0_i\
        );

    \I__3640\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__15440\,
            I => \FTDI.un3_TX_axb_3\
        );

    \I__3638\ : InMux
    port map (
            O => \N__15437\,
            I => \N__15430\
        );

    \I__3637\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__15435\,
            I => \N__15419\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__15430\,
            I => \N__15416\
        );

    \I__3634\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15401\
        );

    \I__3633\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15401\
        );

    \I__3632\ : InMux
    port map (
            O => \N__15427\,
            I => \N__15401\
        );

    \I__3631\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15401\
        );

    \I__3630\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15401\
        );

    \I__3629\ : InMux
    port map (
            O => \N__15424\,
            I => \N__15401\
        );

    \I__3628\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15401\
        );

    \I__3627\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15398\
        );

    \I__3626\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15395\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__15416\,
            I => \N__15390\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__15401\,
            I => \N__15390\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__15398\,
            I => \N__15385\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__15395\,
            I => \N__15382\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__15390\,
            I => \N__15378\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__15389\,
            I => \N__15374\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__15388\,
            I => \N__15371\
        );

    \I__3618\ : Span4Mux_v
    port map (
            O => \N__15385\,
            I => \N__15366\
        );

    \I__3617\ : Span4Mux_h
    port map (
            O => \N__15382\,
            I => \N__15366\
        );

    \I__3616\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15363\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__15378\,
            I => \N__15360\
        );

    \I__3614\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15353\
        );

    \I__3613\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15353\
        );

    \I__3612\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15353\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__15366\,
            I => \N__15348\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__15363\,
            I => \N__15348\
        );

    \I__3609\ : Odrv4
    port map (
            O => \N__15360\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__15353\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__15348\,
            I => \FTDI.TXstateZ0Z_3\
        );

    \I__3606\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__15338\,
            I => \N__15335\
        );

    \I__3604\ : Span4Mux_v
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__15332\,
            I => \FTDI.TXshiftZ0Z_0\
        );

    \I__3602\ : InMux
    port map (
            O => \N__15329\,
            I => \FTDI.un3_TX_cry_3\
        );

    \I__3601\ : IoInMux
    port map (
            O => \N__15326\,
            I => \N__15323\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__3599\ : Span4Mux_s1_v
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__3598\ : Sp12to4
    port map (
            O => \N__15317\,
            I => \N__15314\
        );

    \I__3597\ : Span12Mux_h
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__3596\ : Span12Mux_v
    port map (
            O => \N__15311\,
            I => \N__15308\
        );

    \I__3595\ : Odrv12
    port map (
            O => \N__15308\,
            I => \FTDI_TX_0_i\
        );

    \I__3594\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__15302\,
            I => m7_x1
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__15299\,
            I => \m7_x0_cascade_\
        );

    \I__3591\ : CEMux
    port map (
            O => \N__15296\,
            I => \N__15292\
        );

    \I__3590\ : CEMux
    port map (
            O => \N__15295\,
            I => \N__15289\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__15292\,
            I => \N__15286\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15282\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__15286\,
            I => \N__15279\
        );

    \I__3586\ : CEMux
    port map (
            O => \N__15285\,
            I => \N__15276\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__15282\,
            I => \N__15270\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__15279\,
            I => \N__15265\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__15276\,
            I => \N__15265\
        );

    \I__3582\ : CEMux
    port map (
            O => \N__15275\,
            I => \N__15261\
        );

    \I__3581\ : CEMux
    port map (
            O => \N__15274\,
            I => \N__15258\
        );

    \I__3580\ : CEMux
    port map (
            O => \N__15273\,
            I => \N__15255\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__15270\,
            I => \N__15250\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__15265\,
            I => \N__15250\
        );

    \I__3577\ : CEMux
    port map (
            O => \N__15264\,
            I => \N__15246\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__15261\,
            I => \N__15243\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__15258\,
            I => \N__15238\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__15255\,
            I => \N__15238\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__15250\,
            I => \N__15235\
        );

    \I__3572\ : CEMux
    port map (
            O => \N__15249\,
            I => \N__15232\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15246\,
            I => \N__15229\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__15243\,
            I => \N__15224\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__15238\,
            I => \N__15224\
        );

    \I__3568\ : Sp12to4
    port map (
            O => \N__15235\,
            I => \N__15217\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__15232\,
            I => \N__15217\
        );

    \I__3566\ : Sp12to4
    port map (
            O => \N__15229\,
            I => \N__15217\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__15224\,
            I => \N__15214\
        );

    \I__3564\ : Odrv12
    port map (
            O => \N__15217\,
            I => \RXready_RNIICV7_2\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__15214\,
            I => \RXready_RNIICV7_2\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \testState30_testState30_1_cascade_\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__15206\,
            I => \N__15201\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__15205\,
            I => \N__15196\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15192\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15201\,
            I => \N__15183\
        );

    \I__3557\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15183\
        );

    \I__3556\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15174\
        );

    \I__3555\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15174\
        );

    \I__3554\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15171\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__15192\,
            I => \N__15168\
        );

    \I__3552\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15165\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__15190\,
            I => \N__15162\
        );

    \I__3550\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15156\
        );

    \I__3549\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15153\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__15183\,
            I => \N__15150\
        );

    \I__3547\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15143\
        );

    \I__3546\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15143\
        );

    \I__3545\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15143\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__15179\,
            I => \N__15139\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__15174\,
            I => \N__15129\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__15171\,
            I => \N__15126\
        );

    \I__3541\ : Span4Mux_v
    port map (
            O => \N__15168\,
            I => \N__15123\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__15165\,
            I => \N__15120\
        );

    \I__3539\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15117\
        );

    \I__3538\ : InMux
    port map (
            O => \N__15161\,
            I => \N__15110\
        );

    \I__3537\ : InMux
    port map (
            O => \N__15160\,
            I => \N__15110\
        );

    \I__3536\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15110\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15107\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__15153\,
            I => \N__15100\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__15150\,
            I => \N__15100\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__15143\,
            I => \N__15100\
        );

    \I__3531\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15088\
        );

    \I__3530\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15088\
        );

    \I__3529\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15088\
        );

    \I__3528\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15088\
        );

    \I__3527\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15088\
        );

    \I__3526\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15079\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15079\
        );

    \I__3524\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15079\
        );

    \I__3523\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15079\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__15129\,
            I => \N__15076\
        );

    \I__3521\ : Span4Mux_v
    port map (
            O => \N__15126\,
            I => \N__15071\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__15123\,
            I => \N__15071\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__15120\,
            I => \N__15060\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__15117\,
            I => \N__15060\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__15110\,
            I => \N__15060\
        );

    \I__3516\ : Span4Mux_v
    port map (
            O => \N__15107\,
            I => \N__15060\
        );

    \I__3515\ : Span4Mux_v
    port map (
            O => \N__15100\,
            I => \N__15060\
        );

    \I__3514\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15057\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__15088\,
            I => \N__15052\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__15079\,
            I => \N__15052\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__15076\,
            I => \aZ0Z_5\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__15071\,
            I => \aZ0Z_5\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__15060\,
            I => \aZ0Z_5\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__15057\,
            I => \aZ0Z_5\
        );

    \I__3507\ : Odrv12
    port map (
            O => \N__15052\,
            I => \aZ0Z_5\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__15041\,
            I => \N__15033\
        );

    \I__3505\ : InMux
    port map (
            O => \N__15040\,
            I => \N__15028\
        );

    \I__3504\ : InMux
    port map (
            O => \N__15039\,
            I => \N__15025\
        );

    \I__3503\ : InMux
    port map (
            O => \N__15038\,
            I => \N__15019\
        );

    \I__3502\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15019\
        );

    \I__3501\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15014\
        );

    \I__3500\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15011\
        );

    \I__3499\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15006\
        );

    \I__3498\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15006\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__15028\,
            I => \N__15002\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__15025\,
            I => \N__14995\
        );

    \I__3495\ : InMux
    port map (
            O => \N__15024\,
            I => \N__14992\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__15019\,
            I => \N__14989\
        );

    \I__3493\ : InMux
    port map (
            O => \N__15018\,
            I => \N__14982\
        );

    \I__3492\ : InMux
    port map (
            O => \N__15017\,
            I => \N__14982\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__15014\,
            I => \N__14979\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15011\,
            I => \N__14976\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__15006\,
            I => \N__14973\
        );

    \I__3488\ : InMux
    port map (
            O => \N__15005\,
            I => \N__14970\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__15002\,
            I => \N__14967\
        );

    \I__3486\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14962\
        );

    \I__3485\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14962\
        );

    \I__3484\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14957\
        );

    \I__3483\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14957\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__14995\,
            I => \N__14950\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__14992\,
            I => \N__14950\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__14989\,
            I => \N__14950\
        );

    \I__3479\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14945\
        );

    \I__3478\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14945\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__14982\,
            I => \N__14942\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__14979\,
            I => \N__14933\
        );

    \I__3475\ : Span4Mux_h
    port map (
            O => \N__14976\,
            I => \N__14933\
        );

    \I__3474\ : Span4Mux_h
    port map (
            O => \N__14973\,
            I => \N__14933\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__14970\,
            I => \N__14933\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__14967\,
            I => \bZ0Z_5\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__14962\,
            I => \bZ0Z_5\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__14957\,
            I => \bZ0Z_5\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__14950\,
            I => \bZ0Z_5\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__14945\,
            I => \bZ0Z_5\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__14942\,
            I => \bZ0Z_5\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__14933\,
            I => \bZ0Z_5\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__3464\ : InMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__3461\ : Span4Mux_h
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__14903\,
            I => \ALU.addsub_axb_5_l_ofxZ0\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \N__14894\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__14899\,
            I => \N__14891\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__14898\,
            I => \N__14882\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__14897\,
            I => \N__14879\
        );

    \I__3455\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14869\
        );

    \I__3454\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14869\
        );

    \I__3453\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14863\
        );

    \I__3452\ : InMux
    port map (
            O => \N__14889\,
            I => \N__14857\
        );

    \I__3451\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14848\
        );

    \I__3450\ : InMux
    port map (
            O => \N__14887\,
            I => \N__14848\
        );

    \I__3449\ : InMux
    port map (
            O => \N__14886\,
            I => \N__14848\
        );

    \I__3448\ : InMux
    port map (
            O => \N__14885\,
            I => \N__14848\
        );

    \I__3447\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14842\
        );

    \I__3446\ : InMux
    port map (
            O => \N__14879\,
            I => \N__14842\
        );

    \I__3445\ : InMux
    port map (
            O => \N__14878\,
            I => \N__14833\
        );

    \I__3444\ : InMux
    port map (
            O => \N__14877\,
            I => \N__14833\
        );

    \I__3443\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14833\
        );

    \I__3442\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14828\
        );

    \I__3441\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14825\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14822\
        );

    \I__3439\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14816\
        );

    \I__3438\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14811\
        );

    \I__3437\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14811\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__14863\,
            I => \N__14808\
        );

    \I__3435\ : InMux
    port map (
            O => \N__14862\,
            I => \N__14801\
        );

    \I__3434\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14801\
        );

    \I__3433\ : InMux
    port map (
            O => \N__14860\,
            I => \N__14801\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14796\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__14848\,
            I => \N__14796\
        );

    \I__3430\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14793\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__14842\,
            I => \N__14790\
        );

    \I__3428\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14785\
        );

    \I__3427\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14785\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__14833\,
            I => \N__14782\
        );

    \I__3425\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14777\
        );

    \I__3424\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14777\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14770\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14770\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__14822\,
            I => \N__14770\
        );

    \I__3420\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14767\
        );

    \I__3419\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14764\
        );

    \I__3418\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14761\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__14816\,
            I => \N__14758\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__14811\,
            I => \N__14755\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__14808\,
            I => \N__14747\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__14801\,
            I => \N__14747\
        );

    \I__3413\ : Span4Mux_h
    port map (
            O => \N__14796\,
            I => \N__14742\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__14793\,
            I => \N__14742\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__14790\,
            I => \N__14737\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__14785\,
            I => \N__14734\
        );

    \I__3409\ : Span4Mux_h
    port map (
            O => \N__14782\,
            I => \N__14729\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__14777\,
            I => \N__14729\
        );

    \I__3407\ : Span4Mux_h
    port map (
            O => \N__14770\,
            I => \N__14724\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__14767\,
            I => \N__14724\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__14764\,
            I => \N__14717\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__14761\,
            I => \N__14717\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__14758\,
            I => \N__14717\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__14755\,
            I => \N__14714\
        );

    \I__3401\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14711\
        );

    \I__3400\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14706\
        );

    \I__3399\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14706\
        );

    \I__3398\ : Span4Mux_h
    port map (
            O => \N__14747\,
            I => \N__14701\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__14742\,
            I => \N__14701\
        );

    \I__3396\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14696\
        );

    \I__3395\ : InMux
    port map (
            O => \N__14740\,
            I => \N__14696\
        );

    \I__3394\ : Span4Mux_h
    port map (
            O => \N__14737\,
            I => \N__14689\
        );

    \I__3393\ : Span4Mux_h
    port map (
            O => \N__14734\,
            I => \N__14689\
        );

    \I__3392\ : Span4Mux_h
    port map (
            O => \N__14729\,
            I => \N__14689\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__14724\,
            I => \N__14684\
        );

    \I__3390\ : Span4Mux_h
    port map (
            O => \N__14717\,
            I => \N__14684\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__14714\,
            I => \aZ0Z_0\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__14711\,
            I => \aZ0Z_0\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__14706\,
            I => \aZ0Z_0\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__14701\,
            I => \aZ0Z_0\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__14696\,
            I => \aZ0Z_0\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__14689\,
            I => \aZ0Z_0\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__14684\,
            I => \aZ0Z_0\
        );

    \I__3382\ : InMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__3380\ : Odrv12
    port map (
            O => \N__14663\,
            I => \ALU.regsA_result_cry_13_ma\
        );

    \I__3379\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14652\
        );

    \I__3378\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14649\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__14658\,
            I => \N__14645\
        );

    \I__3376\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14641\
        );

    \I__3375\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14636\
        );

    \I__3374\ : InMux
    port map (
            O => \N__14655\,
            I => \N__14636\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__14652\,
            I => \N__14631\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__14649\,
            I => \N__14631\
        );

    \I__3371\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14628\
        );

    \I__3370\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14623\
        );

    \I__3369\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14623\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14617\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__14636\,
            I => \N__14617\
        );

    \I__3366\ : Span4Mux_v
    port map (
            O => \N__14631\,
            I => \N__14610\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__14628\,
            I => \N__14610\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__14623\,
            I => \N__14610\
        );

    \I__3363\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14607\
        );

    \I__3362\ : Span4Mux_v
    port map (
            O => \N__14617\,
            I => \N__14604\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__14610\,
            I => \N__14600\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__14607\,
            I => \N__14597\
        );

    \I__3359\ : Span4Mux_h
    port map (
            O => \N__14604\,
            I => \N__14594\
        );

    \I__3358\ : InMux
    port map (
            O => \N__14603\,
            I => \N__14591\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__14600\,
            I => \N__14588\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__14597\,
            I => \aZ0Z_13\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__14594\,
            I => \aZ0Z_13\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__14591\,
            I => \aZ0Z_13\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__14588\,
            I => \aZ0Z_13\
        );

    \I__3352\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14575\
        );

    \I__3351\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14572\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__14575\,
            I => \N__14567\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__14572\,
            I => \N__14564\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__14571\,
            I => \N__14561\
        );

    \I__3347\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14556\
        );

    \I__3346\ : Span4Mux_h
    port map (
            O => \N__14567\,
            I => \N__14553\
        );

    \I__3345\ : Span4Mux_v
    port map (
            O => \N__14564\,
            I => \N__14550\
        );

    \I__3344\ : InMux
    port map (
            O => \N__14561\,
            I => \N__14543\
        );

    \I__3343\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14543\
        );

    \I__3342\ : InMux
    port map (
            O => \N__14559\,
            I => \N__14543\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__14556\,
            I => \bZ0Z_13\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__14553\,
            I => \bZ0Z_13\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__14550\,
            I => \bZ0Z_13\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__14543\,
            I => \bZ0Z_13\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__14534\,
            I => \N__14531\
        );

    \I__3336\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14528\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__3334\ : Span4Mux_h
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__14519\,
            I => \ALU.addsub_axb_13_l_ofxZ0\
        );

    \I__3331\ : InMux
    port map (
            O => \N__14516\,
            I => \N__14511\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__14515\,
            I => \N__14507\
        );

    \I__3329\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14504\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__14511\,
            I => \N__14500\
        );

    \I__3327\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14497\
        );

    \I__3326\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14494\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__14504\,
            I => \N__14491\
        );

    \I__3324\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14488\
        );

    \I__3323\ : Span4Mux_h
    port map (
            O => \N__14500\,
            I => \N__14481\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__14497\,
            I => \N__14481\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__14494\,
            I => \N__14481\
        );

    \I__3320\ : Span4Mux_h
    port map (
            O => \N__14491\,
            I => \N__14478\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14475\
        );

    \I__3318\ : Span4Mux_v
    port map (
            O => \N__14481\,
            I => \N__14472\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__14478\,
            I => \RXbuffer_0\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__14475\,
            I => \RXbuffer_0\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__14472\,
            I => \RXbuffer_0\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14460\
        );

    \I__3313\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14452\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__14463\,
            I => \N__14449\
        );

    \I__3311\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14440\
        );

    \I__3310\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14437\
        );

    \I__3309\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14434\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14427\
        );

    \I__3307\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14427\
        );

    \I__3306\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14427\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__14452\,
            I => \N__14423\
        );

    \I__3304\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14420\
        );

    \I__3303\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14417\
        );

    \I__3302\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14412\
        );

    \I__3301\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14412\
        );

    \I__3300\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14405\
        );

    \I__3299\ : InMux
    port map (
            O => \N__14444\,
            I => \N__14405\
        );

    \I__3298\ : InMux
    port map (
            O => \N__14443\,
            I => \N__14405\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__14440\,
            I => \N__14402\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14399\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14396\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__14427\,
            I => \N__14393\
        );

    \I__3293\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14390\
        );

    \I__3292\ : Span4Mux_v
    port map (
            O => \N__14423\,
            I => \N__14379\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__14420\,
            I => \N__14379\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__14417\,
            I => \N__14379\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__14412\,
            I => \N__14379\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__14405\,
            I => \N__14379\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__14402\,
            I => \N__14376\
        );

    \I__3286\ : Span4Mux_h
    port map (
            O => \N__14399\,
            I => \N__14373\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__14396\,
            I => \N__14363\
        );

    \I__3284\ : Span4Mux_h
    port map (
            O => \N__14393\,
            I => \N__14363\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__14390\,
            I => \N__14360\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__14379\,
            I => \N__14357\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__14376\,
            I => \N__14352\
        );

    \I__3280\ : Span4Mux_h
    port map (
            O => \N__14373\,
            I => \N__14352\
        );

    \I__3279\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14349\
        );

    \I__3278\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14346\
        );

    \I__3277\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14339\
        );

    \I__3276\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14339\
        );

    \I__3275\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14339\
        );

    \I__3274\ : Span4Mux_h
    port map (
            O => \N__14363\,
            I => \N__14334\
        );

    \I__3273\ : Span4Mux_h
    port map (
            O => \N__14360\,
            I => \N__14334\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__14357\,
            I => \N__14331\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__14352\,
            I => \opZ0Z_0\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__14349\,
            I => \opZ0Z_0\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__14346\,
            I => \opZ0Z_0\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__14339\,
            I => \opZ0Z_0\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__14334\,
            I => \opZ0Z_0\
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__14331\,
            I => \opZ0Z_0\
        );

    \I__3265\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14314\
        );

    \I__3264\ : InMux
    port map (
            O => \N__14317\,
            I => \N__14311\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__14311\,
            I => \N__14304\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__14308\,
            I => \N__14301\
        );

    \I__3260\ : InMux
    port map (
            O => \N__14307\,
            I => \N__14298\
        );

    \I__3259\ : Span4Mux_v
    port map (
            O => \N__14304\,
            I => \N__14293\
        );

    \I__3258\ : Span4Mux_h
    port map (
            O => \N__14301\,
            I => \N__14288\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14288\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14285\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14282\
        );

    \I__3254\ : Span4Mux_v
    port map (
            O => \N__14293\,
            I => \N__14277\
        );

    \I__3253\ : Span4Mux_v
    port map (
            O => \N__14288\,
            I => \N__14277\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__14285\,
            I => \N__14274\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__14282\,
            I => \RXbuffer_6\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__14277\,
            I => \RXbuffer_6\
        );

    \I__3249\ : Odrv4
    port map (
            O => \N__14274\,
            I => \RXbuffer_6\
        );

    \I__3248\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14263\
        );

    \I__3247\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14260\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__14260\,
            I => \N__14252\
        );

    \I__3244\ : Span4Mux_v
    port map (
            O => \N__14257\,
            I => \N__14249\
        );

    \I__3243\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14244\
        );

    \I__3242\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14244\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__14252\,
            I => \N__14240\
        );

    \I__3240\ : Sp12to4
    port map (
            O => \N__14249\,
            I => \N__14235\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__14244\,
            I => \N__14235\
        );

    \I__3238\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14232\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__14240\,
            I => \bZ0Z_14\
        );

    \I__3236\ : Odrv12
    port map (
            O => \N__14235\,
            I => \bZ0Z_14\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__14232\,
            I => \bZ0Z_14\
        );

    \I__3234\ : CEMux
    port map (
            O => \N__14225\,
            I => \N__14220\
        );

    \I__3233\ : CEMux
    port map (
            O => \N__14224\,
            I => \N__14216\
        );

    \I__3232\ : CEMux
    port map (
            O => \N__14223\,
            I => \N__14212\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__14220\,
            I => \N__14209\
        );

    \I__3230\ : CEMux
    port map (
            O => \N__14219\,
            I => \N__14206\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__14216\,
            I => \N__14203\
        );

    \I__3228\ : CEMux
    port map (
            O => \N__14215\,
            I => \N__14200\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__14212\,
            I => \N__14196\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__14209\,
            I => \N__14193\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14190\
        );

    \I__3224\ : Span4Mux_h
    port map (
            O => \N__14203\,
            I => \N__14185\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__14200\,
            I => \N__14185\
        );

    \I__3222\ : CEMux
    port map (
            O => \N__14199\,
            I => \N__14182\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__14196\,
            I => \N__14179\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__14193\,
            I => \N__14172\
        );

    \I__3219\ : Span4Mux_v
    port map (
            O => \N__14190\,
            I => \N__14172\
        );

    \I__3218\ : Span4Mux_v
    port map (
            O => \N__14185\,
            I => \N__14172\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__14182\,
            I => \N__14169\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__14179\,
            I => \RXready_RNIICV7\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__14172\,
            I => \RXready_RNIICV7\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__14169\,
            I => \RXready_RNIICV7\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__14162\,
            I => \N__14158\
        );

    \I__3212\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14154\
        );

    \I__3211\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14150\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__14157\,
            I => \N__14145\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__14154\,
            I => \N__14142\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__14153\,
            I => \N__14139\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__14150\,
            I => \N__14136\
        );

    \I__3206\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14131\
        );

    \I__3205\ : InMux
    port map (
            O => \N__14148\,
            I => \N__14131\
        );

    \I__3204\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14124\
        );

    \I__3203\ : Span4Mux_v
    port map (
            O => \N__14142\,
            I => \N__14121\
        );

    \I__3202\ : InMux
    port map (
            O => \N__14139\,
            I => \N__14118\
        );

    \I__3201\ : Span4Mux_h
    port map (
            O => \N__14136\,
            I => \N__14113\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__14131\,
            I => \N__14113\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14109\
        );

    \I__3198\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14102\
        );

    \I__3197\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14102\
        );

    \I__3196\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14102\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__14124\,
            I => \N__14099\
        );

    \I__3194\ : Span4Mux_h
    port map (
            O => \N__14121\,
            I => \N__14092\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__14118\,
            I => \N__14092\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__14113\,
            I => \N__14092\
        );

    \I__3191\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14089\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__14109\,
            I => \bZ0Z_10\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__14102\,
            I => \bZ0Z_10\
        );

    \I__3188\ : Odrv4
    port map (
            O => \N__14099\,
            I => \bZ0Z_10\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__14092\,
            I => \bZ0Z_10\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__14089\,
            I => \bZ0Z_10\
        );

    \I__3185\ : InMux
    port map (
            O => \N__14078\,
            I => \N__14075\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__14075\,
            I => \N__14072\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__14072\,
            I => \N__14069\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__14069\,
            I => \N__14066\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__14066\,
            I => \ALU.regsA_result_cry_9_ma\
        );

    \I__3180\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__14060\,
            I => \N__14057\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__14057\,
            I => \N__14053\
        );

    \I__3177\ : IoInMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__3176\ : Span4Mux_h
    port map (
            O => \N__14053\,
            I => \N__14047\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__14050\,
            I => \N__14044\
        );

    \I__3174\ : Sp12to4
    port map (
            O => \N__14047\,
            I => \N__14041\
        );

    \I__3173\ : IoSpan4Mux
    port map (
            O => \N__14044\,
            I => \N__14038\
        );

    \I__3172\ : Span12Mux_v
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__3171\ : Span4Mux_s2_v
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__3170\ : Odrv12
    port map (
            O => \N__14035\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__14032\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3168\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14024\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__3166\ : Span12Mux_v
    port map (
            O => \N__14021\,
            I => \N__14014\
        );

    \I__3165\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14011\
        );

    \I__3164\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14008\
        );

    \I__3163\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14003\
        );

    \I__3162\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14003\
        );

    \I__3161\ : Odrv12
    port map (
            O => \N__14014\,
            I => \FTDI.un3_TX_0\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__14011\,
            I => \FTDI.un3_TX_0\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__14008\,
            I => \FTDI.un3_TX_0\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__14003\,
            I => \FTDI.un3_TX_0\
        );

    \I__3157\ : InMux
    port map (
            O => \N__13994\,
            I => \N__13985\
        );

    \I__3156\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13985\
        );

    \I__3155\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13985\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__13985\,
            I => \FTDI.gap8\
        );

    \I__3153\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13976\
        );

    \I__3152\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13976\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__13976\,
            I => \FTDI.gapZ0Z_1\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__3149\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13961\
        );

    \I__3148\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13961\
        );

    \I__3147\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13961\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__13961\,
            I => \FTDI.gapZ0Z_0\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__13958\,
            I => \N__13953\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__13957\,
            I => \N__13947\
        );

    \I__3143\ : InMux
    port map (
            O => \N__13956\,
            I => \N__13938\
        );

    \I__3142\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13938\
        );

    \I__3141\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13938\
        );

    \I__3140\ : InMux
    port map (
            O => \N__13951\,
            I => \N__13938\
        );

    \I__3139\ : InMux
    port map (
            O => \N__13950\,
            I => \N__13933\
        );

    \I__3138\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13933\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__13938\,
            I => \FTDI.gapZ0Z_2\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__13933\,
            I => \FTDI.gapZ0Z_2\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__3134\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__3132\ : Span4Mux_h
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__13916\,
            I => \ALU.addsub_axb_6_l_ofxZ0\
        );

    \I__3130\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__3128\ : Span4Mux_v
    port map (
            O => \N__13907\,
            I => \N__13902\
        );

    \I__3127\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13899\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__13905\,
            I => \N__13896\
        );

    \I__3125\ : Span4Mux_v
    port map (
            O => \N__13902\,
            I => \N__13893\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__13899\,
            I => \N__13890\
        );

    \I__3123\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13887\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__13893\,
            I => \ALU.mult_AdderTree2_bigtree_600\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__13890\,
            I => \ALU.mult_AdderTree2_bigtree_600\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__13887\,
            I => \ALU.mult_AdderTree2_bigtree_600\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__13880\,
            I => \N__13875\
        );

    \I__3118\ : InMux
    port map (
            O => \N__13879\,
            I => \N__13870\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__13878\,
            I => \N__13860\
        );

    \I__3116\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13855\
        );

    \I__3115\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13855\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__13873\,
            I => \N__13852\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__13870\,
            I => \N__13849\
        );

    \I__3112\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13846\
        );

    \I__3111\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13843\
        );

    \I__3110\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13840\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__13866\,
            I => \N__13837\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__13865\,
            I => \N__13833\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__13864\,
            I => \N__13829\
        );

    \I__3106\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13823\
        );

    \I__3105\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13823\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__13855\,
            I => \N__13820\
        );

    \I__3103\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13817\
        );

    \I__3102\ : Span4Mux_h
    port map (
            O => \N__13849\,
            I => \N__13808\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__13846\,
            I => \N__13808\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__13843\,
            I => \N__13808\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__13840\,
            I => \N__13808\
        );

    \I__3098\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13795\
        );

    \I__3097\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13795\
        );

    \I__3096\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13795\
        );

    \I__3095\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13795\
        );

    \I__3094\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13795\
        );

    \I__3093\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13795\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__13823\,
            I => \aZ0Z_6\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__13820\,
            I => \aZ0Z_6\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__13817\,
            I => \aZ0Z_6\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__13808\,
            I => \aZ0Z_6\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__13795\,
            I => \aZ0Z_6\
        );

    \I__3087\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13777\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__13783\,
            I => \N__13773\
        );

    \I__3085\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13762\
        );

    \I__3084\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13759\
        );

    \I__3083\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13756\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__13777\,
            I => \N__13752\
        );

    \I__3081\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13749\
        );

    \I__3080\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13745\
        );

    \I__3079\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13741\
        );

    \I__3078\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13736\
        );

    \I__3077\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13736\
        );

    \I__3076\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13729\
        );

    \I__3075\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13729\
        );

    \I__3074\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13729\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__13766\,
            I => \N__13718\
        );

    \I__3072\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13713\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__13762\,
            I => \N__13710\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__13759\,
            I => \N__13705\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__13756\,
            I => \N__13705\
        );

    \I__3068\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13702\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__13752\,
            I => \N__13697\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__13749\,
            I => \N__13697\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13694\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__13745\,
            I => \N__13691\
        );

    \I__3063\ : InMux
    port map (
            O => \N__13744\,
            I => \N__13688\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13683\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__13736\,
            I => \N__13683\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__13729\,
            I => \N__13680\
        );

    \I__3059\ : InMux
    port map (
            O => \N__13728\,
            I => \N__13677\
        );

    \I__3058\ : InMux
    port map (
            O => \N__13727\,
            I => \N__13664\
        );

    \I__3057\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13664\
        );

    \I__3056\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13657\
        );

    \I__3055\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13657\
        );

    \I__3054\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13657\
        );

    \I__3053\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13652\
        );

    \I__3052\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13652\
        );

    \I__3051\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13645\
        );

    \I__3050\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13645\
        );

    \I__3049\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13645\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__13713\,
            I => \N__13639\
        );

    \I__3047\ : Span4Mux_h
    port map (
            O => \N__13710\,
            I => \N__13632\
        );

    \I__3046\ : Span4Mux_v
    port map (
            O => \N__13705\,
            I => \N__13632\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__13702\,
            I => \N__13632\
        );

    \I__3044\ : Span4Mux_h
    port map (
            O => \N__13697\,
            I => \N__13627\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__13694\,
            I => \N__13627\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__13691\,
            I => \N__13616\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__13688\,
            I => \N__13616\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__13683\,
            I => \N__13616\
        );

    \I__3039\ : Span4Mux_v
    port map (
            O => \N__13680\,
            I => \N__13616\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__13677\,
            I => \N__13616\
        );

    \I__3037\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13611\
        );

    \I__3036\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13611\
        );

    \I__3035\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13602\
        );

    \I__3034\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13602\
        );

    \I__3033\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13602\
        );

    \I__3032\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13602\
        );

    \I__3031\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13597\
        );

    \I__3030\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13597\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__13664\,
            I => \N__13594\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__13657\,
            I => \N__13587\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13587\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__13645\,
            I => \N__13587\
        );

    \I__3025\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13582\
        );

    \I__3024\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13582\
        );

    \I__3023\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13579\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__13639\,
            I => \N__13574\
        );

    \I__3021\ : Span4Mux_h
    port map (
            O => \N__13632\,
            I => \N__13574\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__13627\,
            I => \N__13567\
        );

    \I__3019\ : Span4Mux_h
    port map (
            O => \N__13616\,
            I => \N__13567\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__13611\,
            I => \N__13567\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__13602\,
            I => \bZ0Z_0\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__13597\,
            I => \bZ0Z_0\
        );

    \I__3015\ : Odrv12
    port map (
            O => \N__13594\,
            I => \bZ0Z_0\
        );

    \I__3014\ : Odrv12
    port map (
            O => \N__13587\,
            I => \bZ0Z_0\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__13582\,
            I => \bZ0Z_0\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__13579\,
            I => \bZ0Z_0\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__13574\,
            I => \bZ0Z_0\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__13567\,
            I => \bZ0Z_0\
        );

    \I__3009\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__13541\,
            I => \ALU.regsA_result_cry_2_c_RNO_1\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__13538\,
            I => \N__13530\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__13537\,
            I => \N__13527\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__13536\,
            I => \N__13524\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__13535\,
            I => \N__13516\
        );

    \I__3001\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13509\
        );

    \I__3000\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13506\
        );

    \I__2999\ : InMux
    port map (
            O => \N__13530\,
            I => \N__13499\
        );

    \I__2998\ : InMux
    port map (
            O => \N__13527\,
            I => \N__13499\
        );

    \I__2997\ : InMux
    port map (
            O => \N__13524\,
            I => \N__13499\
        );

    \I__2996\ : InMux
    port map (
            O => \N__13523\,
            I => \N__13496\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__13522\,
            I => \N__13492\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__13521\,
            I => \N__13489\
        );

    \I__2993\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13485\
        );

    \I__2992\ : InMux
    port map (
            O => \N__13519\,
            I => \N__13482\
        );

    \I__2991\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13475\
        );

    \I__2990\ : InMux
    port map (
            O => \N__13515\,
            I => \N__13475\
        );

    \I__2989\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13475\
        );

    \I__2988\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13472\
        );

    \I__2987\ : InMux
    port map (
            O => \N__13512\,
            I => \N__13469\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__13509\,
            I => \N__13460\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__13506\,
            I => \N__13457\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__13499\,
            I => \N__13454\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13496\,
            I => \N__13451\
        );

    \I__2982\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13448\
        );

    \I__2981\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13441\
        );

    \I__2980\ : InMux
    port map (
            O => \N__13489\,
            I => \N__13441\
        );

    \I__2979\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13441\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__13485\,
            I => \N__13431\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13428\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__13475\,
            I => \N__13425\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__13472\,
            I => \N__13422\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__13469\,
            I => \N__13419\
        );

    \I__2973\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13416\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13411\
        );

    \I__2971\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13411\
        );

    \I__2970\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13404\
        );

    \I__2969\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13404\
        );

    \I__2968\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13404\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__13460\,
            I => \N__13401\
        );

    \I__2966\ : Span4Mux_v
    port map (
            O => \N__13457\,
            I => \N__13390\
        );

    \I__2965\ : Span4Mux_h
    port map (
            O => \N__13454\,
            I => \N__13390\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__13451\,
            I => \N__13390\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13390\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__13441\,
            I => \N__13390\
        );

    \I__2961\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13377\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13377\
        );

    \I__2959\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13377\
        );

    \I__2958\ : InMux
    port map (
            O => \N__13437\,
            I => \N__13377\
        );

    \I__2957\ : InMux
    port map (
            O => \N__13436\,
            I => \N__13377\
        );

    \I__2956\ : InMux
    port map (
            O => \N__13435\,
            I => \N__13377\
        );

    \I__2955\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13374\
        );

    \I__2954\ : Span4Mux_v
    port map (
            O => \N__13431\,
            I => \N__13365\
        );

    \I__2953\ : Span4Mux_v
    port map (
            O => \N__13428\,
            I => \N__13365\
        );

    \I__2952\ : Span4Mux_v
    port map (
            O => \N__13425\,
            I => \N__13365\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__13422\,
            I => \N__13365\
        );

    \I__2950\ : Odrv12
    port map (
            O => \N__13419\,
            I => \aZ0Z_3\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__13416\,
            I => \aZ0Z_3\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__13411\,
            I => \aZ0Z_3\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__13404\,
            I => \aZ0Z_3\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__13401\,
            I => \aZ0Z_3\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__13390\,
            I => \aZ0Z_3\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__13377\,
            I => \aZ0Z_3\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__13374\,
            I => \aZ0Z_3\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__13365\,
            I => \aZ0Z_3\
        );

    \I__2941\ : InMux
    port map (
            O => \N__13346\,
            I => \N__13339\
        );

    \I__2940\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13335\
        );

    \I__2939\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13331\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13326\
        );

    \I__2937\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13326\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__13339\,
            I => \N__13322\
        );

    \I__2935\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13319\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__13335\,
            I => \N__13312\
        );

    \I__2933\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13309\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__13331\,
            I => \N__13306\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__13326\,
            I => \N__13303\
        );

    \I__2930\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13300\
        );

    \I__2929\ : Span4Mux_v
    port map (
            O => \N__13322\,
            I => \N__13291\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__13319\,
            I => \N__13291\
        );

    \I__2927\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13288\
        );

    \I__2926\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13282\
        );

    \I__2925\ : InMux
    port map (
            O => \N__13316\,
            I => \N__13277\
        );

    \I__2924\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13277\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__13312\,
            I => \N__13270\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13270\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__13306\,
            I => \N__13270\
        );

    \I__2920\ : Span4Mux_h
    port map (
            O => \N__13303\,
            I => \N__13265\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__13300\,
            I => \N__13265\
        );

    \I__2918\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13261\
        );

    \I__2917\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13256\
        );

    \I__2916\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13256\
        );

    \I__2915\ : InMux
    port map (
            O => \N__13296\,
            I => \N__13253\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__13291\,
            I => \N__13247\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__13288\,
            I => \N__13247\
        );

    \I__2912\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13244\
        );

    \I__2911\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13239\
        );

    \I__2910\ : InMux
    port map (
            O => \N__13285\,
            I => \N__13239\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__13282\,
            I => \N__13234\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__13277\,
            I => \N__13234\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__13270\,
            I => \N__13229\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__13265\,
            I => \N__13229\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13226\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__13261\,
            I => \N__13223\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13218\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N__13218\
        );

    \I__2901\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13215\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__13247\,
            I => \bZ0Z_3\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__13244\,
            I => \bZ0Z_3\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__13239\,
            I => \bZ0Z_3\
        );

    \I__2897\ : Odrv12
    port map (
            O => \N__13234\,
            I => \bZ0Z_3\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__13229\,
            I => \bZ0Z_3\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__13226\,
            I => \bZ0Z_3\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__13223\,
            I => \bZ0Z_3\
        );

    \I__2893\ : Odrv12
    port map (
            O => \N__13218\,
            I => \bZ0Z_3\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__13215\,
            I => \bZ0Z_3\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__13196\,
            I => \N__13193\
        );

    \I__2890\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__2888\ : Odrv12
    port map (
            O => \N__13187\,
            I => \ALU.addsub_axb_3_l_ofxZ0\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__13184\,
            I => \N__13179\
        );

    \I__2886\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13175\
        );

    \I__2885\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13172\
        );

    \I__2884\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13168\
        );

    \I__2883\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13165\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13160\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__13172\,
            I => \N__13160\
        );

    \I__2880\ : InMux
    port map (
            O => \N__13171\,
            I => \N__13157\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__13168\,
            I => \N__13145\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13142\
        );

    \I__2877\ : Span4Mux_v
    port map (
            O => \N__13160\,
            I => \N__13137\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__13157\,
            I => \N__13137\
        );

    \I__2875\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13132\
        );

    \I__2874\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13132\
        );

    \I__2873\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13129\
        );

    \I__2872\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13126\
        );

    \I__2871\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13115\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13115\
        );

    \I__2869\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13115\
        );

    \I__2868\ : InMux
    port map (
            O => \N__13149\,
            I => \N__13115\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13115\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__13145\,
            I => \N__13108\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__13142\,
            I => \N__13108\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__13137\,
            I => \N__13108\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__13132\,
            I => \bZ0Z_8\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__13129\,
            I => \bZ0Z_8\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__13126\,
            I => \bZ0Z_8\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__13115\,
            I => \bZ0Z_8\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__13108\,
            I => \bZ0Z_8\
        );

    \I__2858\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__13094\,
            I => \ALU.regsA_result_cry_9_ma_2\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__13091\,
            I => \N__13086\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__13090\,
            I => \N__13082\
        );

    \I__2854\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13076\
        );

    \I__2853\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13073\
        );

    \I__2852\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13070\
        );

    \I__2851\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13064\
        );

    \I__2850\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13061\
        );

    \I__2849\ : InMux
    port map (
            O => \N__13080\,
            I => \N__13056\
        );

    \I__2848\ : InMux
    port map (
            O => \N__13079\,
            I => \N__13056\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__13076\,
            I => \N__13049\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13049\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__13070\,
            I => \N__13046\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__13069\,
            I => \N__13040\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__13068\,
            I => \N__13036\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__13067\,
            I => \N__13033\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__13064\,
            I => \N__13027\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__13061\,
            I => \N__13027\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__13024\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13019\
        );

    \I__2837\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13019\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__13049\,
            I => \N__13016\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__13046\,
            I => \N__13013\
        );

    \I__2834\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13010\
        );

    \I__2833\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13007\
        );

    \I__2832\ : InMux
    port map (
            O => \N__13043\,
            I => \N__12994\
        );

    \I__2831\ : InMux
    port map (
            O => \N__13040\,
            I => \N__12994\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13039\,
            I => \N__12994\
        );

    \I__2829\ : InMux
    port map (
            O => \N__13036\,
            I => \N__12994\
        );

    \I__2828\ : InMux
    port map (
            O => \N__13033\,
            I => \N__12994\
        );

    \I__2827\ : InMux
    port map (
            O => \N__13032\,
            I => \N__12994\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__13027\,
            I => \N__12989\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__13024\,
            I => \N__12989\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__13019\,
            I => \bZ0Z_6\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__13016\,
            I => \bZ0Z_6\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__13013\,
            I => \bZ0Z_6\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__13010\,
            I => \bZ0Z_6\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__13007\,
            I => \bZ0Z_6\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__12994\,
            I => \bZ0Z_6\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__12989\,
            I => \bZ0Z_6\
        );

    \I__2817\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12971\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__12971\,
            I => \ALU.regsA_result_cry_7_ma_3\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__12968\,
            I => \N__12963\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12958\
        );

    \I__2813\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12955\
        );

    \I__2812\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12952\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__12962\,
            I => \N__12942\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__12961\,
            I => \N__12935\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__12958\,
            I => \N__12931\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__12955\,
            I => \N__12921\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__12952\,
            I => \N__12921\
        );

    \I__2806\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12914\
        );

    \I__2805\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12914\
        );

    \I__2804\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12914\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12899\
        );

    \I__2802\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12899\
        );

    \I__2801\ : InMux
    port map (
            O => \N__12946\,
            I => \N__12899\
        );

    \I__2800\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12899\
        );

    \I__2799\ : InMux
    port map (
            O => \N__12942\,
            I => \N__12899\
        );

    \I__2798\ : InMux
    port map (
            O => \N__12941\,
            I => \N__12899\
        );

    \I__2797\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12899\
        );

    \I__2796\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12894\
        );

    \I__2795\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12894\
        );

    \I__2794\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12889\
        );

    \I__2793\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12889\
        );

    \I__2792\ : Span12Mux_v
    port map (
            O => \N__12931\,
            I => \N__12886\
        );

    \I__2791\ : InMux
    port map (
            O => \N__12930\,
            I => \N__12875\
        );

    \I__2790\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12875\
        );

    \I__2789\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12875\
        );

    \I__2788\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12875\
        );

    \I__2787\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12875\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__12921\,
            I => \N__12866\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__12914\,
            I => \N__12866\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__12899\,
            I => \N__12866\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__12894\,
            I => \N__12866\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__12889\,
            I => \aZ0Z_7\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__12886\,
            I => \aZ0Z_7\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__12875\,
            I => \aZ0Z_7\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__12866\,
            I => \aZ0Z_7\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__12857\,
            I => \N__12853\
        );

    \I__2777\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12846\
        );

    \I__2776\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12846\
        );

    \I__2775\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12839\
        );

    \I__2774\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12839\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__12846\,
            I => \N__12836\
        );

    \I__2772\ : InMux
    port map (
            O => \N__12845\,
            I => \N__12833\
        );

    \I__2771\ : InMux
    port map (
            O => \N__12844\,
            I => \N__12827\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__12839\,
            I => \N__12824\
        );

    \I__2769\ : Span4Mux_v
    port map (
            O => \N__12836\,
            I => \N__12821\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12818\
        );

    \I__2767\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12813\
        );

    \I__2766\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12813\
        );

    \I__2765\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12810\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__12827\,
            I => \N__12807\
        );

    \I__2763\ : Span4Mux_h
    port map (
            O => \N__12824\,
            I => \N__12798\
        );

    \I__2762\ : Span4Mux_v
    port map (
            O => \N__12821\,
            I => \N__12789\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__12818\,
            I => \N__12789\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12789\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__12810\,
            I => \N__12789\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__12807\,
            I => \N__12786\
        );

    \I__2757\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12781\
        );

    \I__2756\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12781\
        );

    \I__2755\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12772\
        );

    \I__2754\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12772\
        );

    \I__2753\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12772\
        );

    \I__2752\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12772\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__12798\,
            I => \bZ0Z_7\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__12789\,
            I => \bZ0Z_7\
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__12786\,
            I => \bZ0Z_7\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__12781\,
            I => \bZ0Z_7\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__12772\,
            I => \bZ0Z_7\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__2745\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__12755\,
            I => \ALU.regsA_result_cry_8_ma_2\
        );

    \I__2743\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__12746\,
            I => \N__12738\
        );

    \I__2740\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12733\
        );

    \I__2739\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12733\
        );

    \I__2738\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12728\
        );

    \I__2737\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12728\
        );

    \I__2736\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12725\
        );

    \I__2735\ : Span4Mux_h
    port map (
            O => \N__12738\,
            I => \N__12722\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__12733\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__12728\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__12725\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__12722\,
            I => \FTDI.baudAccZ0Z_2\
        );

    \I__2730\ : CEMux
    port map (
            O => \N__12713\,
            I => \N__12709\
        );

    \I__2729\ : CEMux
    port map (
            O => \N__12712\,
            I => \N__12706\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__12709\,
            I => \N__12703\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__12706\,
            I => \N__12700\
        );

    \I__2726\ : Span4Mux_v
    port map (
            O => \N__12703\,
            I => \N__12697\
        );

    \I__2725\ : Span4Mux_h
    port map (
            O => \N__12700\,
            I => \N__12694\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__12697\,
            I => \FTDI.un1_TXstate_0_sqmuxa_0_i\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__12694\,
            I => \FTDI.un1_TXstate_0_sqmuxa_0_i\
        );

    \I__2722\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12686\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__12683\,
            I => \N__12679\
        );

    \I__2719\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12676\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__12679\,
            I => \TXstartZ0\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__12676\,
            I => \TXstartZ0\
        );

    \I__2716\ : CEMux
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2714\ : Sp12to4
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__2713\ : Odrv12
    port map (
            O => \N__12662\,
            I => \un1_testState31_0_0\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__12656\,
            I => \ALU.regsA_result_cry_6_ma_3\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__12653\,
            I => \N__12645\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__12652\,
            I => \N__12642\
        );

    \I__2708\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12633\
        );

    \I__2707\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12633\
        );

    \I__2706\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12630\
        );

    \I__2705\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12627\
        );

    \I__2704\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12622\
        );

    \I__2703\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12619\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__12641\,
            I => \N__12616\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__12640\,
            I => \N__12612\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__12639\,
            I => \N__12609\
        );

    \I__2699\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12604\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12597\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12594\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__12627\,
            I => \N__12591\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__12626\,
            I => \N__12588\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__12625\,
            I => \N__12585\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__12622\,
            I => \N__12582\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__12619\,
            I => \N__12579\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12568\
        );

    \I__2690\ : InMux
    port map (
            O => \N__12615\,
            I => \N__12568\
        );

    \I__2689\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12568\
        );

    \I__2688\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12568\
        );

    \I__2687\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12568\
        );

    \I__2686\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12565\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__12604\,
            I => \N__12562\
        );

    \I__2684\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12559\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12602\,
            I => \N__12552\
        );

    \I__2682\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12552\
        );

    \I__2681\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12552\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__12597\,
            I => \N__12547\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__12594\,
            I => \N__12547\
        );

    \I__2678\ : Span4Mux_h
    port map (
            O => \N__12591\,
            I => \N__12544\
        );

    \I__2677\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12539\
        );

    \I__2676\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12539\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__12582\,
            I => \N__12530\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__12579\,
            I => \N__12530\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12530\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__12565\,
            I => \N__12530\
        );

    \I__2671\ : Odrv12
    port map (
            O => \N__12562\,
            I => \aZ0Z_1\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__12559\,
            I => \aZ0Z_1\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__12552\,
            I => \aZ0Z_1\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__12547\,
            I => \aZ0Z_1\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__12544\,
            I => \aZ0Z_1\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__12539\,
            I => \aZ0Z_1\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__12530\,
            I => \aZ0Z_1\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__2663\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12509\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__12506\,
            I => \ALU.regsA_result_axb_8_l_ofx\
        );

    \I__2660\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__12500\,
            I => \N__12497\
        );

    \I__2658\ : Span4Mux_h
    port map (
            O => \N__12497\,
            I => \N__12494\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__12494\,
            I => \ALU.regsA_result_cry_7_ma\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__2655\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__12485\,
            I => \N__12482\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__12479\,
            I => \ALU.regsA_result_axb_8_l_ofx_1\
        );

    \I__2651\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__12470\,
            I => \N__12467\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__12467\,
            I => \ALU.regsA_result_cry_9_ma_1\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__2646\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__12458\,
            I => \N__12450\
        );

    \I__2644\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12445\
        );

    \I__2643\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12445\
        );

    \I__2642\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12437\
        );

    \I__2641\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12437\
        );

    \I__2640\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12434\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__12450\,
            I => \N__12429\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__12445\,
            I => \N__12429\
        );

    \I__2637\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12424\
        );

    \I__2636\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12424\
        );

    \I__2635\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12421\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__12437\,
            I => \N__12418\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__12434\,
            I => \N__12413\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__12429\,
            I => \N__12413\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__12424\,
            I => \aZ0Z_2\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__12421\,
            I => \aZ0Z_2\
        );

    \I__2629\ : Odrv12
    port map (
            O => \N__12418\,
            I => \aZ0Z_2\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__12413\,
            I => \aZ0Z_2\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__2626\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12398\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__12398\,
            I => \N__12395\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__12392\,
            I => \ALU.regsA_result_axb_9_l_ofx_1\
        );

    \I__2622\ : InMux
    port map (
            O => \N__12389\,
            I => \N__12386\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__12386\,
            I => \ALU.regsA_result_axb_8_l_ofx_2\
        );

    \I__2620\ : InMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__12380\,
            I => \N__12375\
        );

    \I__2618\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12372\
        );

    \I__2617\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12365\
        );

    \I__2616\ : Span4Mux_v
    port map (
            O => \N__12375\,
            I => \N__12362\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__12372\,
            I => \N__12359\
        );

    \I__2614\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12356\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12348\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12343\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12343\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__12365\,
            I => \N__12340\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__12362\,
            I => \N__12337\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__12359\,
            I => \N__12332\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__12356\,
            I => \N__12332\
        );

    \I__2606\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12327\
        );

    \I__2605\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12327\
        );

    \I__2604\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12324\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12319\
        );

    \I__2602\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12319\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__12348\,
            I => \N__12314\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__12343\,
            I => \N__12314\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__12340\,
            I => \N__12311\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__12337\,
            I => \bZ0Z_9\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__12332\,
            I => \bZ0Z_9\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__12327\,
            I => \bZ0Z_9\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__12324\,
            I => \bZ0Z_9\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__12319\,
            I => \bZ0Z_9\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__12314\,
            I => \bZ0Z_9\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__12311\,
            I => \bZ0Z_9\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__12296\,
            I => \N__12293\
        );

    \I__2590\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12290\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__12290\,
            I => \ALU.regsA_result_axb_9_l_ofx_2\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12283\
        );

    \I__2587\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12278\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__12283\,
            I => \N__12275\
        );

    \I__2585\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12272\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12268\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12261\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__12275\,
            I => \N__12261\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12261\
        );

    \I__2580\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12258\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__12268\,
            I => \N__12255\
        );

    \I__2578\ : Span4Mux_v
    port map (
            O => \N__12261\,
            I => \N__12252\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12258\,
            I => \RXbuffer_5\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__12255\,
            I => \RXbuffer_5\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__12252\,
            I => \RXbuffer_5\
        );

    \I__2574\ : CEMux
    port map (
            O => \N__12245\,
            I => \N__12238\
        );

    \I__2573\ : CEMux
    port map (
            O => \N__12244\,
            I => \N__12235\
        );

    \I__2572\ : CEMux
    port map (
            O => \N__12243\,
            I => \N__12232\
        );

    \I__2571\ : CEMux
    port map (
            O => \N__12242\,
            I => \N__12228\
        );

    \I__2570\ : CEMux
    port map (
            O => \N__12241\,
            I => \N__12225\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__12238\,
            I => \N__12222\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__12235\,
            I => \N__12217\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__12232\,
            I => \N__12217\
        );

    \I__2566\ : CEMux
    port map (
            O => \N__12231\,
            I => \N__12214\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__12228\,
            I => \N__12210\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__12225\,
            I => \N__12207\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__12222\,
            I => \N__12200\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__12217\,
            I => \N__12200\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__12214\,
            I => \N__12200\
        );

    \I__2560\ : CEMux
    port map (
            O => \N__12213\,
            I => \N__12196\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__12210\,
            I => \N__12193\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__12207\,
            I => \N__12190\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__12200\,
            I => \N__12187\
        );

    \I__2556\ : CEMux
    port map (
            O => \N__12199\,
            I => \N__12184\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__12196\,
            I => \N__12181\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__12193\,
            I => \N__12176\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__12190\,
            I => \N__12176\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__12187\,
            I => \N__12173\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__12184\,
            I => \N__12170\
        );

    \I__2550\ : Span4Mux_h
    port map (
            O => \N__12181\,
            I => \N__12167\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__12176\,
            I => \RXready_RNIICV7_1\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__12173\,
            I => \RXready_RNIICV7_1\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__12170\,
            I => \RXready_RNIICV7_1\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__12167\,
            I => \RXready_RNIICV7_1\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__2544\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12152\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__12152\,
            I => \N__12149\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__12149\,
            I => \N__12146\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__12146\,
            I => \ALU.regsA_result_cry_1_ma\
        );

    \I__2540\ : InMux
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__2538\ : Span4Mux_v
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__12134\,
            I => \ALU.regsA_result_cry_3_ma_3\
        );

    \I__2536\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__12125\,
            I => \N__12122\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__12122\,
            I => \ALU.regsA_result_cry_2_ma\
        );

    \I__2532\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__12116\,
            I => \N__12111\
        );

    \I__2530\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12108\
        );

    \I__2529\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12105\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__12111\,
            I => \N__12100\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__12108\,
            I => \N__12097\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__12105\,
            I => \N__12094\
        );

    \I__2525\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12091\
        );

    \I__2524\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12088\
        );

    \I__2523\ : Span4Mux_h
    port map (
            O => \N__12100\,
            I => \N__12085\
        );

    \I__2522\ : Sp12to4
    port map (
            O => \N__12097\,
            I => \N__12082\
        );

    \I__2521\ : Span4Mux_v
    port map (
            O => \N__12094\,
            I => \N__12077\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__12091\,
            I => \N__12077\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__12088\,
            I => \RXbuffer_7\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__12085\,
            I => \RXbuffer_7\
        );

    \I__2517\ : Odrv12
    port map (
            O => \N__12082\,
            I => \RXbuffer_7\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__12077\,
            I => \RXbuffer_7\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__12068\,
            I => \N__12058\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__12067\,
            I => \N__12054\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__12066\,
            I => \N__12050\
        );

    \I__2512\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12045\
        );

    \I__2511\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12040\
        );

    \I__2510\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12040\
        );

    \I__2509\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12037\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__12061\,
            I => \N__12030\
        );

    \I__2507\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12027\
        );

    \I__2506\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12022\
        );

    \I__2505\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12019\
        );

    \I__2504\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12014\
        );

    \I__2503\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12014\
        );

    \I__2502\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12010\
        );

    \I__2501\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12007\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__12045\,
            I => \N__12000\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__12040\,
            I => \N__12000\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__12037\,
            I => \N__12000\
        );

    \I__2497\ : InMux
    port map (
            O => \N__12036\,
            I => \N__11995\
        );

    \I__2496\ : InMux
    port map (
            O => \N__12035\,
            I => \N__11995\
        );

    \I__2495\ : InMux
    port map (
            O => \N__12034\,
            I => \N__11990\
        );

    \I__2494\ : InMux
    port map (
            O => \N__12033\,
            I => \N__11987\
        );

    \I__2493\ : InMux
    port map (
            O => \N__12030\,
            I => \N__11984\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__12027\,
            I => \N__11981\
        );

    \I__2491\ : InMux
    port map (
            O => \N__12026\,
            I => \N__11976\
        );

    \I__2490\ : InMux
    port map (
            O => \N__12025\,
            I => \N__11976\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__11971\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__12019\,
            I => \N__11971\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__12014\,
            I => \N__11964\
        );

    \I__2486\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11961\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__11952\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__12007\,
            I => \N__11952\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__12000\,
            I => \N__11952\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11995\,
            I => \N__11952\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__11994\,
            I => \N__11949\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__11993\,
            I => \N__11941\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__11990\,
            I => \N__11933\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11933\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__11984\,
            I => \N__11933\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__11981\,
            I => \N__11926\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__11976\,
            I => \N__11926\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__11971\,
            I => \N__11926\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11970\,
            I => \N__11923\
        );

    \I__2472\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11920\
        );

    \I__2471\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11915\
        );

    \I__2470\ : InMux
    port map (
            O => \N__11967\,
            I => \N__11915\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__11964\,
            I => \N__11908\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__11961\,
            I => \N__11908\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__11952\,
            I => \N__11908\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11949\,
            I => \N__11905\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__11948\,
            I => \N__11901\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__11947\,
            I => \N__11898\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11946\,
            I => \N__11895\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11892\
        );

    \I__2461\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11887\
        );

    \I__2460\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11887\
        );

    \I__2459\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11884\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__11933\,
            I => \N__11879\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__11926\,
            I => \N__11879\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__11923\,
            I => \N__11876\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__11920\,
            I => \N__11873\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__11915\,
            I => \N__11866\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__11908\,
            I => \N__11866\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11866\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11859\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11859\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11859\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__11895\,
            I => \bZ0Z_1\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__11892\,
            I => \bZ0Z_1\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__11887\,
            I => \bZ0Z_1\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__11884\,
            I => \bZ0Z_1\
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__11879\,
            I => \bZ0Z_1\
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__11876\,
            I => \bZ0Z_1\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__11873\,
            I => \bZ0Z_1\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__11866\,
            I => \bZ0Z_1\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__11859\,
            I => \bZ0Z_1\
        );

    \I__2439\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11837\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__11837\,
            I => \ALU.regsA_result_cry_2_ma_5\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__11834\,
            I => \N__11828\
        );

    \I__2436\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11821\
        );

    \I__2435\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11818\
        );

    \I__2434\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11815\
        );

    \I__2433\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11811\
        );

    \I__2432\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11808\
        );

    \I__2431\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11803\
        );

    \I__2430\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11803\
        );

    \I__2429\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11800\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11794\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__11818\,
            I => \N__11789\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__11815\,
            I => \N__11789\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__11814\,
            I => \N__11786\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__11811\,
            I => \N__11776\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__11808\,
            I => \N__11776\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__11803\,
            I => \N__11771\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__11800\,
            I => \N__11771\
        );

    \I__2420\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11766\
        );

    \I__2419\ : InMux
    port map (
            O => \N__11798\,
            I => \N__11766\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11797\,
            I => \N__11763\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__11794\,
            I => \N__11758\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__11789\,
            I => \N__11758\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11753\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11753\
        );

    \I__2413\ : InMux
    port map (
            O => \N__11784\,
            I => \N__11750\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11783\,
            I => \N__11743\
        );

    \I__2411\ : InMux
    port map (
            O => \N__11782\,
            I => \N__11738\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11738\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__11776\,
            I => \N__11731\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__11771\,
            I => \N__11731\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__11766\,
            I => \N__11731\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__11763\,
            I => \N__11724\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__11758\,
            I => \N__11724\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__11753\,
            I => \N__11719\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__11750\,
            I => \N__11719\
        );

    \I__2402\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11716\
        );

    \I__2401\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11711\
        );

    \I__2400\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11711\
        );

    \I__2399\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11708\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N__11705\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11700\
        );

    \I__2396\ : Span4Mux_h
    port map (
            O => \N__11731\,
            I => \N__11700\
        );

    \I__2395\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11695\
        );

    \I__2394\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11695\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__11724\,
            I => \bZ0Z_2\
        );

    \I__2392\ : Odrv12
    port map (
            O => \N__11719\,
            I => \bZ0Z_2\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__11716\,
            I => \bZ0Z_2\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__11711\,
            I => \bZ0Z_2\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__11708\,
            I => \bZ0Z_2\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__11705\,
            I => \bZ0Z_2\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__11700\,
            I => \bZ0Z_2\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__11695\,
            I => \bZ0Z_2\
        );

    \I__2385\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__11675\,
            I => \ALU.regsA_result_cry_3_ma_5\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__11672\,
            I => \N__11669\
        );

    \I__2382\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__11666\,
            I => \ALU.regsA_result_cry_4_ma_4\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__11663\,
            I => \N__11654\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__11662\,
            I => \N__11647\
        );

    \I__2378\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11641\
        );

    \I__2377\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11638\
        );

    \I__2376\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11635\
        );

    \I__2375\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11630\
        );

    \I__2374\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11630\
        );

    \I__2373\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11627\
        );

    \I__2372\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11620\
        );

    \I__2371\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11620\
        );

    \I__2370\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11620\
        );

    \I__2369\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11617\
        );

    \I__2368\ : InMux
    port map (
            O => \N__11647\,
            I => \N__11612\
        );

    \I__2367\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11612\
        );

    \I__2366\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11607\
        );

    \I__2365\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11603\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__11641\,
            I => \N__11595\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__11638\,
            I => \N__11595\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__11635\,
            I => \N__11595\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__11630\,
            I => \N__11592\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__11627\,
            I => \N__11587\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__11620\,
            I => \N__11587\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__11617\,
            I => \N__11580\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__11612\,
            I => \N__11580\
        );

    \I__2356\ : InMux
    port map (
            O => \N__11611\,
            I => \N__11577\
        );

    \I__2355\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11574\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11571\
        );

    \I__2353\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11568\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__11603\,
            I => \N__11565\
        );

    \I__2351\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11562\
        );

    \I__2350\ : Span4Mux_v
    port map (
            O => \N__11595\,
            I => \N__11555\
        );

    \I__2349\ : Span4Mux_v
    port map (
            O => \N__11592\,
            I => \N__11555\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__11587\,
            I => \N__11555\
        );

    \I__2347\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11550\
        );

    \I__2346\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11550\
        );

    \I__2345\ : Span4Mux_h
    port map (
            O => \N__11580\,
            I => \N__11547\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11542\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11542\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__11571\,
            I => \N__11535\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__11568\,
            I => \N__11535\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__11565\,
            I => \N__11535\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__11562\,
            I => \bZ0Z_4\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__11555\,
            I => \bZ0Z_4\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__11550\,
            I => \bZ0Z_4\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__11547\,
            I => \bZ0Z_4\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__11542\,
            I => \bZ0Z_4\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__11535\,
            I => \bZ0Z_4\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__11519\,
            I => \ALU.regsA_result_cry_5_ma_4\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__11516\,
            I => \FTDI.N_23_cascade_\
        );

    \I__2330\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11498\
        );

    \I__2329\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11498\
        );

    \I__2328\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11498\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11510\,
            I => \N__11498\
        );

    \I__2326\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11498\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__11498\,
            I => \FTDI.RXstateZ0Z_0\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__11495\,
            I => \N__11485\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__11494\,
            I => \N__11481\
        );

    \I__2322\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11476\
        );

    \I__2321\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11476\
        );

    \I__2320\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11461\
        );

    \I__2319\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11461\
        );

    \I__2318\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11461\
        );

    \I__2317\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11461\
        );

    \I__2316\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11461\
        );

    \I__2315\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11461\
        );

    \I__2314\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11461\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__11476\,
            I => \FTDI.RXstateZ0Z_3\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__11461\,
            I => \FTDI.RXstateZ0Z_3\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__11456\,
            I => \N__11453\
        );

    \I__2310\ : InMux
    port map (
            O => \N__11453\,
            I => \N__11444\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11444\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11437\
        );

    \I__2307\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11437\
        );

    \I__2306\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11437\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__11444\,
            I => \FTDI.RXstateZ0Z_2\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__11437\,
            I => \FTDI.RXstateZ0Z_2\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__11432\,
            I => \N__11428\
        );

    \I__2302\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11423\
        );

    \I__2301\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11423\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__11423\,
            I => \FTDI.N_28\
        );

    \I__2299\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11410\
        );

    \I__2298\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11410\
        );

    \I__2297\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11401\
        );

    \I__2296\ : InMux
    port map (
            O => \N__11417\,
            I => \N__11401\
        );

    \I__2295\ : InMux
    port map (
            O => \N__11416\,
            I => \N__11401\
        );

    \I__2294\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11401\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__11410\,
            I => \FTDI.RXstateZ0Z_1\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__11401\,
            I => \FTDI.RXstateZ0Z_1\
        );

    \I__2291\ : CEMux
    port map (
            O => \N__11396\,
            I => \N__11391\
        );

    \I__2290\ : CEMux
    port map (
            O => \N__11395\,
            I => \N__11388\
        );

    \I__2289\ : CEMux
    port map (
            O => \N__11394\,
            I => \N__11384\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__11391\,
            I => \N__11381\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__11388\,
            I => \N__11378\
        );

    \I__2286\ : CEMux
    port map (
            O => \N__11387\,
            I => \N__11375\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__11384\,
            I => \N__11371\
        );

    \I__2284\ : Span4Mux_v
    port map (
            O => \N__11381\,
            I => \N__11368\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__11378\,
            I => \N__11363\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__11375\,
            I => \N__11363\
        );

    \I__2281\ : CEMux
    port map (
            O => \N__11374\,
            I => \N__11360\
        );

    \I__2280\ : Span4Mux_h
    port map (
            O => \N__11371\,
            I => \N__11357\
        );

    \I__2279\ : Span4Mux_h
    port map (
            O => \N__11368\,
            I => \N__11354\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__11363\,
            I => \N__11349\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11349\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__11357\,
            I => \N__11346\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__11354\,
            I => \N__11341\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__11349\,
            I => \N__11341\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__11346\,
            I => \RXready_RNIICV7_0\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__11341\,
            I => \RXready_RNIICV7_0\
        );

    \I__2271\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__11333\,
            I => \N__11328\
        );

    \I__2269\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11325\
        );

    \I__2268\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11322\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__11328\,
            I => \N__11315\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__11325\,
            I => \N__11315\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__11322\,
            I => \N__11311\
        );

    \I__2264\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11308\
        );

    \I__2263\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11305\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__11315\,
            I => \N__11302\
        );

    \I__2261\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11299\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__11311\,
            I => \N__11294\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__11308\,
            I => \N__11294\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__11305\,
            I => \RXbuffer_1\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__11302\,
            I => \RXbuffer_1\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__11299\,
            I => \RXbuffer_1\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__11294\,
            I => \RXbuffer_1\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__11285\,
            I => \N__11273\
        );

    \I__2253\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11266\
        );

    \I__2252\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11266\
        );

    \I__2251\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11257\
        );

    \I__2250\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11257\
        );

    \I__2249\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11257\
        );

    \I__2248\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11254\
        );

    \I__2247\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11241\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11241\
        );

    \I__2245\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11241\
        );

    \I__2244\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11241\
        );

    \I__2243\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11241\
        );

    \I__2242\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11241\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__11266\,
            I => \N__11238\
        );

    \I__2240\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11235\
        );

    \I__2239\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11232\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11223\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__11254\,
            I => \N__11223\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__11241\,
            I => \N__11223\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__11238\,
            I => \N__11216\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__11235\,
            I => \N__11216\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__11232\,
            I => \N__11216\
        );

    \I__2232\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11213\
        );

    \I__2231\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11210\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__11223\,
            I => \N__11207\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__11216\,
            I => \N__11204\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__11213\,
            I => \N__11197\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__11210\,
            I => \N__11197\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__11207\,
            I => \N__11194\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__11204\,
            I => \N__11191\
        );

    \I__2224\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11186\
        );

    \I__2223\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11186\
        );

    \I__2222\ : Span4Mux_h
    port map (
            O => \N__11197\,
            I => \N__11181\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__11194\,
            I => \N__11181\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__11191\,
            I => \opZ0Z_1\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__11186\,
            I => \opZ0Z_1\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__11181\,
            I => \opZ0Z_1\
        );

    \I__2217\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11171\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__2214\ : Span4Mux_h
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__11162\,
            I => \ALU.addsub_4\
        );

    \I__2212\ : InMux
    port map (
            O => \N__11159\,
            I => \N__11156\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__11156\,
            I => \ALU.mult_4\
        );

    \I__2210\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__2208\ : Sp12to4
    port map (
            O => \N__11147\,
            I => \N__11144\
        );

    \I__2207\ : Span12Mux_v
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__2206\ : Odrv12
    port map (
            O => \N__11141\,
            I => res_4
        );

    \I__2205\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__2203\ : Span12Mux_v
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__2202\ : Odrv12
    port map (
            O => \N__11129\,
            I => \ALU.regsA_result_cry_2_ma_0\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__2200\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__11117\,
            I => \N__11114\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__11114\,
            I => \N__11111\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__11111\,
            I => \ALU.regsA_result_cry_10_ma_1\
        );

    \I__2195\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11100\
        );

    \I__2194\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11100\
        );

    \I__2193\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11096\
        );

    \I__2192\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11091\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11088\
        );

    \I__2190\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11085\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__11096\,
            I => \N__11081\
        );

    \I__2188\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11078\
        );

    \I__2187\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11075\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__11091\,
            I => \N__11072\
        );

    \I__2185\ : Span12Mux_h
    port map (
            O => \N__11088\,
            I => \N__11067\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__11085\,
            I => \N__11067\
        );

    \I__2183\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11064\
        );

    \I__2182\ : Span4Mux_h
    port map (
            O => \N__11081\,
            I => \N__11061\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__11078\,
            I => \N__11058\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__11075\,
            I => \N__11053\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__11072\,
            I => \N__11053\
        );

    \I__2178\ : Span12Mux_v
    port map (
            O => \N__11067\,
            I => \N__11050\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__11064\,
            I => \RXbuffer_2\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__11061\,
            I => \RXbuffer_2\
        );

    \I__2175\ : Odrv12
    port map (
            O => \N__11058\,
            I => \RXbuffer_2\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__11053\,
            I => \RXbuffer_2\
        );

    \I__2173\ : Odrv12
    port map (
            O => \N__11050\,
            I => \RXbuffer_2\
        );

    \I__2172\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__2170\ : Odrv12
    port map (
            O => \N__11033\,
            I => \TXbufferZ0Z_7\
        );

    \I__2169\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__11027\,
            I => \FTDI.TXshiftZ0Z_7\
        );

    \I__2167\ : InMux
    port map (
            O => \N__11024\,
            I => \N__11020\
        );

    \I__2166\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11017\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__11020\,
            I => \N__11012\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__11012\
        );

    \I__2163\ : Span4Mux_h
    port map (
            O => \N__11012\,
            I => \N__11009\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__11006\,
            I => \N__11003\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__11003\,
            I => \RX_c\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__11000\,
            I => \FTDI.m13_ns_1_cascade_\
        );

    \I__2158\ : CEMux
    port map (
            O => \N__10997\,
            I => \N__10994\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__10994\,
            I => \N__10990\
        );

    \I__2156\ : CEMux
    port map (
            O => \N__10993\,
            I => \N__10987\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__10990\,
            I => \N__10984\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10981\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__10984\,
            I => \N__10978\
        );

    \I__2152\ : Span4Mux_h
    port map (
            O => \N__10981\,
            I => \N__10975\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__10978\,
            I => \FTDI.N_201_2\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__10975\,
            I => \FTDI.N_201_2\
        );

    \I__2149\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__10964\,
            I => \N__10960\
        );

    \I__2146\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__2145\ : Span4Mux_h
    port map (
            O => \N__10960\,
            I => \N__10950\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10957\,
            I => \N__10950\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10947\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10944\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__10950\,
            I => \N__10939\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10936\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__10944\,
            I => \N__10933\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10930\
        );

    \I__2137\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10927\
        );

    \I__2136\ : Span4Mux_h
    port map (
            O => \N__10939\,
            I => \N__10924\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__10936\,
            I => \N__10917\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__10933\,
            I => \N__10917\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__10930\,
            I => \N__10917\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__10927\,
            I => \RXbuffer_4\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__10924\,
            I => \RXbuffer_4\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__10917\,
            I => \RXbuffer_4\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__10910\,
            I => \N__10907\
        );

    \I__2128\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10904\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__10904\,
            I => \ALU.regsA_result_axb_5_l_ofx_2\
        );

    \I__2126\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__10892\,
            I => \ALU.addsub_axb_4_l_ofxZ0\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10886\,
            I => \ALU.regsA_result_cry_4_ma_2\
        );

    \I__2120\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10880\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__10880\,
            I => \ALU.regsA_result_cry_5_ma_2\
        );

    \I__2118\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__10874\,
            I => \ALU.regsA_result_cry_6_ma_1\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__2115\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__10859\,
            I => \ALU.regsA_result_axb_9_l_ofx\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__2110\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10849\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10844\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__10849\,
            I => \N__10840\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__10848\,
            I => \N__10837\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__10847\,
            I => \N__10834\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10830\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__10843\,
            I => \N__10824\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__10840\,
            I => \N__10819\
        );

    \I__2102\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10814\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10814\
        );

    \I__2100\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10811\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__10830\,
            I => \N__10808\
        );

    \I__2098\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10803\
        );

    \I__2097\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10803\
        );

    \I__2096\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10800\
        );

    \I__2095\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10793\
        );

    \I__2094\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10793\
        );

    \I__2093\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10793\
        );

    \I__2092\ : Span4Mux_h
    port map (
            O => \N__10819\,
            I => \N__10786\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__10814\,
            I => \N__10786\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__10811\,
            I => \N__10786\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__10808\,
            I => \aZ0Z_4\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__10803\,
            I => \aZ0Z_4\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__10800\,
            I => \aZ0Z_4\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__10793\,
            I => \aZ0Z_4\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__10786\,
            I => \aZ0Z_4\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__2083\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__10769\,
            I => \ALU.regsA_result_axb_9_l_ofx_0\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__10754\,
            I => \ALU.mult_AdderTree2_bigtree_642\
        );

    \I__2076\ : InMux
    port map (
            O => \N__10751\,
            I => \bfn_15_14_0_\
        );

    \I__2075\ : InMux
    port map (
            O => \N__10748\,
            I => \ALU.regsA_result_cry_9\
        );

    \I__2074\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__10739\,
            I => \ALU.regsA_result_cry_9_THRU_CO\
        );

    \I__2071\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__10727\,
            I => \ALU.regsA_result_cry_9_ma_0\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__2066\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__10718\,
            I => \ALU.regsA_result_cry_2_ma_3\
        );

    \I__2064\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__10712\,
            I => \ALU.regsA_result_cry_7_ma_1\
        );

    \I__2062\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__10703\,
            I => \ALU.regsA_result_axb_10\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__2058\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__10694\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_4\
        );

    \I__2056\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__10688\,
            I => \N__10685\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__10685\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_6\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__2052\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__10676\,
            I => \ALU.regsA_result_axb_4_l_ofx_2\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__2049\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__10667\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_5\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__2046\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__10658\,
            I => \ALU.regsA_result_axb_2_l_ofx_5\
        );

    \I__2044\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__10646\,
            I => \ALU.mult_AdderTree2_bigtree_635\
        );

    \I__2040\ : InMux
    port map (
            O => \N__10643\,
            I => \ALU.regsA_result_cry_1_9\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__2038\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__10634\,
            I => \ALU.regsA_result_axb_3_l_ofx_5\
        );

    \I__2036\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__10622\,
            I => \ALU.mult_AdderTree2_bigtree_636\
        );

    \I__2032\ : InMux
    port map (
            O => \N__10619\,
            I => \ALU.regsA_result_cry_2_11\
        );

    \I__2031\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__10613\,
            I => \ALU.regsA_result_axb_4_l_ofx_4\
        );

    \I__2029\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__10601\,
            I => \ALU.mult_AdderTree2_bigtree_637\
        );

    \I__2025\ : InMux
    port map (
            O => \N__10598\,
            I => \ALU.regsA_result_cry_3_11\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2023\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10589\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__10589\,
            I => \ALU.regsA_result_axb_5_l_ofx_4\
        );

    \I__2021\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__10580\,
            I => \N__10577\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__10577\,
            I => \ALU.mult_AdderTree2_bigtree_638\
        );

    \I__2017\ : InMux
    port map (
            O => \N__10574\,
            I => \ALU.regsA_result_cry_4_10\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__10571\,
            I => \N__10568\
        );

    \I__2015\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10565\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__10565\,
            I => \ALU.regsA_result_axb_6_l_ofx_3\
        );

    \I__2013\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10559\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__10559\,
            I => \N__10556\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__10556\,
            I => \N__10553\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__10553\,
            I => \ALU.mult_AdderTree2_bigtree_639\
        );

    \I__2009\ : InMux
    port map (
            O => \N__10550\,
            I => \ALU.regsA_result_cry_5_10\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__10547\,
            I => \N__10544\
        );

    \I__2007\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__10541\,
            I => \ALU.regsA_result_axb_7_l_ofx_3\
        );

    \I__2005\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__10529\,
            I => \ALU.mult_AdderTree2_bigtree_640\
        );

    \I__2001\ : InMux
    port map (
            O => \N__10526\,
            I => \ALU.regsA_result_cry_6_9\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__1999\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10517\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__1997\ : Span4Mux_h
    port map (
            O => \N__10514\,
            I => \N__10511\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__10511\,
            I => \ALU.mult_AdderTree2_bigtree_641\
        );

    \I__1995\ : InMux
    port map (
            O => \N__10508\,
            I => \ALU.regsA_result_cry_7_8\
        );

    \I__1994\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10500\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__10504\,
            I => \N__10496\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__10503\,
            I => \N__10492\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__10500\,
            I => \N__10488\
        );

    \I__1990\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10477\
        );

    \I__1989\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10477\
        );

    \I__1988\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10477\
        );

    \I__1987\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10477\
        );

    \I__1986\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10477\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__10488\,
            I => \a_fastZ0Z_4\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__10477\,
            I => \a_fastZ0Z_4\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__10472\,
            I => \N__10467\
        );

    \I__1982\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10462\
        );

    \I__1981\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10462\
        );

    \I__1980\ : InMux
    port map (
            O => \N__10467\,
            I => \N__10459\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10456\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__10456\,
            I => \N__10448\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__10453\,
            I => \N__10448\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__10448\,
            I => \ALU.mult_AdderTree2_bigtree_796\
        );

    \I__1974\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__1971\ : Span4Mux_h
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__10430\,
            I => \ALU.mult_AdderTree2_bigtree_634\
        );

    \I__1968\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__10421\,
            I => \N__10414\
        );

    \I__1965\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10411\
        );

    \I__1964\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10408\
        );

    \I__1963\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10405\
        );

    \I__1962\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10402\
        );

    \I__1961\ : Span4Mux_h
    port map (
            O => \N__10414\,
            I => \N__10395\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__10411\,
            I => \N__10395\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10395\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__10405\,
            I => \RXbuffer_3\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__10402\,
            I => \RXbuffer_3\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__10395\,
            I => \RXbuffer_3\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__1954\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__10373\,
            I => \ALU.mult_AdderTree2_bigtree_599\
        );

    \I__1949\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1946\ : Odrv4
    port map (
            O => \N__10361\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_3\
        );

    \I__1945\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__10349\,
            I => \ALU.regsA_result_axb_2_l_ofx_3\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__1940\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__10334\,
            I => \ALU.regsA_result_axb_3_l_ofx_3\
        );

    \I__1936\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__10322\,
            I => \ALU.regsA_result_cry_0_c_RNO\
        );

    \I__1932\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__10316\,
            I => \FTDI.TXshiftZ0Z_6\
        );

    \I__1930\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__10307\,
            I => \TXbufferZ0Z_5\
        );

    \I__1927\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__10301\,
            I => \FTDI.TXshiftZ0Z_5\
        );

    \I__1925\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10295\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__10295\,
            I => \ALU.regsA_result_cry_11_ma_0\
        );

    \I__1923\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10288\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__10291\,
            I => \N__10283\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__10288\,
            I => \N__10280\
        );

    \I__1920\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10277\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10272\
        );

    \I__1918\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10268\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__10280\,
            I => \N__10263\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10263\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__10276\,
            I => \N__10259\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10255\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10250\
        );

    \I__1912\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10250\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__10268\,
            I => \N__10247\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__10263\,
            I => \N__10244\
        );

    \I__1909\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10237\
        );

    \I__1908\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10237\
        );

    \I__1907\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10237\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__10255\,
            I => \bZ0Z_11\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__10250\,
            I => \bZ0Z_11\
        );

    \I__1904\ : Odrv12
    port map (
            O => \N__10247\,
            I => \bZ0Z_11\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__10244\,
            I => \bZ0Z_11\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__10237\,
            I => \bZ0Z_11\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__10226\,
            I => \N__10223\
        );

    \I__1900\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10220\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__10220\,
            I => \ALU.regsA_result_axb_11_l_ofx_0\
        );

    \I__1898\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__10214\,
            I => \ALU.regsA_result_cry_10_ma_0\
        );

    \I__1896\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__10208\,
            I => \TXbufferZ0Z_1\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__10199\,
            I => \TXbufferZ0Z_2\
        );

    \I__1891\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__10193\,
            I => \FTDI.TXshiftZ0Z_2\
        );

    \I__1889\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__10184\,
            I => \TXbufferZ0Z_6\
        );

    \I__1886\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__10178\,
            I => \TXbufferZ0Z_4\
        );

    \I__1884\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__10172\,
            I => \FTDI.TXshiftZ0Z_1\
        );

    \I__1882\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__10163\,
            I => \TXbufferZ0Z_0\
        );

    \I__1879\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__10157\,
            I => \FTDI.TXshiftZ0Z_4\
        );

    \I__1877\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10151\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__10151\,
            I => \TXbufferZ0Z_3\
        );

    \I__1875\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__10145\,
            I => \FTDI.TXshiftZ0Z_3\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1872\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10136\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__10133\,
            I => \ALU.regsA_result_axb_6_l_ofx_1\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1868\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__10124\,
            I => \ALU.mult_AdderTree2_bigtree_604\
        );

    \I__1866\ : InMux
    port map (
            O => \N__10121\,
            I => \ALU.regsA_result_cry_5_8\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__1864\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__10112\,
            I => \ALU.regsA_result_axb_7_l_ofx_1\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__1861\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__10103\,
            I => \ALU.mult_AdderTree2_bigtree_605\
        );

    \I__1859\ : InMux
    port map (
            O => \N__10100\,
            I => \ALU.regsA_result_cry_6_7\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__10091\,
            I => \ALU.regsA_result_axb_8_l_ofx_0\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__1854\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__10079\,
            I => \ALU.regsA_result_cry_8_ma_0\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1850\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__10070\,
            I => \ALU.mult_AdderTree2_bigtree_606\
        );

    \I__1848\ : InMux
    port map (
            O => \N__10067\,
            I => \ALU.regsA_result_cry_7_6\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__1846\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__10058\,
            I => \ALU.mult_AdderTree2_bigtree_607\
        );

    \I__1844\ : InMux
    port map (
            O => \N__10055\,
            I => \bfn_14_16_0_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__10049\,
            I => \ALU.mult_AdderTree2_bigtree_608\
        );

    \I__1841\ : InMux
    port map (
            O => \N__10046\,
            I => \ALU.regsA_result_cry_9_4\
        );

    \I__1840\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10040\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__10040\,
            I => \ALU.mult_AdderTree2_bigtree_609\
        );

    \I__1838\ : InMux
    port map (
            O => \N__10037\,
            I => \ALU.regsA_result_cry_10_3\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__1836\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10028\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__10022\,
            I => \ALU.regsA_result_axb_12_1\
        );

    \I__1832\ : InMux
    port map (
            O => \N__10019\,
            I => \ALU.regsA_result_cry_11_1\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__10016\,
            I => \N__10013\
        );

    \I__1830\ : InMux
    port map (
            O => \N__10013\,
            I => \N__10010\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__10010\,
            I => \N__10007\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__10007\,
            I => \N__10004\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__10004\,
            I => \ALU.regsA_result_axb_12\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__1825\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__9995\,
            I => \ALU.regsA_result_axb_10_l_ofx_0\
        );

    \I__1823\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__9986\,
            I => \ALU.regsA_result_cry_8_ma_1\
        );

    \I__1820\ : InMux
    port map (
            O => \N__9983\,
            I => \ALU.regsA_result_cry_1_7\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__1818\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__9974\,
            I => \ALU.mult_AdderTree2_bigtree_601\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9971\,
            I => \ALU.regsA_result_cry_2_9\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__9962\,
            I => \ALU.mult_AdderTree2_bigtree_602\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9959\,
            I => \ALU.regsA_result_cry_3_9\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1810\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9950\,
            I => \ALU.mult_AdderTree2_bigtree_603\
        );

    \I__1808\ : InMux
    port map (
            O => \N__9947\,
            I => \ALU.regsA_result_cry_4_8\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1806\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__9938\,
            I => \N__9935\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__9932\,
            I => \ALU.regsA_result_axb_6_l_ofx\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__1801\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__9917\,
            I => \ALU.regsA_result_cry_5_ma\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__9905\,
            I => \ALU.regsA_result_axb_6_l_ofx_2\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__9893\,
            I => \ALU.regsA_result_cry_7_ma_2\
        );

    \I__1789\ : InMux
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__1787\ : Span4Mux_h
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__9881\,
            I => \ALU.regsA_result_axb_7_l_ofx_2\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__9869\,
            I => \ALU.regsA_result_cry_6_ma\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9863\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__9863\,
            I => \ALU.regsA_result_cry_2_ma_4\
        );

    \I__1779\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__9857\,
            I => \ALU.regsA_result_cry_3_ma_4\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__9854\,
            I => \N__9851\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__9848\,
            I => \ALU.regsA_result_cry_4_ma_3\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__9845\,
            I => \N__9842\
        );

    \I__1773\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__9833\,
            I => \ALU.mult_AdderTree2_bigtree_831\
        );

    \I__1769\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9825\
        );

    \I__1768\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9822\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__9828\,
            I => \N__9819\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__9825\,
            I => \N__9816\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9822\,
            I => \N__9813\
        );

    \I__1764\ : InMux
    port map (
            O => \N__9819\,
            I => \N__9810\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__9816\,
            I => \ALU.mult_AdderTree2_bigtree_530\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__9813\,
            I => \ALU.mult_AdderTree2_bigtree_530\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__9810\,
            I => \ALU.mult_AdderTree2_bigtree_530\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9798\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9795\
        );

    \I__1758\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9792\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__9798\,
            I => \N__9786\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__9795\,
            I => \N__9783\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9780\
        );

    \I__1754\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9777\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__9790\,
            I => \N__9774\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__9789\,
            I => \N__9770\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__9786\,
            I => \N__9764\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__9783\,
            I => \N__9764\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__9780\,
            I => \N__9759\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__9777\,
            I => \N__9759\
        );

    \I__1747\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9750\
        );

    \I__1746\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9750\
        );

    \I__1745\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9750\
        );

    \I__1744\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9750\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__9764\,
            I => \a_2_repZ0Z1\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__9759\,
            I => \a_2_repZ0Z1\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__9750\,
            I => \a_2_repZ0Z1\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__9740\,
            I => \ALU.regsA_result_cry_0_c_RNO_0\
        );

    \I__1738\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9734\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__9734\,
            I => \N__9731\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__9731\,
            I => \ALU.regsA_result_cry_4_ma\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1734\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__1732\ : Span4Mux_h
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__9716\,
            I => \ALU.regsA_result_cry_6_ma_2\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__1729\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__9707\,
            I => \ALU.regsA_result_axb_2_l_ofx_4\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__1726\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__9698\,
            I => \ALU.regsA_result_axb_3_l_ofx_4\
        );

    \I__1724\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__9692\,
            I => \ALU.regsA_result_axb_4_l_ofx_3\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__1721\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__9683\,
            I => \ALU.regsA_result_axb_5_l_ofx_3\
        );

    \I__1719\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__9674\,
            I => \ALU.mult_AdderTree2_bigtree_564\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__1715\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9664\
        );

    \I__1714\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__9664\,
            I => \a_fastZ0Z_2\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__9661\,
            I => \a_fastZ0Z_2\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__1710\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__9650\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_4\
        );

    \I__1708\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9644\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__9644\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_5\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__9641\,
            I => \N__9638\
        );

    \I__1705\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__9635\,
            I => \N__9632\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__9629\,
            I => \ALU.regsA_result_axb_11_l_ofx\
        );

    \I__1701\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__9617\,
            I => \N__9614\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__9614\,
            I => \ALU.regsA_result_cry_10_ma\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__9611\,
            I => \N__9608\
        );

    \I__1695\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__9605\,
            I => \N__9602\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__9602\,
            I => \ALU.regsA_result_axb_11_l_ofx_1\
        );

    \I__1692\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__9596\,
            I => \N__9590\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__9595\,
            I => \N__9587\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__9594\,
            I => \N__9584\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__9593\,
            I => \N__9578\
        );

    \I__1687\ : Span4Mux_h
    port map (
            O => \N__9590\,
            I => \N__9574\
        );

    \I__1686\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9565\
        );

    \I__1685\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9565\
        );

    \I__1684\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9565\
        );

    \I__1683\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9565\
        );

    \I__1682\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9558\
        );

    \I__1681\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9558\
        );

    \I__1680\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9558\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__9574\,
            I => \bZ0Z_12\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__9565\,
            I => \bZ0Z_12\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__9558\,
            I => \bZ0Z_12\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__1675\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__9545\,
            I => \N__9542\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__9539\,
            I => \ALU.regsA_result_axb_12_l_ofx_0\
        );

    \I__1671\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9530\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__9530\,
            I => \ALU.regsA_result_axb_10_l_ofx_1\
        );

    \I__1668\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9524\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__1666\ : Span4Mux_v
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__9518\,
            I => \ALU.regsA_result_cry_11_ma_1\
        );

    \I__1664\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__9512\,
            I => \ALU.mult_AdderTree2_bigtree_840\
        );

    \I__1662\ : InMux
    port map (
            O => \N__9509\,
            I => \ALU.regsA_result_cry_10_1\
        );

    \I__1661\ : InMux
    port map (
            O => \N__9506\,
            I => \ALU.regsA_result_cry_11\
        );

    \I__1660\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__9497\,
            I => \ALU.regsA_result_cry_11_THRU_CO\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__1656\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__9485\,
            I => \ALU.regsA_result_axb_10_l_ofx\
        );

    \I__1653\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__9479\,
            I => \N__9476\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__9473\,
            I => \ALU.addsub_3\
        );

    \I__1649\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9467\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__1647\ : Odrv12
    port map (
            O => \N__9464\,
            I => \ALU.mult_3\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__1645\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__9449\,
            I => res_11
        );

    \I__1641\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__9443\,
            I => res_3
        );

    \I__1639\ : IoInMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1637\ : IoSpan4Mux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__1636\ : Span4Mux_s3_h
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1635\ : Sp12to4
    port map (
            O => \N__9428\,
            I => \N__9424\
        );

    \I__1634\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9421\
        );

    \I__1633\ : Span12Mux_s10_h
    port map (
            O => \N__9424\,
            I => \N__9418\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__1631\ : Odrv12
    port map (
            O => \N__9418\,
            I => \GPIO1_c\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__9415\,
            I => \GPIO1_c\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__1628\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__9401\,
            I => res_9
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__1624\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__9392\,
            I => \N__9389\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__9389\,
            I => res_12
        );

    \I__1621\ : CEMux
    port map (
            O => \N__9386\,
            I => \N__9382\
        );

    \I__1620\ : CEMux
    port map (
            O => \N__9385\,
            I => \N__9379\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__9382\,
            I => \TXstate_fast_RNIP6NA1_3\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__9379\,
            I => \TXstate_fast_RNIP6NA1_3\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__1616\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__9368\,
            I => \ALU.mult_AdderTree2_bigtree_832\
        );

    \I__1614\ : InMux
    port map (
            O => \N__9365\,
            I => \ALU.regsA_result_cry_2_4\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__1612\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__9356\,
            I => \ALU.mult_AdderTree2_bigtree_833\
        );

    \I__1610\ : InMux
    port map (
            O => \N__9353\,
            I => \ALU.regsA_result_cry_3_5\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__1608\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__9344\,
            I => \ALU.mult_AdderTree2_bigtree_834\
        );

    \I__1606\ : InMux
    port map (
            O => \N__9341\,
            I => \ALU.regsA_result_cry_4_4\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__1604\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__9332\,
            I => \ALU.mult_AdderTree2_bigtree_835\
        );

    \I__1602\ : InMux
    port map (
            O => \N__9329\,
            I => \ALU.regsA_result_cry_5_5\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__1600\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__9320\,
            I => \ALU.mult_AdderTree2_bigtree_836\
        );

    \I__1598\ : InMux
    port map (
            O => \N__9317\,
            I => \ALU.regsA_result_cry_6_4\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__1596\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__9308\,
            I => \ALU.mult_AdderTree2_bigtree_837\
        );

    \I__1594\ : InMux
    port map (
            O => \N__9305\,
            I => \ALU.regsA_result_cry_7_4\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__9296\,
            I => \ALU.mult_AdderTree2_bigtree_838\
        );

    \I__1590\ : InMux
    port map (
            O => \N__9293\,
            I => \ALU.regsA_result_cry_8_1\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__9284\,
            I => \ALU.mult_AdderTree2_bigtree_839\
        );

    \I__1586\ : InMux
    port map (
            O => \N__9281\,
            I => \bfn_13_16_0_\
        );

    \I__1585\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__9275\,
            I => \ALU.mult_AdderTree2_bigtree_538\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__1582\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__9263\,
            I => \ALU.mult_AdderTree2_bigtree_571\
        );

    \I__1579\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__9257\,
            I => \ALU.mult_AdderTree2_bigtree_802\
        );

    \I__1577\ : InMux
    port map (
            O => \N__9254\,
            I => \bfn_13_14_0_\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__9248\,
            I => \ALU.mult_AdderTree2_bigtree_539\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__9236\,
            I => \ALU.mult_AdderTree2_bigtree_572\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__9230\,
            I => \ALU.mult_AdderTree2_bigtree_803\
        );

    \I__1568\ : InMux
    port map (
            O => \N__9227\,
            I => \ALU.regsA_result_cry_8_0\
        );

    \I__1567\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9221\,
            I => \ALU.mult_AdderTree2_bigtree_540\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__9212\,
            I => \N__9209\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__9209\,
            I => \ALU.mult_AdderTree2_bigtree_573\
        );

    \I__1561\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__9197\,
            I => \ALU.mult_AdderTree2_bigtree_804\
        );

    \I__1557\ : InMux
    port map (
            O => \N__9194\,
            I => \ALU.regsA_result_cry_9_1\
        );

    \I__1556\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__9188\,
            I => \ALU.mult_AdderTree2_bigtree_541\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__1553\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__9176\,
            I => \ALU.mult_AdderTree2_bigtree_574\
        );

    \I__1550\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__9167\,
            I => \ALU.mult_AdderTree2_bigtree_805\
        );

    \I__1547\ : InMux
    port map (
            O => \N__9164\,
            I => \ALU.regsA_result_cry_10_0\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__9158\,
            I => \ALU.mult_AdderTree2_bigtree_542\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__1543\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__9146\,
            I => \ALU.mult_AdderTree2_bigtree_575\
        );

    \I__1540\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__9137\,
            I => \ALU.mult_AdderTree2_bigtree_806\
        );

    \I__1537\ : InMux
    port map (
            O => \N__9134\,
            I => \ALU.regsA_result_cry_11_2\
        );

    \I__1536\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__9128\,
            I => \ALU.mult_AdderTree2_bigtree_543\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__1533\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__1531\ : Span4Mux_h
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__9113\,
            I => \ALU.mult_AdderTree2_bigtree_576\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__1528\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__9101\,
            I => \ALU.mult_AdderTree2_bigtree_807\
        );

    \I__1525\ : InMux
    port map (
            O => \N__9098\,
            I => \ALU.regsA_result_cry_12\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__9092\,
            I => \ALU.regsA_result_axb_14\
        );

    \I__1522\ : InMux
    port map (
            O => \N__9089\,
            I => \ALU.regsA_result_cry_13\
        );

    \I__1521\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__9080\,
            I => \ALU.regsA_result_axb_12_0\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__9071\,
            I => \ALU.mult_AdderTree2_bigtree_531\
        );

    \I__1515\ : InMux
    port map (
            O => \N__9068\,
            I => \ALU.regsA_result_cry_0_1\
        );

    \I__1514\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__9062\,
            I => \ALU.mult_AdderTree2_bigtree_532\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__1511\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__9050\,
            I => \ALU.mult_AdderTree2_bigtree_565\
        );

    \I__1508\ : InMux
    port map (
            O => \N__9047\,
            I => \ALU.regsA_result_cry_1_2\
        );

    \I__1507\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__9041\,
            I => \ALU.mult_AdderTree2_bigtree_533\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1504\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__9029\,
            I => \ALU.mult_AdderTree2_bigtree_566\
        );

    \I__1501\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__9020\,
            I => \ALU.mult_AdderTree2_bigtree_797\
        );

    \I__1498\ : InMux
    port map (
            O => \N__9017\,
            I => \ALU.regsA_result_cry_2_3\
        );

    \I__1497\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__9011\,
            I => \ALU.mult_AdderTree2_bigtree_534\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__1494\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__8999\,
            I => \ALU.mult_AdderTree2_bigtree_567\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__8990\,
            I => \ALU.mult_AdderTree2_bigtree_798\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8987\,
            I => \ALU.regsA_result_cry_3_3\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__8981\,
            I => \ALU.mult_AdderTree2_bigtree_535\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__1484\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__8969\,
            I => \ALU.mult_AdderTree2_bigtree_568\
        );

    \I__1481\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__1479\ : Span12Mux_v
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__1478\ : Odrv12
    port map (
            O => \N__8957\,
            I => \ALU.mult_AdderTree2_bigtree_799\
        );

    \I__1477\ : InMux
    port map (
            O => \N__8954\,
            I => \ALU.regsA_result_cry_4_2\
        );

    \I__1476\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__8948\,
            I => \ALU.mult_AdderTree2_bigtree_536\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1473\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__8936\,
            I => \ALU.mult_AdderTree2_bigtree_569\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__8927\,
            I => \ALU.mult_AdderTree2_bigtree_800\
        );

    \I__1467\ : InMux
    port map (
            O => \N__8924\,
            I => \ALU.regsA_result_cry_5_3\
        );

    \I__1466\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__8918\,
            I => \ALU.mult_AdderTree2_bigtree_537\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1461\ : Odrv12
    port map (
            O => \N__8906\,
            I => \ALU.mult_AdderTree2_bigtree_570\
        );

    \I__1460\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__8894\,
            I => \ALU.mult_AdderTree2_bigtree_801\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8891\,
            I => \ALU.regsA_result_cry_6_2\
        );

    \I__1455\ : InMux
    port map (
            O => \N__8888\,
            I => \ALU.regsA_result_cry_7_7\
        );

    \I__1454\ : InMux
    port map (
            O => \N__8885\,
            I => \bfn_13_12_0_\
        );

    \I__1453\ : InMux
    port map (
            O => \N__8882\,
            I => \ALU.regsA_result_cry_9_5\
        );

    \I__1452\ : InMux
    port map (
            O => \N__8879\,
            I => \ALU.regsA_result_cry_10_4\
        );

    \I__1451\ : InMux
    port map (
            O => \N__8876\,
            I => \ALU.regsA_result_cry_11_4\
        );

    \I__1450\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__8867\,
            I => \ALU.regsA_result_cry_13_ma_0\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__1446\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__8855\,
            I => \ALU.regsA_result_axb_13_l_ofx_0\
        );

    \I__1443\ : InMux
    port map (
            O => \N__8852\,
            I => \ALU.regsA_result_cry_12_1\
        );

    \I__1442\ : InMux
    port map (
            O => \N__8849\,
            I => \ALU.regsA_result_cry_13_0\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1440\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__8840\,
            I => \ALU.regsA_result_cry_13_0_THRU_CO\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__8834\,
            I => \ALU.regsA_result_cry_12_ma_0\
        );

    \I__1436\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__8828\,
            I => \ALU.regsA_result_cry_0_0_c_RNO_0\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1432\ : Odrv4
    port map (
            O => \N__8819\,
            I => \ALU.regsA_result_cry_12_ma\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1430\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__8807\,
            I => \ALU.regsA_result_axb_13_l_ofx\
        );

    \I__1427\ : InMux
    port map (
            O => \N__8804\,
            I => \ALU.regsA_result_cry_1_8\
        );

    \I__1426\ : InMux
    port map (
            O => \N__8801\,
            I => \ALU.regsA_result_cry_2_10\
        );

    \I__1425\ : InMux
    port map (
            O => \N__8798\,
            I => \ALU.regsA_result_cry_3_10\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__8789\,
            I => \ALU.regsA_result_cry_5_ma_3\
        );

    \I__1421\ : InMux
    port map (
            O => \N__8786\,
            I => \ALU.regsA_result_cry_4_9\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8783\,
            I => \ALU.regsA_result_cry_5_9\
        );

    \I__1419\ : InMux
    port map (
            O => \N__8780\,
            I => \ALU.regsA_result_cry_6_8\
        );

    \I__1418\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__1416\ : Odrv12
    port map (
            O => \N__8771\,
            I => res_6
        );

    \I__1415\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__8765\,
            I => res_14
        );

    \I__1413\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__1411\ : Odrv12
    port map (
            O => \N__8756\,
            I => res_15
        );

    \I__1410\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__8750\,
            I => res_7
        );

    \I__1408\ : InMux
    port map (
            O => \N__8747\,
            I => \N__8740\
        );

    \I__1407\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8736\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__8745\,
            I => \N__8733\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__8744\,
            I => \N__8730\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__8743\,
            I => \N__8727\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__8740\,
            I => \N__8724\
        );

    \I__1402\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8720\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8716\
        );

    \I__1400\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8709\
        );

    \I__1399\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8709\
        );

    \I__1398\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8709\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__8724\,
            I => \N__8706\
        );

    \I__1396\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8703\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8700\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__8719\,
            I => \N__8693\
        );

    \I__1393\ : Span4Mux_h
    port map (
            O => \N__8716\,
            I => \N__8686\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8686\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__8706\,
            I => \N__8683\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__8703\,
            I => \N__8678\
        );

    \I__1389\ : Span4Mux_h
    port map (
            O => \N__8700\,
            I => \N__8678\
        );

    \I__1388\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8675\
        );

    \I__1387\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8662\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8662\
        );

    \I__1385\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8662\
        );

    \I__1384\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8662\
        );

    \I__1383\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8662\
        );

    \I__1382\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8662\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__8686\,
            I => \aZ0Z_11\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__8683\,
            I => \aZ0Z_11\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__8678\,
            I => \aZ0Z_11\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__8675\,
            I => \aZ0Z_11\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__8662\,
            I => \aZ0Z_11\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1375\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__8636\,
            I => \ALU.addsub_axb_11_l_ofxZ0\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__1369\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1367\ : Span4Mux_v
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__8621\,
            I => \ALU.regsA_result_axb_12_l_ofx\
        );

    \I__1365\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__8612\,
            I => \ALU.regsA_result_cry_11_ma\
        );

    \I__1362\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__8603\,
            I => \N__8599\
        );

    \I__1359\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8596\
        );

    \I__1358\ : Span4Mux_v
    port map (
            O => \N__8599\,
            I => \N__8591\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__8596\,
            I => \N__8591\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__8591\,
            I => \ALU.mult_AdderTree2_bigtree_938\
        );

    \I__1355\ : InMux
    port map (
            O => \N__8588\,
            I => \ALU.regsA_result_cry_9_0\
        );

    \I__1354\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8578\
        );

    \I__1352\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8575\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__8578\,
            I => \N__8572\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__8575\,
            I => \N__8569\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__8572\,
            I => \N__8564\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__8569\,
            I => \N__8564\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__8564\,
            I => \ALU.mult_AdderTree2_bigtree_939\
        );

    \I__1346\ : InMux
    port map (
            O => \N__8561\,
            I => \ALU.regsA_result_cry_10\
        );

    \I__1345\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1343\ : Span4Mux_h
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__8546\,
            I => \ALU.regsA_result_axb_8\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1339\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__8531\,
            I => \ALU.regsA_result_cry_7_THRU_CO\
        );

    \I__1335\ : InMux
    port map (
            O => \N__8528\,
            I => \ALU.regsA_result_cry_11_0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__8516\,
            I => \ALU.regsA_result_axb_8_0\
        );

    \I__1330\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__8510\,
            I => \ALU.mult_5\
        );

    \I__1328\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__8501\,
            I => \ALU.addsub_5\
        );

    \I__1325\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__8492\,
            I => \ALU.addsub_7\
        );

    \I__1322\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__8486\,
            I => \ALU.mult_7\
        );

    \I__1320\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__8480\,
            I => overflow
        );

    \I__1318\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__8471\,
            I => \N_91\
        );

    \I__1315\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__8465\,
            I => res_13
        );

    \I__1313\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__8459\,
            I => res_5
        );

    \I__1311\ : IoInMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__1309\ : IoSpan4Mux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__1308\ : Span4Mux_s3_h
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1307\ : Span4Mux_h
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__1306\ : Span4Mux_h
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1305\ : Sp12to4
    port map (
            O => \N__8438\,
            I => \N__8434\
        );

    \I__1304\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8431\
        );

    \I__1303\ : Span12Mux_v
    port map (
            O => \N__8434\,
            I => \N__8426\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__8431\,
            I => \N__8426\
        );

    \I__1301\ : Odrv12
    port map (
            O => \N__8426\,
            I => \GPIO2_c\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1299\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__8417\,
            I => res_10
        );

    \I__1297\ : InMux
    port map (
            O => \N__8414\,
            I => \ALU.regsA_result_cry_0\
        );

    \I__1296\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__8402\,
            I => \ALU.mult_6\
        );

    \I__1292\ : InMux
    port map (
            O => \N__8399\,
            I => \ALU.regsA_result_cry_1_0\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8396\,
            I => \ALU.regsA_result_cry_2_1\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1289\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__8387\,
            I => \N__8383\
        );

    \I__1287\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8380\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__8383\,
            I => \N__8377\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__8380\,
            I => \ALU.mult_AdderTree2_bigtree_932\
        );

    \I__1284\ : Odrv4
    port map (
            O => \N__8377\,
            I => \ALU.mult_AdderTree2_bigtree_932\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8372\,
            I => \ALU.regsA_result_cry_3_1\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__1281\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8363\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__8363\,
            I => \N__8360\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__8357\,
            I => \ALU.mult_AdderTree2_bigtree_933\
        );

    \I__1277\ : InMux
    port map (
            O => \N__8354\,
            I => \ALU.regsA_result_cry_4_0\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__8351\,
            I => \N__8347\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__8350\,
            I => \N__8344\
        );

    \I__1274\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8341\
        );

    \I__1273\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8338\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8335\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8332\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__8335\,
            I => \N__8329\
        );

    \I__1269\ : Span4Mux_h
    port map (
            O => \N__8332\,
            I => \N__8326\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__8329\,
            I => \ALU.mult_AdderTree2_bigtree_934\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__8326\,
            I => \ALU.mult_AdderTree2_bigtree_934\
        );

    \I__1266\ : InMux
    port map (
            O => \N__8321\,
            I => \ALU.regsA_result_cry_5_1\
        );

    \I__1265\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8314\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__8317\,
            I => \N__8311\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8308\
        );

    \I__1262\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8305\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__8305\,
            I => \N__8299\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__8302\,
            I => \N__8296\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__8299\,
            I => \N__8293\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__8296\,
            I => \ALU.mult_AdderTree2_bigtree_935\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__8293\,
            I => \ALU.mult_AdderTree2_bigtree_935\
        );

    \I__1255\ : InMux
    port map (
            O => \N__8288\,
            I => \ALU.regsA_result_cry_6_0\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__1253\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8278\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__8281\,
            I => \N__8275\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__8278\,
            I => \N__8272\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8269\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__8272\,
            I => \N__8266\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__8269\,
            I => \N__8263\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__8266\,
            I => \ALU.mult_AdderTree2_bigtree_936\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__8263\,
            I => \ALU.mult_AdderTree2_bigtree_936\
        );

    \I__1245\ : InMux
    port map (
            O => \N__8258\,
            I => \bfn_12_16_0_\
        );

    \I__1244\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8251\
        );

    \I__1243\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__8248\,
            I => \N__8242\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__8245\,
            I => \N__8239\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__8242\,
            I => \N__8236\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__8239\,
            I => \ALU.mult_AdderTree2_bigtree_937\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__8236\,
            I => \ALU.mult_AdderTree2_bigtree_937\
        );

    \I__1236\ : InMux
    port map (
            O => \N__8231\,
            I => \ALU.regsA_result_cry_8\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__8225\,
            I => \ALU.regsA_result_axb_14_l_ofx\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1232\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__8216\,
            I => \ALU.addsub_axb_7_l_ofxZ0\
        );

    \I__1230\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8210\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1228\ : Odrv12
    port map (
            O => \N__8207\,
            I => \ALU.regsA_result_cry_8_ma\
        );

    \I__1227\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__8201\,
            I => \ALU.regsA_result_axb_14_0\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1224\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__8192\,
            I => \ALU.regsA_result_cry_14_ma\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1221\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__8183\,
            I => \ALU.addsub_axb_1_l_ofxZ0\
        );

    \I__1219\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8177\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__8177\,
            I => \N__8173\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__8176\,
            I => \N__8170\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__8173\,
            I => \N__8165\
        );

    \I__1215\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8158\
        );

    \I__1214\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8158\
        );

    \I__1213\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8158\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__8165\,
            I => \N__8155\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__8158\,
            I => \N__8152\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__8155\,
            I => \bZ0Z_15\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__8152\,
            I => \bZ0Z_15\
        );

    \I__1208\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__8144\,
            I => \ALU.overflow_RNOZ0Z_15\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__1205\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__8135\,
            I => \ALU.addsub_axb_0_l_ofxZ0\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__8132\,
            I => \N__8129\
        );

    \I__1202\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8126\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__8126\,
            I => \ALU.regsA_result_axb_7_l_ofx\
        );

    \I__1200\ : InMux
    port map (
            O => \N__8123\,
            I => \ALU.regsA_result_cry_6_5\
        );

    \I__1199\ : InMux
    port map (
            O => \N__8120\,
            I => \bfn_12_13_0_\
        );

    \I__1198\ : InMux
    port map (
            O => \N__8117\,
            I => \ALU.regsA_result_cry_8_2\
        );

    \I__1197\ : InMux
    port map (
            O => \N__8114\,
            I => \ALU.regsA_result_cry_9_3\
        );

    \I__1196\ : InMux
    port map (
            O => \N__8111\,
            I => \ALU.regsA_result_cry_10_2\
        );

    \I__1195\ : InMux
    port map (
            O => \N__8108\,
            I => \ALU.regsA_result_cry_11_3\
        );

    \I__1194\ : InMux
    port map (
            O => \N__8105\,
            I => \ALU.regsA_result_cry_12_0\
        );

    \I__1193\ : InMux
    port map (
            O => \N__8102\,
            I => \ALU.regsA_result_cry_13_1\
        );

    \I__1192\ : InMux
    port map (
            O => \N__8099\,
            I => \ALU.regsA_result_cry_14\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1190\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__8090\,
            I => \ALU.regsA_result_cry_0_0_c_RNO\
        );

    \I__1188\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__8084\,
            I => \ALU.regsA_result_axb_1_l_ofx\
        );

    \I__1186\ : InMux
    port map (
            O => \N__8081\,
            I => \ALU.regsA_result_cry_0_2\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1184\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__8072\,
            I => \ALU.regsA_result_axb_2_l_ofx\
        );

    \I__1182\ : InMux
    port map (
            O => \N__8069\,
            I => \ALU.regsA_result_cry_1_3\
        );

    \I__1181\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__8063\,
            I => \ALU.regsA_result_cry_3_ma\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1178\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__8054\,
            I => \ALU.regsA_result_axb_3_l_ofx\
        );

    \I__1176\ : InMux
    port map (
            O => \N__8051\,
            I => \ALU.regsA_result_cry_2_5\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1174\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__8042\,
            I => \ALU.regsA_result_axb_4_l_ofx\
        );

    \I__1172\ : InMux
    port map (
            O => \N__8039\,
            I => \ALU.regsA_result_cry_3_6\
        );

    \I__1171\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__8033\,
            I => \ALU.regsA_result_axb_5_l_ofx\
        );

    \I__1169\ : InMux
    port map (
            O => \N__8030\,
            I => \ALU.regsA_result_cry_4_5\
        );

    \I__1168\ : InMux
    port map (
            O => \N__8027\,
            I => \ALU.regsA_result_cry_5_6\
        );

    \I__1167\ : InMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__8018\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_2\
        );

    \I__1164\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__8006\,
            I => \ALU.regsA_result_cry_2_ma_2\
        );

    \I__1160\ : InMux
    port map (
            O => \N__8003\,
            I => \N__8000\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__7997\,
            I => \ALU.regsA_result_cry_3_ma_2\
        );

    \I__1157\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__7988\,
            I => \ALU.regsA_result_cry_4_ma_1\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7981\
        );

    \I__1153\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7978\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__7981\,
            I => \N__7973\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7970\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__7977\,
            I => \N__7967\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__7976\,
            I => \N__7964\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__7973\,
            I => \N__7957\
        );

    \I__1147\ : Span4Mux_h
    port map (
            O => \N__7970\,
            I => \N__7957\
        );

    \I__1146\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7954\
        );

    \I__1145\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7949\
        );

    \I__1144\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7949\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__7962\,
            I => \N__7946\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__7957\,
            I => \N__7942\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__7954\,
            I => \N__7939\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7936\
        );

    \I__1139\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7931\
        );

    \I__1138\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7931\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__7942\,
            I => \aZ0Z_14\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__7939\,
            I => \aZ0Z_14\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__7936\,
            I => \aZ0Z_14\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__7931\,
            I => \aZ0Z_14\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__7910\,
            I => \ALU.addsub_axb_14_l_ofxZ0\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__7907\,
            I => \N__7903\
        );

    \I__1127\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7900\
        );

    \I__1126\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7897\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__7900\,
            I => \N__7892\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7897\,
            I => \N__7889\
        );

    \I__1123\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7886\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__7895\,
            I => \N__7883\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__7892\,
            I => \N__7870\
        );

    \I__1120\ : Span4Mux_h
    port map (
            O => \N__7889\,
            I => \N__7870\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7870\
        );

    \I__1118\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7865\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7865\
        );

    \I__1116\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7862\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__7880\,
            I => \N__7859\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \N__7856\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__7878\,
            I => \N__7852\
        );

    \I__1112\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7848\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__7870\,
            I => \N__7843\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__7865\,
            I => \N__7843\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7840\
        );

    \I__1108\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7829\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7829\
        );

    \I__1106\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7829\
        );

    \I__1105\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7829\
        );

    \I__1104\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7829\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7848\,
            I => \aZ0Z_8\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__7843\,
            I => \aZ0Z_8\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__7840\,
            I => \aZ0Z_8\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__7829\,
            I => \aZ0Z_8\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1098\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__1096\ : Span4Mux_v
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__7808\,
            I => \ALU.addsub_axb_8_l_ofxZ0\
        );

    \I__1094\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__7799\,
            I => \N__7796\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__7796\,
            I => \ALU.addsub_axb_9_l_ofxZ0\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__7793\,
            I => \N__7790\
        );

    \I__1089\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7785\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7782\
        );

    \I__1087\ : InMux
    port map (
            O => \N__7788\,
            I => \N__7778\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__7785\,
            I => \N__7775\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__7782\,
            I => \N__7772\
        );

    \I__1084\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7769\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__7778\,
            I => \N__7764\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__7775\,
            I => \N__7751\
        );

    \I__1081\ : Span4Mux_h
    port map (
            O => \N__7772\,
            I => \N__7751\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__7769\,
            I => \N__7751\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__7768\,
            I => \N__7744\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__7767\,
            I => \N__7740\
        );

    \I__1077\ : Span12Mux_s11_h
    port map (
            O => \N__7764\,
            I => \N__7736\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7725\
        );

    \I__1075\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7725\
        );

    \I__1074\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7725\
        );

    \I__1073\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7725\
        );

    \I__1072\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7725\
        );

    \I__1071\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7722\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__7751\,
            I => \N__7719\
        );

    \I__1069\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7714\
        );

    \I__1068\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7714\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7701\
        );

    \I__1066\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7701\
        );

    \I__1065\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7701\
        );

    \I__1064\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7701\
        );

    \I__1063\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7701\
        );

    \I__1062\ : InMux
    port map (
            O => \N__7739\,
            I => \N__7701\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__7736\,
            I => \aZ0Z_9\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__7725\,
            I => \aZ0Z_9\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__7722\,
            I => \aZ0Z_9\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__7719\,
            I => \aZ0Z_9\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7714\,
            I => \aZ0Z_9\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__7701\,
            I => \aZ0Z_9\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1054\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__7682\,
            I => \ALU.regsA_result_cry_5_ma_1\
        );

    \I__1052\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7676\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__7676\,
            I => \ALU.addsub_15\
        );

    \I__1050\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__7670\,
            I => \ALU.mult_15\
        );

    \I__1048\ : InMux
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__7658\,
            I => \ALU.addsub_6\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__7655\,
            I => \ALU.mult_2_cascade_\
        );

    \I__1043\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1041\ : Span4Mux_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__7643\,
            I => \ALU.addsub_2\
        );

    \I__1039\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7634\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__7634\,
            I => \ALU.regsA_result_cry_7_ma_0\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1035\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__7625\,
            I => \ALU.regsA_result_axb_7_l_ofx_0\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1032\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__7616\,
            I => \ALU.regsA_result_axb_8_1\
        );

    \I__1030\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7609\
        );

    \I__1029\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7606\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7603\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1026\ : Span4Mux_h
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__7600\,
            I => \ALU.mult_ab_128\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__7597\,
            I => \ALU.mult_ab_128\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1022\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__7586\,
            I => \ALU.addsub_8\
        );

    \I__1020\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__7574\,
            I => res_8
        );

    \I__1016\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__7568\,
            I => \ALU.addsub_11\
        );

    \I__1014\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__7562\,
            I => \ALU.mult_11\
        );

    \I__1012\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__7553\,
            I => \ALU.addsub_0\
        );

    \I__1009\ : IoInMux
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__7547\,
            I => \N__7543\
        );

    \I__1007\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7540\
        );

    \I__1006\ : Span12Mux_s4_v
    port map (
            O => \N__7543\,
            I => \N__7537\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__7540\,
            I => \N__7534\
        );

    \I__1004\ : Span12Mux_v
    port map (
            O => \N__7537\,
            I => \N__7531\
        );

    \I__1003\ : Span4Mux_h
    port map (
            O => \N__7534\,
            I => \N__7528\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__7531\,
            I => \GPIO0_c\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__7528\,
            I => \GPIO0_c\
        );

    \I__1000\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__7520\,
            I => \ALU.addsub_13\
        );

    \I__998\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__7514\,
            I => \ALU.mult_13\
        );

    \I__996\ : InMux
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__7505\,
            I => \ALU.addsub_12\
        );

    \I__993\ : InMux
    port map (
            O => \N__7502\,
            I => \N__7499\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__7499\,
            I => \ALU.mult_12\
        );

    \I__991\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__7493\,
            I => \ALU.mult_1\
        );

    \I__989\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__7484\,
            I => \ALU.addsub_1\
        );

    \I__986\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__7475\,
            I => \ALU.addsub_9\
        );

    \I__983\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__7469\,
            I => \ALU.mult_9\
        );

    \I__981\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__7460\,
            I => \ALU.addsub_10\
        );

    \I__978\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__7454\,
            I => \ALU.mult_10\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__7451\,
            I => \N__7447\
        );

    \I__975\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7442\
        );

    \I__974\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7437\
        );

    \I__973\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7437\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__7445\,
            I => \N__7432\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__7442\,
            I => \N__7427\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__7437\,
            I => \N__7427\
        );

    \I__969\ : InMux
    port map (
            O => \N__7436\,
            I => \N__7422\
        );

    \I__968\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7422\
        );

    \I__967\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7416\
        );

    \I__966\ : Sp12to4
    port map (
            O => \N__7427\,
            I => \N__7411\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__7422\,
            I => \N__7411\
        );

    \I__964\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7404\
        );

    \I__963\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7404\
        );

    \I__962\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7404\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__7416\,
            I => \aZ0Z_10\
        );

    \I__960\ : Odrv12
    port map (
            O => \N__7411\,
            I => \aZ0Z_10\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__7404\,
            I => \aZ0Z_10\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__957\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7391\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__7391\,
            I => \ALU.addsub_axb_10_l_ofxZ0\
        );

    \I__955\ : InMux
    port map (
            O => \N__7388\,
            I => \ALU.addsub_cry_9\
        );

    \I__954\ : InMux
    port map (
            O => \N__7385\,
            I => \ALU.addsub_cry_10\
        );

    \I__953\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7378\
        );

    \I__952\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7375\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__7378\,
            I => \N__7369\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7366\
        );

    \I__949\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7363\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__7373\,
            I => \N__7358\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__7372\,
            I => \N__7354\
        );

    \I__946\ : Span4Mux_v
    port map (
            O => \N__7369\,
            I => \N__7350\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__7366\,
            I => \N__7345\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__7363\,
            I => \N__7345\
        );

    \I__943\ : InMux
    port map (
            O => \N__7362\,
            I => \N__7342\
        );

    \I__942\ : InMux
    port map (
            O => \N__7361\,
            I => \N__7339\
        );

    \I__941\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7334\
        );

    \I__940\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7334\
        );

    \I__939\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7329\
        );

    \I__938\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7329\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__7350\,
            I => \aZ0Z_12\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__7345\,
            I => \aZ0Z_12\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__7342\,
            I => \aZ0Z_12\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__7339\,
            I => \aZ0Z_12\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7334\,
            I => \aZ0Z_12\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__7329\,
            I => \aZ0Z_12\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__7316\,
            I => \N__7313\
        );

    \I__930\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__928\ : Odrv12
    port map (
            O => \N__7307\,
            I => \ALU.addsub_axb_12_l_ofxZ0\
        );

    \I__927\ : InMux
    port map (
            O => \N__7304\,
            I => \ALU.addsub_cry_11\
        );

    \I__926\ : InMux
    port map (
            O => \N__7301\,
            I => \ALU.addsub_cry_12\
        );

    \I__925\ : InMux
    port map (
            O => \N__7298\,
            I => \ALU.addsub_cry_13\
        );

    \I__924\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7291\
        );

    \I__923\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7286\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7283\
        );

    \I__921\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7276\
        );

    \I__920\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7276\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7273\
        );

    \I__918\ : Span12Mux_v
    port map (
            O => \N__7283\,
            I => \N__7270\
        );

    \I__917\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7265\
        );

    \I__916\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7265\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7262\
        );

    \I__914\ : Odrv12
    port map (
            O => \N__7273\,
            I => \aZ0Z_15\
        );

    \I__913\ : Odrv12
    port map (
            O => \N__7270\,
            I => \aZ0Z_15\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__7265\,
            I => \aZ0Z_15\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__7262\,
            I => \aZ0Z_15\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \N__7250\
        );

    \I__909\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__7244\,
            I => \ALU.addsub_axb_15_l_ofxZ0\
        );

    \I__906\ : InMux
    port map (
            O => \N__7241\,
            I => \bfn_11_16_0_\
        );

    \I__905\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__7235\,
            I => \ALU.mult_16\
        );

    \I__903\ : InMux
    port map (
            O => \N__7232\,
            I => \ALU.addsub_cry_15\
        );

    \I__902\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__7226\,
            I => \ALU.addsub_14\
        );

    \I__900\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__7220\,
            I => \ALU.mult_14\
        );

    \I__898\ : InMux
    port map (
            O => \N__7217\,
            I => \ALU.addsub_cry_0\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__896\ : InMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__7208\,
            I => \ALU.addsub_axb_2_l_ofxZ0\
        );

    \I__894\ : InMux
    port map (
            O => \N__7205\,
            I => \ALU.addsub_cry_1\
        );

    \I__893\ : InMux
    port map (
            O => \N__7202\,
            I => \ALU.addsub_cry_2\
        );

    \I__892\ : InMux
    port map (
            O => \N__7199\,
            I => \ALU.addsub_cry_3\
        );

    \I__891\ : InMux
    port map (
            O => \N__7196\,
            I => \ALU.addsub_cry_4\
        );

    \I__890\ : InMux
    port map (
            O => \N__7193\,
            I => \ALU.addsub_cry_5\
        );

    \I__889\ : InMux
    port map (
            O => \N__7190\,
            I => \bfn_11_15_0_\
        );

    \I__888\ : InMux
    port map (
            O => \N__7187\,
            I => \ALU.addsub_cry_7\
        );

    \I__887\ : InMux
    port map (
            O => \N__7184\,
            I => \ALU.addsub_cry_8\
        );

    \I__886\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7178\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7178\,
            I => \ALU.regsA_result_axb_6\
        );

    \I__884\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7172\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__7172\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_0\
        );

    \I__882\ : InMux
    port map (
            O => \N__7169\,
            I => \ALU.addsub_cry_0_c_THRU_CO\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__880\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7160\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__7160\,
            I => \ALU.regsA_result_axb_6_l_ofx_0\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__877\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__7151\,
            I => \ALU.mult_AdderTree2_bigtree_674\
        );

    \I__875\ : InMux
    port map (
            O => \N__7148\,
            I => \ALU.regsA_result_cry_5_7\
        );

    \I__874\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7142\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__7142\,
            I => \ALU.mult_AdderTree2_bigtree_675\
        );

    \I__872\ : InMux
    port map (
            O => \N__7139\,
            I => \ALU.regsA_result_cry_6_6\
        );

    \I__871\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__7133\,
            I => \ALU.regsA_result_cry_5_0_THRU_CO\
        );

    \I__869\ : InMux
    port map (
            O => \N__7130\,
            I => \ALU.regsA_result_cry_7_0\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__7127\,
            I => \N__7124\
        );

    \I__867\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__7121\,
            I => \ALU.regsA_result_axb_8_2\
        );

    \I__865\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7112\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__7112\,
            I => \ALU.regsA_result_cry_6_ma_0\
        );

    \I__862\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__7106\,
            I => \N__7101\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__7105\,
            I => \N__7098\
        );

    \I__859\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7095\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__7101\,
            I => \N__7092\
        );

    \I__857\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7089\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__7095\,
            I => \ALU.mult_AdderTree2_bigtree_670\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__7092\,
            I => \ALU.mult_AdderTree2_bigtree_670\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__7089\,
            I => \ALU.mult_AdderTree2_bigtree_670\
        );

    \I__853\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__7076\,
            I => \ALU.regsA_result_cry_2_c_RNO_0\
        );

    \I__850\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__7070\,
            I => \ALU.regsA_result_cry_3_ma_0\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__7067\,
            I => \N__7064\
        );

    \I__847\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__7061\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_1\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__844\ : InMux
    port map (
            O => \N__7055\,
            I => \N__7052\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__7052\,
            I => \ALU.regsA_result_axb_2_l_ofx_2\
        );

    \I__842\ : InMux
    port map (
            O => \N__7049\,
            I => \ALU.regsA_result_cry_1_6\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__840\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__7040\,
            I => \ALU.regsA_result_axb_3_l_ofx_2\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__837\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__7031\,
            I => \ALU.mult_AdderTree2_bigtree_671\
        );

    \I__835\ : InMux
    port map (
            O => \N__7028\,
            I => \ALU.regsA_result_cry_2_8\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__833\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__7019\,
            I => \ALU.regsA_result_axb_4_l_ofx_1\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__830\ : InMux
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__7010\,
            I => \ALU.mult_AdderTree2_bigtree_672\
        );

    \I__828\ : InMux
    port map (
            O => \N__7007\,
            I => \ALU.regsA_result_cry_3_8\
        );

    \I__827\ : InMux
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__6998\,
            I => \ALU.regsA_result_axb_5_l_ofx_1\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__823\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6989\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__6989\,
            I => \ALU.mult_AdderTree2_bigtree_673\
        );

    \I__821\ : InMux
    port map (
            O => \N__6986\,
            I => \ALU.regsA_result_cry_4_7\
        );

    \I__820\ : InMux
    port map (
            O => \N__6983\,
            I => \bfn_10_17_0_\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__818\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6973\
        );

    \I__817\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__6973\,
            I => \a_fastZ0Z_10\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__6970\,
            I => \a_fastZ0Z_10\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__6965\,
            I => \N__6962\
        );

    \I__813\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6959\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__6959\,
            I => \ALU.regsA_result_axb_2_l_ofx_1\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__6956\,
            I => \N__6953\
        );

    \I__810\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__6950\,
            I => \ALU.regsA_result_axb_3_l_ofx_1\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__807\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6941\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__6941\,
            I => \N__6938\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__6938\,
            I => \ALU.regsA_result_axb_5_l_ofx_0\
        );

    \I__804\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__6932\,
            I => \N__6929\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__6929\,
            I => \ALU.mult_AdderTree2_bigtree_669\
        );

    \I__801\ : InMux
    port map (
            O => \N__6926\,
            I => \ALU.regsA_result_cry_0_0\
        );

    \I__800\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__798\ : Span4Mux_h
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__797\ : Odrv4
    port map (
            O => \N__6914\,
            I => \ALU.regsA_result_cry_5_c_RNI073QE\
        );

    \I__796\ : InMux
    port map (
            O => \N__6911\,
            I => \ALU.regsA_result_cry_1_1\
        );

    \I__795\ : InMux
    port map (
            O => \N__6908\,
            I => \N__6905\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__6902\,
            I => \ALU.regsA_result_cry_2_c_RNIHNOEF\
        );

    \I__792\ : InMux
    port map (
            O => \N__6899\,
            I => \ALU.regsA_result_cry_2_2\
        );

    \I__791\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__6893\,
            I => \ALU.regsA_result_cry_7_c_RNI8EG3H\
        );

    \I__789\ : InMux
    port map (
            O => \N__6890\,
            I => \ALU.regsA_result_cry_3_2\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__787\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__6881\,
            I => \N__6878\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__6875\,
            I => \ALU.regsA_result_cry_4_c_RNIA939H\
        );

    \I__783\ : InMux
    port map (
            O => \N__6872\,
            I => \ALU.regsA_result_cry_4_1\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__6869\,
            I => \N__6866\
        );

    \I__781\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__779\ : Span4Mux_v
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__6857\,
            I => \ALU.regsA_result_cry_5_c_RNIKCNNP\
        );

    \I__777\ : InMux
    port map (
            O => \N__6854\,
            I => \ALU.regsA_result_cry_5_2\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__775\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__6839\,
            I => \ALU.regsA_result_cry_6_c_RNICICNO\
        );

    \I__771\ : InMux
    port map (
            O => \N__6836\,
            I => \ALU.regsA_result_cry_6_1\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__6833\,
            I => \N__6829\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__6832\,
            I => \N__6826\
        );

    \I__768\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6818\
        );

    \I__767\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6818\
        );

    \I__766\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6818\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__6818\,
            I => \FTDI.baudAccZ0Z_0\
        );

    \I__764\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6809\
        );

    \I__763\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6809\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__6806\,
            I => \FTDI.baudAccZ0Z_1\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__6803\,
            I => \FTDI.N_170_0_cascade_\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__6800\,
            I => \FTDI.TXstate_cnst_0_0_2_cascade_\
        );

    \I__758\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6793\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__6796\,
            I => \N__6789\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6786\
        );

    \I__755\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6781\
        );

    \I__754\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6781\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__6786\,
            I => \ALU.mult_AdderTree2_bigtree_870\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__6781\,
            I => \ALU.mult_AdderTree2_bigtree_870\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__6776\,
            I => \N__6772\
        );

    \I__750\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6765\
        );

    \I__749\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6758\
        );

    \I__748\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6758\
        );

    \I__747\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6758\
        );

    \I__746\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6753\
        );

    \I__745\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6753\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__6765\,
            I => \FTDI.TXstateZ0Z_1\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__6758\,
            I => \FTDI.TXstateZ0Z_1\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__6753\,
            I => \FTDI.TXstateZ0Z_1\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__6746\,
            I => \N__6742\
        );

    \I__740\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6739\
        );

    \I__739\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6736\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__6739\,
            I => \FTDI.TXstate_fastZ0Z_3\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__6736\,
            I => \FTDI.TXstate_fastZ0Z_3\
        );

    \I__736\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6714\
        );

    \I__735\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6714\
        );

    \I__734\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6714\
        );

    \I__733\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6714\
        );

    \I__732\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6714\
        );

    \I__731\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6709\
        );

    \I__730\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6709\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__6714\,
            I => \FTDI.TXstateZ0Z_0\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__6709\,
            I => \FTDI.TXstateZ0Z_0\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__6704\,
            I => \FTDI_TXready_cascade_\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__6701\,
            I => \un1_testState31_0_cascade_\
        );

    \I__725\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6695\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__6695\,
            I => \ALU.mult_AdderTree2_bigtree_741\
        );

    \I__723\ : InMux
    port map (
            O => \N__6692\,
            I => \ALU.regsA_result_cry_2_6\
        );

    \I__722\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__720\ : Span4Mux_h
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__6680\,
            I => \ALU.regsA_result_axb_2\
        );

    \I__718\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__6671\,
            I => \ALU.regsA_result_cry_1_THRU_CO\
        );

    \I__715\ : InMux
    port map (
            O => \N__6668\,
            I => \ALU.regsA_result_cry_3\
        );

    \I__714\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6662\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__6659\,
            I => \ALU.regsA_result_axb_4_0\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__710\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__6650\,
            I => \ALU.regsA_result_axb_3_l_ofx_0\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__707\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__6641\,
            I => \ALU.regsA_result_axb_4\
        );

    \I__705\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6634\
        );

    \I__704\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6631\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__6634\,
            I => \ALU.mult_AdderTree2_bigtree_873\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__6631\,
            I => \ALU.mult_AdderTree2_bigtree_873\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__700\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__6620\,
            I => \ALU.regsA_result_cry_2_c_RNIC59KA\
        );

    \I__698\ : InMux
    port map (
            O => \N__6617\,
            I => \ALU.regsA_result_cry_2\
        );

    \I__697\ : InMux
    port map (
            O => \N__6614\,
            I => \ALU.regsA_result_cry_3_0\
        );

    \I__696\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__6608\,
            I => \ALU.regsA_result_cry_3_0_THRU_CO\
        );

    \I__694\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__6602\,
            I => \ALU.mult_AdderTree2_bigtree_739\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__691\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__6593\,
            I => \ALU.mult_AdderTree2_bigtree_774\
        );

    \I__689\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__6587\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_3\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__686\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__6578\,
            I => \ALU.regsA_result_cry_1_0_c_RNO\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__683\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__6569\,
            I => \ALU.regsA_result_axb_2_l_ofx_0\
        );

    \I__681\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6559\
        );

    \I__680\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6559\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__6564\,
            I => \N__6556\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__677\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__6553\,
            I => \ALU.mult_AdderTree2_bigtree_740\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__6550\,
            I => \ALU.mult_AdderTree2_bigtree_740\
        );

    \I__674\ : InMux
    port map (
            O => \N__6545\,
            I => \ALU.regsA_result_cry_1_4\
        );

    \I__673\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6539\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__6539\,
            I => \ALU.regsA_result_cry_5_ma_0\
        );

    \I__671\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__6533\,
            I => \N__6530\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__6530\,
            I => \ALU.mult_AdderTree2_bigtree_704\
        );

    \I__668\ : InMux
    port map (
            O => \N__6527\,
            I => \ALU.regsA_result_cry_2_0\
        );

    \I__667\ : InMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__6521\,
            I => \ALU.mult_AdderTree2_bigtree_705\
        );

    \I__665\ : InMux
    port map (
            O => \N__6518\,
            I => \ALU.regsA_result_cry_3_4\
        );

    \I__664\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__6509\,
            I => \ALU.mult_AdderTree2_bigtree_706\
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__6506\,
            I => \N__6503\
        );

    \I__660\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__6500\,
            I => \ALU.mult_AdderTree2_bigtree_871\
        );

    \I__658\ : InMux
    port map (
            O => \N__6497\,
            I => \ALU.regsA_result_cry_4_3\
        );

    \I__657\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__6491\,
            I => \ALU.mult_AdderTree2_bigtree_707\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__6488\,
            I => \N__6484\
        );

    \I__654\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6481\
        );

    \I__653\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6478\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__6481\,
            I => \ALU.mult_AdderTree2_bigtree_872\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__6478\,
            I => \ALU.mult_AdderTree2_bigtree_872\
        );

    \I__650\ : InMux
    port map (
            O => \N__6473\,
            I => \ALU.regsA_result_cry_5_4\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__648\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__6464\,
            I => \ALU.mult_AdderTree2_bigtree_708\
        );

    \I__646\ : InMux
    port map (
            O => \N__6461\,
            I => \ALU.regsA_result_cry_6_3\
        );

    \I__645\ : InMux
    port map (
            O => \N__6458\,
            I => \ALU.regsA_result_cry_7_1\
        );

    \I__644\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__6452\,
            I => \ALU.regsA_result_cry_2_c_RNO\
        );

    \I__642\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__6446\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__6443\,
            I => \N__6440\
        );

    \I__639\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6437\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__6437\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_0_1\
        );

    \I__637\ : InMux
    port map (
            O => \N__6434\,
            I => \N__6431\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__6431\,
            I => \N__6428\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__6428\,
            I => \ALU.regsA_result_cry_2_ma_1\
        );

    \I__634\ : InMux
    port map (
            O => \N__6425\,
            I => \ALU.regsA_result_cry_1_5\
        );

    \I__633\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6419\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__6416\,
            I => \ALU.regsA_result_cry_3_ma_1\
        );

    \I__630\ : InMux
    port map (
            O => \N__6413\,
            I => \ALU.regsA_result_cry_2_7\
        );

    \I__629\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__6407\,
            I => \ALU.regsA_result_cry_4_ma_0\
        );

    \I__627\ : InMux
    port map (
            O => \N__6404\,
            I => \ALU.regsA_result_cry_3_7\
        );

    \I__626\ : InMux
    port map (
            O => \N__6401\,
            I => \ALU.regsA_result_cry_4_6\
        );

    \I__625\ : InMux
    port map (
            O => \N__6398\,
            I => \ALU.regsA_result_cry_5_0\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__623\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__6389\,
            I => \ALU.regsA_result_axb_4_l_ofx_0\
        );

    \I__621\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6383\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__6383\,
            I => \FTDI.TXstate_RNIE1MMZ0Z_2\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__6380\,
            I => \FTDI.TXstate_RNIE1MMZ0Z_2_cascade_\
        );

    \I__618\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__6374\,
            I => \ALU.regsA_result_cry_4_c_RNO\
        );

    \I__616\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__6368\,
            I => \ALU.regsA_result_cry_1_0_c_RNIKGQO9\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__6365\,
            I => \FTDI.i2_mux_cascade_\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__6362\,
            I => \N__6359\
        );

    \I__612\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6356\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__6356\,
            I => \ALU.regsA_result_cry_1_0_c_RNO_2\
        );

    \I__610\ : InMux
    port map (
            O => \N__6353\,
            I => \ALU.regsA_result_cry_1\
        );

    \I__609\ : InMux
    port map (
            O => \N__6350\,
            I => \ALU.regsA_result_cry_4\
        );

    \I__608\ : InMux
    port map (
            O => \N__6347\,
            I => \ALU.regsA_result_cry_5\
        );

    \I__607\ : InMux
    port map (
            O => \N__6344\,
            I => \ALU.regsA_result_cry_6\
        );

    \I__606\ : InMux
    port map (
            O => \N__6341\,
            I => \ALU.regsA_result_cry_7\
        );

    \I__605\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__6335\,
            I => \clkdivZ0Z_17\
        );

    \I__603\ : InMux
    port map (
            O => \N__6332\,
            I => clkdiv_cry_16
        );

    \I__602\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__6326\,
            I => \clkdivZ0Z_18\
        );

    \I__600\ : InMux
    port map (
            O => \N__6323\,
            I => clkdiv_cry_17
        );

    \I__599\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__6317\,
            I => \clkdivZ0Z_19\
        );

    \I__597\ : InMux
    port map (
            O => \N__6314\,
            I => clkdiv_cry_18
        );

    \I__596\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__6308\,
            I => \clkdivZ0Z_20\
        );

    \I__594\ : InMux
    port map (
            O => \N__6305\,
            I => clkdiv_cry_19
        );

    \I__593\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6299\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__6299\,
            I => \clkdivZ0Z_21\
        );

    \I__591\ : InMux
    port map (
            O => \N__6296\,
            I => clkdiv_cry_20
        );

    \I__590\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__6290\,
            I => \clkdivZ0Z_22\
        );

    \I__588\ : InMux
    port map (
            O => \N__6287\,
            I => clkdiv_cry_21
        );

    \I__587\ : InMux
    port map (
            O => \N__6284\,
            I => clkdiv_cry_22
        );

    \I__586\ : IoInMux
    port map (
            O => \N__6281\,
            I => \N__6278\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__584\ : Span12Mux_s10_v
    port map (
            O => \N__6275\,
            I => \N__6271\
        );

    \I__583\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6268\
        );

    \I__582\ : Odrv12
    port map (
            O => \N__6271\,
            I => \GPIO3_c\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__6268\,
            I => \GPIO3_c\
        );

    \I__580\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6260\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__6260\,
            I => \clkdivZ0Z_8\
        );

    \I__578\ : InMux
    port map (
            O => \N__6257\,
            I => \bfn_1_14_0_\
        );

    \I__577\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__6251\,
            I => \clkdivZ0Z_9\
        );

    \I__575\ : InMux
    port map (
            O => \N__6248\,
            I => clkdiv_cry_8
        );

    \I__574\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__6242\,
            I => \clkdivZ0Z_10\
        );

    \I__572\ : InMux
    port map (
            O => \N__6239\,
            I => clkdiv_cry_9
        );

    \I__571\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__6233\,
            I => \clkdivZ0Z_11\
        );

    \I__569\ : InMux
    port map (
            O => \N__6230\,
            I => clkdiv_cry_10
        );

    \I__568\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6224\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__6224\,
            I => \clkdivZ0Z_12\
        );

    \I__566\ : InMux
    port map (
            O => \N__6221\,
            I => clkdiv_cry_11
        );

    \I__565\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__6215\,
            I => \clkdivZ0Z_13\
        );

    \I__563\ : InMux
    port map (
            O => \N__6212\,
            I => clkdiv_cry_12
        );

    \I__562\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__6206\,
            I => \clkdivZ0Z_14\
        );

    \I__560\ : InMux
    port map (
            O => \N__6203\,
            I => clkdiv_cry_13
        );

    \I__559\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__6197\,
            I => \clkdivZ0Z_15\
        );

    \I__557\ : InMux
    port map (
            O => \N__6194\,
            I => clkdiv_cry_14
        );

    \I__556\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__6188\,
            I => \clkdivZ0Z_16\
        );

    \I__554\ : InMux
    port map (
            O => \N__6185\,
            I => \bfn_1_15_0_\
        );

    \I__553\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6179\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__6179\,
            I => \clkdivZ0Z_0\
        );

    \I__551\ : InMux
    port map (
            O => \N__6176\,
            I => \bfn_1_13_0_\
        );

    \I__550\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__6170\,
            I => \clkdivZ0Z_1\
        );

    \I__548\ : InMux
    port map (
            O => \N__6167\,
            I => clkdiv_cry_0
        );

    \I__547\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6161\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__6161\,
            I => \clkdivZ0Z_2\
        );

    \I__545\ : InMux
    port map (
            O => \N__6158\,
            I => clkdiv_cry_1
        );

    \I__544\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__6152\,
            I => \clkdivZ0Z_3\
        );

    \I__542\ : InMux
    port map (
            O => \N__6149\,
            I => clkdiv_cry_2
        );

    \I__541\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6143\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__6143\,
            I => \clkdivZ0Z_4\
        );

    \I__539\ : InMux
    port map (
            O => \N__6140\,
            I => clkdiv_cry_3
        );

    \I__538\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__6134\,
            I => \clkdivZ0Z_5\
        );

    \I__536\ : InMux
    port map (
            O => \N__6131\,
            I => clkdiv_cry_4
        );

    \I__535\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6125\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__6125\,
            I => \clkdivZ0Z_6\
        );

    \I__533\ : InMux
    port map (
            O => \N__6122\,
            I => clkdiv_cry_5
        );

    \I__532\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6116\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__6116\,
            I => \clkdivZ0Z_7\
        );

    \I__530\ : InMux
    port map (
            O => \N__6113\,
            I => clkdiv_cry_6
        );

    \INVFTDI.gap_1C\ : INV
    port map (
            O => \INVFTDI.gap_1C_net\,
            I => \N__16076\
        );

    \INVFTDI.RXstate_2C\ : INV
    port map (
            O => \INVFTDI.RXstate_2C_net\,
            I => \N__16074\
        );

    \INVFTDI.RXstate_3C\ : INV
    port map (
            O => \INVFTDI.RXstate_3C_net\,
            I => \N__16073\
        );

    \INVFTDI.TXshift_7C\ : INV
    port map (
            O => \INVFTDI.TXshift_7C_net\,
            I => \N__16110\
        );

    \INVFTDI.RXbuffer_5C\ : INV
    port map (
            O => \INVFTDI.RXbuffer_5C_net\,
            I => \N__16078\
        );

    \INVFTDI.RXbuffer_2C\ : INV
    port map (
            O => \INVFTDI.RXbuffer_2C_net\,
            I => \N__16075\
        );

    \INVFTDI.TXshift_1C\ : INV
    port map (
            O => \INVFTDI.TXshift_1C_net\,
            I => \N__16112\
        );

    \INVFTDI.TXstate_2C\ : INV
    port map (
            O => \INVFTDI.TXstate_2C_net\,
            I => \N__16117\
        );

    \INVFTDI.baudAcc_0C\ : INV
    port map (
            O => \INVFTDI.baudAcc_0C_net\,
            I => \N__16113\
        );

    \INVFTDI.TXstate_0C\ : INV
    port map (
            O => \INVFTDI.TXstate_0C_net\,
            I => \N__16121\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.addsub_cry_6\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.addsub_cry_14\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_7_9\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_7_2\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_9_2\,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_7_3\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_8_5\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_8_3\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_8_4\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.regsA_result_cry_7_5\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_7,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_15,
            carryinitout => \bfn_1_15_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \clkdiv_0_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6182\,
            in2 => \_gnd_net_\,
            in3 => \N__6176\,
            lcout => \clkdivZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => clkdiv_cry_0,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_1_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6173\,
            in2 => \_gnd_net_\,
            in3 => \N__6167\,
            lcout => \clkdivZ0Z_1\,
            ltout => OPEN,
            carryin => clkdiv_cry_0,
            carryout => clkdiv_cry_1,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_2_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6164\,
            in2 => \_gnd_net_\,
            in3 => \N__6158\,
            lcout => \clkdivZ0Z_2\,
            ltout => OPEN,
            carryin => clkdiv_cry_1,
            carryout => clkdiv_cry_2,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_3_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6155\,
            in2 => \_gnd_net_\,
            in3 => \N__6149\,
            lcout => \clkdivZ0Z_3\,
            ltout => OPEN,
            carryin => clkdiv_cry_2,
            carryout => clkdiv_cry_3,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_4_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6146\,
            in2 => \_gnd_net_\,
            in3 => \N__6140\,
            lcout => \clkdivZ0Z_4\,
            ltout => OPEN,
            carryin => clkdiv_cry_3,
            carryout => clkdiv_cry_4,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_5_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6137\,
            in2 => \_gnd_net_\,
            in3 => \N__6131\,
            lcout => \clkdivZ0Z_5\,
            ltout => OPEN,
            carryin => clkdiv_cry_4,
            carryout => clkdiv_cry_5,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_6_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6128\,
            in2 => \_gnd_net_\,
            in3 => \N__6122\,
            lcout => \clkdivZ0Z_6\,
            ltout => OPEN,
            carryin => clkdiv_cry_5,
            carryout => clkdiv_cry_6,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_7_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6119\,
            in2 => \_gnd_net_\,
            in3 => \N__6113\,
            lcout => \clkdivZ0Z_7\,
            ltout => OPEN,
            carryin => clkdiv_cry_6,
            carryout => clkdiv_cry_7,
            clk => \N__16122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_8_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6263\,
            in2 => \_gnd_net_\,
            in3 => \N__6257\,
            lcout => \clkdivZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => clkdiv_cry_8,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_9_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6254\,
            in2 => \_gnd_net_\,
            in3 => \N__6248\,
            lcout => \clkdivZ0Z_9\,
            ltout => OPEN,
            carryin => clkdiv_cry_8,
            carryout => clkdiv_cry_9,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_10_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6245\,
            in2 => \_gnd_net_\,
            in3 => \N__6239\,
            lcout => \clkdivZ0Z_10\,
            ltout => OPEN,
            carryin => clkdiv_cry_9,
            carryout => clkdiv_cry_10,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_11_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6236\,
            in2 => \_gnd_net_\,
            in3 => \N__6230\,
            lcout => \clkdivZ0Z_11\,
            ltout => OPEN,
            carryin => clkdiv_cry_10,
            carryout => clkdiv_cry_11,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_12_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6227\,
            in2 => \_gnd_net_\,
            in3 => \N__6221\,
            lcout => \clkdivZ0Z_12\,
            ltout => OPEN,
            carryin => clkdiv_cry_11,
            carryout => clkdiv_cry_12,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_13_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6218\,
            in2 => \_gnd_net_\,
            in3 => \N__6212\,
            lcout => \clkdivZ0Z_13\,
            ltout => OPEN,
            carryin => clkdiv_cry_12,
            carryout => clkdiv_cry_13,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_14_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6209\,
            in2 => \_gnd_net_\,
            in3 => \N__6203\,
            lcout => \clkdivZ0Z_14\,
            ltout => OPEN,
            carryin => clkdiv_cry_13,
            carryout => clkdiv_cry_14,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_15_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6200\,
            in2 => \_gnd_net_\,
            in3 => \N__6194\,
            lcout => \clkdivZ0Z_15\,
            ltout => OPEN,
            carryin => clkdiv_cry_14,
            carryout => clkdiv_cry_15,
            clk => \N__16123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_16_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6191\,
            in2 => \_gnd_net_\,
            in3 => \N__6185\,
            lcout => \clkdivZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => clkdiv_cry_16,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_17_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6338\,
            in2 => \_gnd_net_\,
            in3 => \N__6332\,
            lcout => \clkdivZ0Z_17\,
            ltout => OPEN,
            carryin => clkdiv_cry_16,
            carryout => clkdiv_cry_17,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_18_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6329\,
            in2 => \_gnd_net_\,
            in3 => \N__6323\,
            lcout => \clkdivZ0Z_18\,
            ltout => OPEN,
            carryin => clkdiv_cry_17,
            carryout => clkdiv_cry_18,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_19_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6320\,
            in2 => \_gnd_net_\,
            in3 => \N__6314\,
            lcout => \clkdivZ0Z_19\,
            ltout => OPEN,
            carryin => clkdiv_cry_18,
            carryout => clkdiv_cry_19,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_20_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6311\,
            in2 => \_gnd_net_\,
            in3 => \N__6305\,
            lcout => \clkdivZ0Z_20\,
            ltout => OPEN,
            carryin => clkdiv_cry_19,
            carryout => clkdiv_cry_20,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_21_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6302\,
            in2 => \_gnd_net_\,
            in3 => \N__6296\,
            lcout => \clkdivZ0Z_21\,
            ltout => OPEN,
            carryin => clkdiv_cry_20,
            carryout => clkdiv_cry_21,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_22_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6293\,
            in2 => \_gnd_net_\,
            in3 => \N__6287\,
            lcout => \clkdivZ0Z_22\,
            ltout => OPEN,
            carryin => clkdiv_cry_21,
            carryout => clkdiv_cry_22,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_23_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6274\,
            in2 => \_gnd_net_\,
            in3 => \N__6284\,
            lcout => \GPIO3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_14_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14318\,
            lcout => \aZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16108\,
            ce => \N__12244\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__7282\,
            in1 => \N__7945\,
            in2 => \N__13783\,
            in3 => \N__12025\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_8_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__12026\,
            in1 => \N__7281\,
            in2 => \N__7962\,
            in3 => \N__11833\,
            lcout => \ALU.regsA_result_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_15_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12119\,
            lcout => \aZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16108\,
            ce => \N__12244\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6590\,
            in2 => \N__6362\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \ALU.regsA_result_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_1_THRU_LUT4_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6353\,
            lcout => \ALU.regsA_result_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6377\,
            in2 => \N__6796\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \ALU.regsA_result_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNIA939H_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__8255\,
            in1 => \N__6605\,
            in2 => \N__6506\,
            in3 => \N__6350\,
            lcout => \ALU.regsA_result_cry_4_c_RNIA939H\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4\,
            carryout => \ALU.regsA_result_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_5_c_RNIKCNNP_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__8609\,
            in1 => \N__6371\,
            in2 => \N__6488\,
            in3 => \N__6347\,
            lcout => \ALU.regsA_result_cry_5_c_RNIKCNNP\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5\,
            carryout => \ALU.regsA_result_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_6_c_RNICICNO_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__8585\,
            in1 => \N__6637\,
            in2 => \N__6626\,
            in3 => \N__6344\,
            lcout => \ALU.regsA_result_cry_6_c_RNICICNO\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6\,
            carryout => \ALU.regsA_result_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_7_THRU_LUT4_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6341\,
            lcout => \ALU.regsA_result_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_2_regsA_result_cry_4_c_RNO_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7361\,
            in1 => \N__6792\,
            in2 => \_gnd_net_\,
            in3 => \N__13724\,
            lcout => \ALU.regsA_result_cry_4_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNIKGQO9_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001101100"
        )
    port map (
            in0 => \N__13725\,
            in1 => \N__6565\,
            in2 => \N__7976\,
            in3 => \N__6487\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNIKGQO9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNO_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__6566\,
            in1 => \N__7963\,
            in2 => \_gnd_net_\,
            in3 => \N__13723\,
            lcout => \ALU.regsA_result_cry_2_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_12_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10970\,
            lcout => \aZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16116\,
            ce => \N__12242\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__13782\,
            in1 => \N__14660\,
            in2 => \N__12067\,
            in3 => \N__7353\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_2_l_ofx_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__12057\,
            in1 => \N__14659\,
            in2 => \N__7372\,
            in3 => \N__11831\,
            lcout => \ALU.regsA_result_axb_2_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_0_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001111"
        )
    port map (
            in0 => \N__14020\,
            in1 => \N__6770\,
            in2 => \N__15388\,
            in3 => \N__6727\,
            lcout => OPEN,
            ltout => \FTDI.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__6728\,
            in1 => \_gnd_net_\,
            in2 => \N__6365\,
            in3 => \N__12745\,
            lcout => \FTDI.TXstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_fast_3_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000100"
        )
    port map (
            in0 => \N__6731\,
            in1 => \N__6386\,
            in2 => \N__6776\,
            in3 => \N__6745\,
            lcout => \FTDI.TXstate_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNIE1MM_2_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12741\,
            in2 => \_gnd_net_\,
            in3 => \N__14019\,
            lcout => \FTDI.TXstate_RNIE1MMZ0Z_2\,
            ltout => \FTDI.TXstate_RNIE1MMZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_3_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100010000"
        )
    port map (
            in0 => \N__6730\,
            in1 => \N__6775\,
            in2 => \N__6380\,
            in3 => \N__15377\,
            lcout => \FTDI.TXstateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_1_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010011000100"
        )
    port map (
            in0 => \N__12744\,
            in1 => \N__6771\,
            in2 => \N__15389\,
            in3 => \N__6729\,
            lcout => \FTDI.TXstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_15_l_ofx_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__14464\,
            in1 => \N__8180\,
            in2 => \_gnd_net_\,
            in3 => \N__7294\,
            lcout => \ALU.addsub_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_RNO_0_0_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7583\,
            in1 => \N__7546\,
            in2 => \_gnd_net_\,
            in3 => \N__15914\,
            lcout => \N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_1_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__8697\,
            in1 => \N__13768\,
            in2 => \N__6980\,
            in3 => \N__12062\,
            lcout => \ALU.mult_AdderTree2_bigtree_704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__8698\,
            in1 => \N__13769\,
            in2 => \N__12066\,
            in3 => \N__6976\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_11_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10427\,
            lcout => \aZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16099\,
            ce => \N__12241\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNO_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__8691\,
            in1 => \N__13767\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_ma_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8692\,
            in2 => \_gnd_net_\,
            in3 => \N__12053\,
            lcout => \ALU.regsA_result_cry_2_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_ma_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11824\,
            in1 => \_gnd_net_\,
            in2 => \N__8719\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_3_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_ma_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8696\,
            in2 => \_gnd_net_\,
            in3 => \N__13344\,
            lcout => \ALU.regsA_result_cry_4_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6449\,
            in2 => \N__6443\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \ALU.regsA_result_cry_1_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_1_0_c_RNI2J0N2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6434\,
            in2 => \N__6965\,
            in3 => \N__6425\,
            lcout => \ALU.mult_AdderTree2_bigtree_705\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_5\,
            carryout => \ALU.regsA_result_cry_2_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_2_0_c_RNI6Q6R2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6422\,
            in2 => \N__6956\,
            in3 => \N__6413\,
            lcout => \ALU.mult_AdderTree2_bigtree_706\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_7\,
            carryout => \ALU.regsA_result_cry_3_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_3_0_c_RNIA1DV2_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6410\,
            in2 => \N__6395\,
            in3 => \N__6404\,
            lcout => \ALU.mult_AdderTree2_bigtree_707\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_7\,
            carryout => \ALU.regsA_result_cry_4_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_4_0_c_RNIE8JJ2_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6542\,
            in2 => \N__6947\,
            in3 => \N__6401\,
            lcout => \ALU.mult_AdderTree2_bigtree_708\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_6\,
            carryout => \ALU.regsA_result_cry_5_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_5_0_THRU_LUT4_0_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6398\,
            lcout => \ALU.regsA_result_cry_5_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_4_l_ofx_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11657\,
            in1 => \N__8723\,
            in2 => \N__7445\,
            in3 => \N__13317\,
            lcout => \ALU.regsA_result_axb_4_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_cry_5_ma_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11658\,
            in2 => \_gnd_net_\,
            in3 => \N__8699\,
            lcout => \ALU.regsA_result_cry_5_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7082\,
            in2 => \N__7105\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \ALU.regsA_result_cry_2_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNIHNOEF_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__8318\,
            in1 => \N__6536\,
            in2 => \N__7037\,
            in3 => \N__6527\,
            lcout => \ALU.regsA_result_cry_2_c_RNIHNOEF\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_0\,
            carryout => \ALU.regsA_result_cry_3_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_3_c_RNIHID36_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6524\,
            in2 => \N__7016\,
            in3 => \N__6518\,
            lcout => \ALU.mult_AdderTree2_bigtree_870\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_4\,
            carryout => \ALU.regsA_result_cry_4_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_4_c_RNIQ2RR5_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6515\,
            in2 => \N__6995\,
            in3 => \N__6497\,
            lcout => \ALU.mult_AdderTree2_bigtree_871\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_3\,
            carryout => \ALU.regsA_result_cry_5_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_5_c_RNI3J846_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6494\,
            in2 => \N__7157\,
            in3 => \N__6473\,
            lcout => \ALU.mult_AdderTree2_bigtree_872\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_4\,
            carryout => \ALU.regsA_result_cry_6_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_6_c_RNIC3MS5_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7145\,
            in2 => \N__6470\,
            in3 => \N__6461\,
            lcout => \ALU.mult_AdderTree2_bigtree_873\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_3\,
            carryout => \ALU.regsA_result_cry_7_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_2_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6611\,
            in1 => \N__6665\,
            in2 => \N__7127\,
            in3 => \N__6458\,
            lcout => \ALU.regsA_result_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6455\,
            in2 => \N__6564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \ALU.regsA_result_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_4_regsA_result_cry_2_c_RNIC59KA_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__6638\,
            in1 => \N__6698\,
            in2 => \N__6599\,
            in3 => \N__6617\,
            lcout => \ALU.regsA_result_cry_2_c_RNIC59KA\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2\,
            carryout => \ALU.regsA_result_cry_3_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_3_0_THRU_LUT4_0_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6614\,
            lcout => \ALU.regsA_result_cry_3_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_1_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__12064\,
            in1 => \N__7362\,
            in2 => \N__13766\,
            in3 => \N__14648\,
            lcout => \ALU.mult_AdderTree2_bigtree_739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_axb_1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__7290\,
            in1 => \N__13717\,
            in2 => \N__7977\,
            in3 => \N__12063\,
            lcout => \ALU.mult_AdderTree2_bigtree_774\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_8_regsA_result_cry_1_0_c_RNO_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13716\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_5_l_ofx_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__7788\,
            in1 => \N__11661\,
            in2 => \N__15041\,
            in3 => \N__7881\,
            lcout => \ALU.regsA_result_axb_5_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7175\,
            in2 => \N__6584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \ALU.regsA_result_cry_1_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNI9GUP2_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11138\,
            in2 => \N__6575\,
            in3 => \N__6545\,
            lcout => \ALU.mult_AdderTree2_bigtree_740\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_4\,
            carryout => \ALU.regsA_result_cry_2_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_0_c_RNIDN4U2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7073\,
            in2 => \N__6656\,
            in3 => \N__6692\,
            lcout => \ALU.mult_AdderTree2_bigtree_741\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_6\,
            carryout => \ALU.regsA_result_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_4_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6689\,
            in1 => \N__6677\,
            in2 => \N__6647\,
            in3 => \N__6668\,
            lcout => \ALU.regsA_result_axb_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_axb_3_l_ofx_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13342\,
            in1 => \N__7357\,
            in2 => \N__11834\,
            in3 => \N__14656\,
            lcout => \ALU.regsA_result_axb_3_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_9_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__14655\,
            in1 => \N__11659\,
            in2 => \N__7373\,
            in3 => \N__13343\,
            lcout => \ALU.regsA_result_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_FirstStep_AB_1_128_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7896\,
            lcout => \ALU.mult_ab_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_2_l_ofx_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__14446\,
            in1 => \N__11832\,
            in2 => \_gnd_net_\,
            in3 => \N__9803\,
            lcout => \ALU.addsub_axb_2_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_0_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6825\,
            in2 => \_gnd_net_\,
            in3 => \N__16173\,
            lcout => \FTDI.baudAccZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_1_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__16174\,
            in1 => \_gnd_net_\,
            in2 => \N__6832\,
            in3 => \N__6814\,
            lcout => \FTDI.baudAccZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_10_l_ofx_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14447\,
            in1 => \_gnd_net_\,
            in2 => \N__7451\,
            in3 => \N__14161\,
            lcout => \ALU.addsub_axb_10_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_1_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__7789\,
            in1 => \N__13771\,
            in2 => \N__7907\,
            in3 => \N__12048\,
            lcout => \ALU.mult_AdderTree2_bigtree_669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_2_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__16175\,
            in1 => \_gnd_net_\,
            in2 => \N__6833\,
            in3 => \N__6815\,
            lcout => \FTDI.baudAccZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.baudAcc_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNI073QE_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__7109\,
            in1 => \N__7446\,
            in2 => \N__8351\,
            in3 => \N__13770\,
            lcout => \ALU.regsA_result_cry_5_c_RNI073QE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_1_2_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12742\,
            in1 => \N__6769\,
            in2 => \_gnd_net_\,
            in3 => \N__6726\,
            lcout => OPEN,
            ltout => \FTDI.N_170_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_RNO_0_2_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001011111"
        )
    port map (
            in0 => \N__15381\,
            in1 => \N__12743\,
            in2 => \N__6803\,
            in3 => \N__14018\,
            lcout => OPEN,
            ltout => \FTDI.TXstate_cnst_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12689\,
            in2 => \N__6800\,
            in3 => \N__16172\,
            lcout => \FTDI.un3_TX_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXstate_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNI8EG3H_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__7374\,
            in1 => \N__13780\,
            in2 => \N__8285\,
            in3 => \N__6797\,
            lcout => \ALU.regsA_result_cry_7_c_RNI8EG3H\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_fast_RNIRJI91_3_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14017\,
            in1 => \N__6768\,
            in2 => \N__6746\,
            in3 => \N__6725\,
            lcout => \FTDI_TXready\,
            ltout => \FTDI_TXready_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXstart_esr_RNO_0_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__15778\,
            in1 => \N__15661\,
            in2 => \N__6704\,
            in3 => \N__15902\,
            lcout => OPEN,
            ltout => \un1_testState31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXstart_esr_RNO_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__15947\,
            in1 => \_gnd_net_\,
            in2 => \N__6701\,
            in3 => \_gnd_net_\,
            lcout => \un1_testState31_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_4_m1_forloop_1_1_regsA_result_cry_0_c_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7613\,
            in2 => \N__8393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \ALU.regsA_result_cry_0_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_9_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6935\,
            in2 => \N__8369\,
            in3 => \N__6926\,
            lcout => \ALU.mult_9\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_0_0\,
            carryout => \ALU.regsA_result_cry_1_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_10_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6923\,
            in2 => \N__8350\,
            in3 => \N__6911\,
            lcout => \ALU.mult_10\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_1\,
            carryout => \ALU.regsA_result_cry_2_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_11_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6908\,
            in2 => \N__8317\,
            in3 => \N__6899\,
            lcout => \ALU.mult_11\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_2\,
            carryout => \ALU.regsA_result_cry_3_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_12_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6896\,
            in2 => \N__8281\,
            in3 => \N__6890\,
            lcout => \ALU.mult_12\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_2\,
            carryout => \ALU.regsA_result_cry_4_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_13_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8254\,
            in2 => \N__6887\,
            in3 => \N__6872\,
            lcout => \ALU.mult_13\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_1\,
            carryout => \ALU.regsA_result_cry_5_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_14_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8602\,
            in2 => \N__6869\,
            in3 => \N__6854\,
            lcout => \ALU.mult_14\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_2\,
            carryout => \ALU.regsA_result_cry_6_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_15_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8581\,
            in2 => \N__6851\,
            in3 => \N__6836\,
            lcout => \ALU.mult_15\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_1\,
            carryout => \ALU.regsA_result_cry_7_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8525\,
            in2 => \_gnd_net_\,
            in3 => \N__6983\,
            lcout => \ALU.mult_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_fast_10_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11095\,
            lcout => \a_fastZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16088\,
            ce => \N__12245\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_2_l_ofx_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__12065\,
            in1 => \N__11825\,
            in2 => \N__8743\,
            in3 => \N__7419\,
            lcout => \ALU.regsA_result_axb_2_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_10_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16094\,
            ce => \N__12199\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_3_l_ofx_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13334\,
            in1 => \N__11826\,
            in2 => \N__8744\,
            in3 => \N__7420\,
            lcout => \ALU.regsA_result_axb_3_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_6_regsA_result_axb_5_l_ofx_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__11611\,
            in1 => \N__7421\,
            in2 => \N__8745\,
            in3 => \N__15039\,
            lcout => \ALU.regsA_result_axb_5_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_8_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14514\,
            lcout => \aZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16100\,
            ce => \N__12243\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__7763\,
            in1 => \N__13744\,
            in2 => \N__12061\,
            in3 => \N__7851\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_2_l_ofx_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__12034\,
            in1 => \N__7759\,
            in2 => \N__7878\,
            in3 => \N__11785\,
            lcout => \ALU.regsA_result_axb_2_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_3_l_ofx_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__7760\,
            in1 => \N__13315\,
            in2 => \N__11814\,
            in3 => \N__7855\,
            lcout => \ALU.regsA_result_axb_3_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_4_l_ofx_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__13316\,
            in1 => \N__7761\,
            in2 => \N__7879\,
            in3 => \N__11602\,
            lcout => \ALU.regsA_result_axb_4_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_6_l_ofx_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15040\,
            in1 => \N__7762\,
            in2 => \N__7880\,
            in3 => \N__13081\,
            lcout => \ALU.regsA_result_axb_6_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8024\,
            in2 => \N__7067\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \ALU.regsA_result_cry_1_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNI6MAO2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8015\,
            in2 => \N__7058\,
            in3 => \N__7049\,
            lcout => \ALU.mult_AdderTree2_bigtree_670\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_6\,
            carryout => \ALU.regsA_result_cry_2_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_0_c_RNIATGS2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8003\,
            in2 => \N__7046\,
            in3 => \N__7028\,
            lcout => \ALU.mult_AdderTree2_bigtree_671\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_8\,
            carryout => \ALU.regsA_result_cry_3_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_0_c_RNIE4N03_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7994\,
            in2 => \N__7025\,
            in3 => \N__7007\,
            lcout => \ALU.mult_AdderTree2_bigtree_672\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_8\,
            carryout => \ALU.regsA_result_cry_4_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_0_c_RNIIBTK2_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7004\,
            in2 => \N__7688\,
            in3 => \N__6986\,
            lcout => \ALU.mult_AdderTree2_bigtree_673\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_7\,
            carryout => \ALU.regsA_result_cry_5_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_0_c_RNIMI3P2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7118\,
            in2 => \N__7166\,
            in3 => \N__7148\,
            lcout => \ALU.mult_AdderTree2_bigtree_674\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_7\,
            carryout => \ALU.regsA_result_cry_6_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_0_c_RNIQP9T2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7640\,
            in2 => \N__7631\,
            in3 => \N__7139\,
            lcout => \ALU.mult_AdderTree2_bigtree_675\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_6\,
            carryout => \ALU.regsA_result_cry_7_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_5_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__7136\,
            in1 => \N__7181\,
            in2 => \N__7622\,
            in3 => \N__7130\,
            lcout => \ALU.regsA_result_axb_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_7_l_ofx_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14867\,
            in1 => \N__13183\,
            in2 => \N__12626\,
            in3 => \N__12844\,
            lcout => \ALU.regsA_result_axb_7_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_12_l_ofx_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__7382\,
            in1 => \N__14459\,
            in2 => \_gnd_net_\,
            in3 => \N__9599\,
            lcout => \ALU.addsub_axb_12_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_2_l_ofx_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14866\,
            in1 => \N__13345\,
            in2 => \N__12625\,
            in3 => \N__11798\,
            lcout => \ALU.regsA_result_axb_2_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_6_ma_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7781\,
            in2 => \_gnd_net_\,
            in3 => \N__15031\,
            lcout => \ALU.regsA_result_cry_6_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_3_regsA_result_cry_2_c_RNO_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13722\,
            in1 => \N__7104\,
            in2 => \_gnd_net_\,
            in3 => \N__7435\,
            lcout => \ALU.regsA_result_cry_2_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_3_ma_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11799\,
            in1 => \_gnd_net_\,
            in2 => \N__14658\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_3_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_10_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__15032\,
            in1 => \N__7436\,
            in2 => \N__13091\,
            in3 => \N__8739\,
            lcout => \ALU.regsA_result_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_1_0_c_RNO_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14644\,
            in1 => \N__13721\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11336\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16109\,
            ce => \N__15295\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__12036\,
            in1 => \N__13755\,
            in2 => \N__14898\,
            in3 => \N__12608\,
            lcout => \ALU.regsA_result_cry_0_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_1_l_ofx_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14876\,
            in1 => \N__11827\,
            in2 => \N__12639\,
            in3 => \N__12035\,
            lcout => \ALU.regsA_result_axb_1_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_3_l_ofx_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14877\,
            in1 => \N__11660\,
            in2 => \N__12640\,
            in3 => \N__13325\,
            lcout => \ALU.regsA_result_axb_3_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_4_l_ofx_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__15038\,
            in1 => \N__11606\,
            in2 => \N__14897\,
            in3 => \N__12615\,
            lcout => \ALU.regsA_result_axb_4_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_5_l_ofx_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14878\,
            in1 => \N__13089\,
            in2 => \N__12641\,
            in3 => \N__15037\,
            lcout => \ALU.regsA_result_axb_5_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_0_c_THRU_CRY_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14448\,
            in2 => \N__14463\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \ALU.addsub_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_0_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14889\,
            in2 => \N__8141\,
            in3 => \N__7169\,
            lcout => \ALU.addsub_0\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_0_c_THRU_CO\,
            carryout => \ALU.addsub_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_1_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12603\,
            in2 => \N__8189\,
            in3 => \N__7217\,
            lcout => \ALU.addsub_1\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_0\,
            carryout => \ALU.addsub_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_2_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9802\,
            in2 => \N__7214\,
            in3 => \N__7205\,
            lcout => \ALU.addsub_2\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_1\,
            carryout => \ALU.addsub_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_3_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13523\,
            in2 => \N__13196\,
            in3 => \N__7202\,
            lcout => \ALU.addsub_3\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_2\,
            carryout => \ALU.addsub_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_4_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10901\,
            in2 => \N__10856\,
            in3 => \N__7199\,
            lcout => \ALU.addsub_4\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_3\,
            carryout => \ALU.addsub_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_5_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15204\,
            in2 => \N__14918\,
            in3 => \N__7196\,
            lcout => \ALU.addsub_5\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_4\,
            carryout => \ALU.addsub_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_6_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13879\,
            in2 => \N__13928\,
            in3 => \N__7193\,
            lcout => \ALU.addsub_6\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_5\,
            carryout => \ALU.addsub_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_7_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12967\,
            in2 => \N__8222\,
            in3 => \N__7190\,
            lcout => \ALU.addsub_7\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \ALU.addsub_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_8_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7906\,
            in2 => \N__7820\,
            in3 => \N__7187\,
            lcout => \ALU.addsub_8\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_7\,
            carryout => \ALU.addsub_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_9_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7805\,
            in2 => \N__7793\,
            in3 => \N__7184\,
            lcout => \ALU.addsub_9\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_8\,
            carryout => \ALU.addsub_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_10_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7450\,
            in2 => \N__7397\,
            in3 => \N__7388\,
            lcout => \ALU.addsub_10\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_9\,
            carryout => \ALU.addsub_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_11_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8747\,
            in2 => \N__8651\,
            in3 => \N__7385\,
            lcout => \ALU.addsub_11\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_10\,
            carryout => \ALU.addsub_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_12_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7381\,
            in2 => \N__7316\,
            in3 => \N__7304\,
            lcout => \ALU.addsub_12\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_11\,
            carryout => \ALU.addsub_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_13_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14657\,
            in2 => \N__14534\,
            in3 => \N__7301\,
            lcout => \ALU.addsub_13\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_12\,
            carryout => \ALU.addsub_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_14_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7984\,
            in2 => \N__7922\,
            in3 => \N__7298\,
            lcout => \ALU.addsub_14\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_13\,
            carryout => \ALU.addsub_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_0_15_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7295\,
            in2 => \N__7253\,
            in3 => \N__7241\,
            lcout => \ALU.addsub_15\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \ALU.addsub_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__11271\,
            in1 => \N__7238\,
            in2 => \N__14465\,
            in3 => \N__7232\,
            lcout => overflow,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_1_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__12049\,
            in1 => \N__12638\,
            in2 => \N__14899\,
            in3 => \N__13781\,
            lcout => \ALU.mult_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_14_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11276\,
            in1 => \N__7229\,
            in2 => \_gnd_net_\,
            in3 => \N__7223\,
            lcout => res_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_8_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__7612\,
            in1 => \N__11278\,
            in2 => \N__7592\,
            in3 => \N__8386\,
            lcout => res_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_11_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11272\,
            in1 => \N__7571\,
            in2 => \_gnd_net_\,
            in3 => \N__7565\,
            lcout => res_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__13784\,
            in1 => \N__7559\,
            in2 => \N__14900\,
            in3 => \N__11277\,
            lcout => \GPIO0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_13_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__7523\,
            in1 => \_gnd_net_\,
            in2 => \N__11285\,
            in3 => \N__7517\,
            lcout => res_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_12_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11280\,
            in1 => \N__7511\,
            in2 => \_gnd_net_\,
            in3 => \N__7502\,
            lcout => res_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_1_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11284\,
            in1 => \N__7496\,
            in2 => \_gnd_net_\,
            in3 => \N__7490\,
            lcout => \GPIO1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_9_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11282\,
            in1 => \N__7481\,
            in2 => \_gnd_net_\,
            in3 => \N__7472\,
            lcout => res_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_10_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11283\,
            in1 => \N__7466\,
            in2 => \_gnd_net_\,
            in3 => \N__7457\,
            lcout => res_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_15_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11281\,
            in1 => \N__7679\,
            in2 => \_gnd_net_\,
            in3 => \N__7673\,
            lcout => res_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_15_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12104\,
            lcout => \bZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16083\,
            ce => \N__14225\,
            sr => \_gnd_net_\
        );

    \ALU.res_6_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11231\,
            in1 => \N__7667\,
            in2 => \_gnd_net_\,
            in3 => \N__8411\,
            lcout => res_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9801\,
            in1 => \N__9829\,
            in2 => \_gnd_net_\,
            in3 => \N__13765\,
            lcout => OPEN,
            ltout => \ALU.mult_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11230\,
            in2 => \N__7655\,
            in3 => \N__7652\,
            lcout => \GPIO2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_ma_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11610\,
            in2 => \_gnd_net_\,
            in3 => \N__13513\,
            lcout => \ALU.regsA_result_cry_5_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_7_ma_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7758\,
            in2 => \_gnd_net_\,
            in3 => \N__13085\,
            lcout => \ALU.regsA_result_cry_7_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_axb_7_l_ofx_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__7748\,
            in1 => \N__12851\,
            in2 => \N__13090\,
            in3 => \N__7882\,
            lcout => \ALU.regsA_result_axb_7_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_11_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__12852\,
            in1 => \N__7747\,
            in2 => \N__7895\,
            in3 => \N__13178\,
            lcout => \ALU.regsA_result_axb_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_9_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11332\,
            lcout => \aZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16095\,
            ce => \N__12231\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_1_0_c_RNO_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13728\,
            in2 => \_gnd_net_\,
            in3 => \N__7739\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_2_ma_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7767\,
            in3 => \N__12033\,
            lcout => \ALU.regsA_result_cry_2_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_3_ma_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11784\,
            in2 => \_gnd_net_\,
            in3 => \N__7743\,
            lcout => \ALU.regsA_result_cry_3_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_4_ma_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13318\,
            in2 => \N__7768\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_4_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_14_l_ofx_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__7985\,
            in1 => \N__14267\,
            in2 => \_gnd_net_\,
            in3 => \N__14457\,
            lcout => \ALU.addsub_axb_14_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_8_l_ofx_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14455\,
            in1 => \N__7877\,
            in2 => \_gnd_net_\,
            in3 => \N__13182\,
            lcout => \ALU.addsub_axb_8_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_9_l_ofx_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__7750\,
            in1 => \N__14456\,
            in2 => \_gnd_net_\,
            in3 => \N__12383\,
            lcout => \ALU.addsub_axb_9_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_5_regsA_result_cry_5_ma_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11586\,
            in2 => \_gnd_net_\,
            in3 => \N__7749\,
            lcout => \ALU.regsA_result_cry_5_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_4_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10955\,
            lcout => \bZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16101\,
            ce => \N__11394\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_ma_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11585\,
            in2 => \_gnd_net_\,
            in3 => \N__14868\,
            lcout => \ALU.regsA_result_cry_3_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8831\,
            in2 => \N__8096\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \ALU.regsA_result_cry_0_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNI9TCO2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8087\,
            in2 => \N__12158\,
            in3 => \N__8081\,
            lcout => \ALU.mult_AdderTree2_bigtree_530\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_0_2\,
            carryout => \ALU.regsA_result_cry_1_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_0_c_RNID4JS2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12131\,
            in2 => \N__8078\,
            in3 => \N__8069\,
            lcout => \ALU.mult_AdderTree2_bigtree_531\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_3\,
            carryout => \ALU.regsA_result_cry_2_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_0_c_RNIHBP03_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8066\,
            in2 => \N__8060\,
            in3 => \N__8051\,
            lcout => \ALU.mult_AdderTree2_bigtree_532\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_5\,
            carryout => \ALU.regsA_result_cry_3_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_3_0_c_RNILIVK2_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9737\,
            in2 => \N__8048\,
            in3 => \N__8039\,
            lcout => \ALU.mult_AdderTree2_bigtree_533\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_6\,
            carryout => \ALU.regsA_result_cry_4_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_0_c_RNIPP5P2_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8036\,
            in2 => \N__9929\,
            in3 => \N__8030\,
            lcout => \ALU.mult_AdderTree2_bigtree_534\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_5\,
            carryout => \ALU.regsA_result_cry_5_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_0_c_RNIT0CT2_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9878\,
            in2 => \N__9944\,
            in3 => \N__8027\,
            lcout => \ALU.mult_AdderTree2_bigtree_535\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_6\,
            carryout => \ALU.regsA_result_cry_6_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_0_c_RNI18I13_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12503\,
            in2 => \N__8132\,
            in3 => \N__8123\,
            lcout => \ALU.mult_AdderTree2_bigtree_536\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_5\,
            carryout => \ALU.regsA_result_cry_7_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_0_c_RNI5FOL2_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8213\,
            in2 => \N__12515\,
            in3 => \N__8120\,
            lcout => \ALU.mult_AdderTree2_bigtree_537\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \ALU.regsA_result_cry_8_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_0_c_RNIN2AT1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14078\,
            in2 => \N__10871\,
            in3 => \N__8117\,
            lcout => \ALU.mult_AdderTree2_bigtree_538\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_8_2\,
            carryout => \ALU.regsA_result_cry_9_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_0_c_RNI206J1_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9626\,
            in2 => \N__9494\,
            in3 => \N__8114\,
            lcout => \ALU.mult_AdderTree2_bigtree_539\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_9_3\,
            carryout => \ALU.regsA_result_cry_10_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_0_c_RNIDUIG1_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8618\,
            in2 => \N__9641\,
            in3 => \N__8111\,
            lcout => \ALU.mult_AdderTree2_bigtree_540\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_10_2\,
            carryout => \ALU.regsA_result_cry_11_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_0_c_RNIH5PK1_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8825\,
            in2 => \N__8633\,
            in3 => \N__8108\,
            lcout => \ALU.mult_AdderTree2_bigtree_541\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_11_3\,
            carryout => \ALU.regsA_result_cry_12_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_0_c_RNILCVO1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14669\,
            in2 => \N__8816\,
            in3 => \N__8105\,
            lcout => \ALU.mult_AdderTree2_bigtree_542\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_12_0\,
            carryout => \ALU.regsA_result_cry_13_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_0_c_RNIPJ5D1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8228\,
            in2 => \N__8198\,
            in3 => \N__8102\,
            lcout => \ALU.mult_AdderTree2_bigtree_543\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_13_1\,
            carryout => \ALU.regsA_result_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_7_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8204\,
            in1 => \N__8147\,
            in2 => \N__8846\,
            in3 => \N__8099\,
            lcout => \ALU.regsA_result_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_14_l_ofx_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14255\,
            in1 => \N__12600\,
            in2 => \N__8176\,
            in3 => \N__14888\,
            lcout => \ALU.regsA_result_axb_14_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_7_l_ofx_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__12966\,
            in1 => \N__14445\,
            in2 => \_gnd_net_\,
            in3 => \N__12845\,
            lcout => \ALU.addsub_axb_7_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_8_ma_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12378\,
            in1 => \N__14885\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_8_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_14_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__13519\,
            in1 => \N__14578\,
            in2 => \N__12464\,
            in3 => \N__14256\,
            lcout => \ALU.regsA_result_axb_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_14_ma_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14886\,
            lcout => \ALU.regsA_result_cry_14_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_1_l_ofx_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__12602\,
            in1 => \_gnd_net_\,
            in2 => \N__12068\,
            in3 => \N__14444\,
            lcout => \ALU.addsub_axb_1_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_15_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12601\,
            lcout => \ALU.overflow_RNOZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_0_l_ofx_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__14887\,
            in1 => \N__14443\,
            in2 => \_gnd_net_\,
            in3 => \N__13776\,
            lcout => \ALU.addsub_axb_0_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10331\,
            in2 => \N__10472\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \ALU.regsA_result_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_5_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9026\,
            in2 => \N__10388\,
            in3 => \N__8414\,
            lcout => \ALU.mult_5\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_0\,
            carryout => \ALU.regsA_result_cry_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_6_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8996\,
            in2 => \N__9845\,
            in3 => \N__8399\,
            lcout => \ALU.mult_6\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_0\,
            carryout => \ALU.regsA_result_cry_2_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_7_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8966\,
            in2 => \N__9374\,
            in3 => \N__8396\,
            lcout => \ALU.mult_7\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_1\,
            carryout => \ALU.regsA_result_cry_3_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_3_c_RNI2M12C_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8933\,
            in2 => \N__9362\,
            in3 => \N__8372\,
            lcout => \ALU.mult_AdderTree2_bigtree_932\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_1\,
            carryout => \ALU.regsA_result_cry_4_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_4_c_RNILOTIB_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8903\,
            in2 => \N__9350\,
            in3 => \N__8354\,
            lcout => \ALU.mult_AdderTree2_bigtree_933\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_0\,
            carryout => \ALU.regsA_result_cry_5_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_5_c_RNIM757B_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9260\,
            in2 => \N__9338\,
            in3 => \N__8321\,
            lcout => \ALU.mult_AdderTree2_bigtree_934\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_1\,
            carryout => \ALU.regsA_result_cry_6_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_6_c_RNIG0NPA_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9233\,
            in2 => \N__9326\,
            in3 => \N__8288\,
            lcout => \ALU.mult_AdderTree2_bigtree_935\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_0\,
            carryout => \ALU.regsA_result_cry_7_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_7_c_RNIHGF5A_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9206\,
            in2 => \N__9314\,
            in3 => \N__8258\,
            lcout => \ALU.mult_AdderTree2_bigtree_936\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \ALU.regsA_result_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_8_c_RNI026D9_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9173\,
            in2 => \N__9302\,
            in3 => \N__8231\,
            lcout => \ALU.mult_AdderTree2_bigtree_937\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_8\,
            carryout => \ALU.regsA_result_cry_9_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_9_c_RNIQQNF9_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9143\,
            in2 => \N__9290\,
            in3 => \N__8588\,
            lcout => \ALU.mult_AdderTree2_bigtree_938\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_9_0\,
            carryout => \ALU.regsA_result_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_10_c_RNIGPFR7_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9515\,
            in2 => \N__9110\,
            in3 => \N__8561\,
            lcout => \ALU.mult_AdderTree2_bigtree_939\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_10\,
            carryout => \ALU.regsA_result_cry_11_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_1_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8558\,
            in1 => \N__9086\,
            in2 => \N__8543\,
            in3 => \N__8528\,
            lcout => \ALU.regsA_result_axb_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_5_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8513\,
            in1 => \N__11265\,
            in2 => \_gnd_net_\,
            in3 => \N__8507\,
            lcout => res_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_7_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11279\,
            in1 => \N__8498\,
            in2 => \_gnd_net_\,
            in3 => \N__8489\,
            lcout => res_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_0_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__15908\,
            in1 => \N__8483\,
            in2 => \N__15674\,
            in3 => \N__8477\,
            lcout => \TXbufferZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16119\,
            ce => \N__9386\,
            sr => \_gnd_net_\
        );

    \TXbuffer_5_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__15906\,
            in1 => \N__8468\,
            in2 => \N__15675\,
            in3 => \N__8462\,
            lcout => \TXbufferZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16119\,
            ce => \N__9386\,
            sr => \_gnd_net_\
        );

    \TXbuffer_2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__8437\,
            in1 => \N__15651\,
            in2 => \N__8423\,
            in3 => \N__15909\,
            lcout => \TXbufferZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16119\,
            ce => \N__9386\,
            sr => \_gnd_net_\
        );

    \TXbuffer_6_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__8777\,
            in1 => \N__15910\,
            in2 => \N__15680\,
            in3 => \N__8768\,
            lcout => \TXbufferZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16119\,
            ce => \N__9386\,
            sr => \_gnd_net_\
        );

    \TXbuffer_7_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__15907\,
            in1 => \N__8762\,
            in2 => \N__15676\,
            in3 => \N__8753\,
            lcout => \TXbufferZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16119\,
            ce => \N__9386\,
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_11_l_ofx_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__8746\,
            in1 => \N__14458\,
            in2 => \_gnd_net_\,
            in3 => \N__10275\,
            lcout => \ALU.addsub_axb_11_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_12_l_ofx_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__14570\,
            in1 => \N__12650\,
            in2 => \N__9594\,
            in3 => \N__14862\,
            lcout => \ALU.regsA_result_axb_12_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_12_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10963\,
            lcout => \bZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16090\,
            ce => \N__14223\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_11_ma_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__9582\,
            in1 => \N__14860\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_11_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_13_ma_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9583\,
            in2 => \_gnd_net_\,
            in3 => \N__13466\,
            lcout => \ALU.regsA_result_cry_13_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_13_l_ofx_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13467\,
            in1 => \N__14560\,
            in2 => \N__9595\,
            in3 => \N__12453\,
            lcout => \ALU.regsA_result_axb_13_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_13_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12287\,
            lcout => \bZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16090\,
            ce => \N__14223\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_12_ma_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14559\,
            in2 => \_gnd_net_\,
            in3 => \N__14861\,
            lcout => \ALU.regsA_result_cry_12_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_13_l_ofx_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__12651\,
            in1 => \N__14890\,
            in2 => \N__14571\,
            in3 => \N__14266\,
            lcout => \ALU.regsA_result_axb_13_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9647\,
            in2 => \N__9656\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \ALU.regsA_result_cry_1_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNIF6113_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9866\,
            in2 => \N__9713\,
            in3 => \N__8804\,
            lcout => \ALU.mult_AdderTree2_bigtree_565\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_8\,
            carryout => \ALU.regsA_result_cry_2_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_0_c_RNIJD753_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9860\,
            in2 => \N__9704\,
            in3 => \N__8801\,
            lcout => \ALU.mult_AdderTree2_bigtree_566\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_10\,
            carryout => \ALU.regsA_result_cry_3_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_0_c_RNINKDP2_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9695\,
            in2 => \N__9854\,
            in3 => \N__8798\,
            lcout => \ALU.mult_AdderTree2_bigtree_567\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_10\,
            carryout => \ALU.regsA_result_cry_4_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_0_c_RNIRRJT2_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8795\,
            in2 => \N__9689\,
            in3 => \N__8786\,
            lcout => \ALU.mult_AdderTree2_bigtree_568\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_9\,
            carryout => \ALU.regsA_result_cry_5_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_5_0_c_RNI1R903_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9914\,
            in2 => \N__9728\,
            in3 => \N__8783\,
            lcout => \ALU.mult_AdderTree2_bigtree_569\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_9\,
            carryout => \ALU.regsA_result_cry_6_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_0_c_RNI52GK2_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9890\,
            in2 => \N__9902\,
            in3 => \N__8780\,
            lcout => \ALU.mult_AdderTree2_bigtree_570\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_8\,
            carryout => \ALU.regsA_result_cry_7_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_0_c_RNI99MO2_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9992\,
            in2 => \N__12491\,
            in3 => \N__8888\,
            lcout => \ALU.mult_AdderTree2_bigtree_571\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_7_7\,
            carryout => \ALU.regsA_result_cry_8_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_0_c_RNIDGSS2_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12476\,
            in2 => \N__12404\,
            in3 => \N__8885\,
            lcout => \ALU.mult_AdderTree2_bigtree_572\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \ALU.regsA_result_cry_9_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_0_c_RNIODOI2_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9536\,
            in2 => \N__11126\,
            in3 => \N__8882\,
            lcout => \ALU.mult_AdderTree2_bigtree_573\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_9_5\,
            carryout => \ALU.regsA_result_cry_10_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_0_c_RNIHP7H1_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9527\,
            in2 => \N__9611\,
            in3 => \N__8879\,
            lcout => \ALU.mult_AdderTree2_bigtree_574\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_10_4\,
            carryout => \ALU.regsA_result_cry_11_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_0_c_RNIL0EL1_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8837\,
            in2 => \N__9551\,
            in3 => \N__8876\,
            lcout => \ALU.mult_AdderTree2_bigtree_575\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_11_4\,
            carryout => \ALU.regsA_result_cry_12_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_0_c_RNIP7K91_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8873\,
            in2 => \N__8864\,
            in3 => \N__8852\,
            lcout => \ALU.mult_AdderTree2_bigtree_576\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_12_1\,
            carryout => \ALU.regsA_result_cry_13_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_13_0_THRU_LUT4_0_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8849\,
            lcout => \ALU.regsA_result_cry_13_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_12_ma_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10287\,
            in2 => \_gnd_net_\,
            in3 => \N__13468\,
            lcout => \ALU.regsA_result_cry_12_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_0_0_c_RNO_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12013\,
            in1 => \N__14819\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9743\,
            in2 => \N__9828\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \ALU.regsA_result_cry_0_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_3_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9680\,
            in2 => \N__9077\,
            in3 => \N__9068\,
            lcout => \ALU.mult_3\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_0_1\,
            carryout => \ALU.regsA_result_cry_1_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_1_c_RNITU8C6_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9065\,
            in2 => \N__9059\,
            in3 => \N__9047\,
            lcout => \ALU.mult_AdderTree2_bigtree_796\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_2\,
            carryout => \ALU.regsA_result_cry_2_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_2_c_RNI6FM46_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9044\,
            in2 => \N__9038\,
            in3 => \N__9017\,
            lcout => \ALU.mult_AdderTree2_bigtree_797\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_3\,
            carryout => \ALU.regsA_result_cry_3_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_3_c_RNIFV3T5_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9014\,
            in2 => \N__9008\,
            in3 => \N__8987\,
            lcout => \ALU.mult_AdderTree2_bigtree_798\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_3\,
            carryout => \ALU.regsA_result_cry_4_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_4_c_RNIOFH56_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8984\,
            in2 => \N__8978\,
            in3 => \N__8954\,
            lcout => \ALU.mult_AdderTree2_bigtree_799\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_2\,
            carryout => \ALU.regsA_result_cry_5_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_5_c_RNI3OEC6_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8951\,
            in2 => \N__8945\,
            in3 => \N__8924\,
            lcout => \ALU.mult_AdderTree2_bigtree_800\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_3\,
            carryout => \ALU.regsA_result_cry_6_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_6_c_RNIC8SK5_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8921\,
            in2 => \N__8915\,
            in3 => \N__8891\,
            lcout => \ALU.mult_AdderTree2_bigtree_801\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_2\,
            carryout => \ALU.regsA_result_cry_7_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_7_c_RNI35L05_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9278\,
            in2 => \N__9272\,
            in3 => \N__9254\,
            lcout => \ALU.mult_AdderTree2_bigtree_802\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \ALU.regsA_result_cry_8_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_8_c_RNIJBOQ4_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9251\,
            in2 => \N__9245\,
            in3 => \N__9227\,
            lcout => \ALU.mult_AdderTree2_bigtree_803\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_8_0\,
            carryout => \ALU.regsA_result_cry_9_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_9_c_RNIA92E4_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9224\,
            in2 => \N__9218\,
            in3 => \N__9194\,
            lcout => \ALU.mult_AdderTree2_bigtree_804\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_9_1\,
            carryout => \ALU.regsA_result_cry_10_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_10_c_RNIF8AD3_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9191\,
            in2 => \N__9185\,
            in3 => \N__9164\,
            lcout => \ALU.mult_AdderTree2_bigtree_805\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_10_0\,
            carryout => \ALU.regsA_result_cry_11_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_11_c_RNIOONL3_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9161\,
            in2 => \N__9155\,
            in3 => \N__9134\,
            lcout => \ALU.mult_AdderTree2_bigtree_806\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_11_2\,
            carryout => \ALU.regsA_result_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_12_c_RNI195U2_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9131\,
            in2 => \N__9125\,
            in3 => \N__9098\,
            lcout => \ALU.mult_AdderTree2_bigtree_807\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_12\,
            carryout => \ALU.regsA_result_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_3_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9503\,
            in1 => \N__9095\,
            in2 => \N__10016\,
            in3 => \N__9089\,
            lcout => \ALU.regsA_result_axb_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13550\,
            in2 => \N__13905\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \ALU.regsA_result_cry_2_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNIS7EJ4_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10445\,
            in2 => \N__9980\,
            in3 => \N__9365\,
            lcout => \ALU.mult_AdderTree2_bigtree_832\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_4\,
            carryout => \ALU.regsA_result_cry_3_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_3_c_RNIV8BJ5_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10655\,
            in2 => \N__9968\,
            in3 => \N__9353\,
            lcout => \ALU.mult_AdderTree2_bigtree_833\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_5\,
            carryout => \ALU.regsA_result_cry_4_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_4_c_RNI8POR5_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10631\,
            in2 => \N__9956\,
            in3 => \N__9341\,
            lcout => \ALU.mult_AdderTree2_bigtree_834\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_4\,
            carryout => \ALU.regsA_result_cry_5_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_5_c_RNIH9646_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10610\,
            in2 => \N__10130\,
            in3 => \N__9329\,
            lcout => \ALU.mult_AdderTree2_bigtree_835\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_5\,
            carryout => \ALU.regsA_result_cry_6_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_6_c_RNIQPJS5_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10586\,
            in2 => \N__10109\,
            in3 => \N__9317\,
            lcout => \ALU.mult_AdderTree2_bigtree_836\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_4\,
            carryout => \ALU.regsA_result_cry_7_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_7_c_RNI3A1L5_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10562\,
            in2 => \N__10076\,
            in3 => \N__9305\,
            lcout => \ALU.mult_AdderTree2_bigtree_837\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_7_4\,
            carryout => \ALU.regsA_result_cry_8_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_8_c_RNICQET5_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10538\,
            in2 => \N__10064\,
            in3 => \N__9293\,
            lcout => \ALU.mult_AdderTree2_bigtree_838\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_8_1\,
            carryout => \ALU.regsA_result_cry_9_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_9_c_RNIS0IN5_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10052\,
            in2 => \N__10523\,
            in3 => \N__9281\,
            lcout => \ALU.mult_AdderTree2_bigtree_839\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \ALU.regsA_result_cry_10_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_10_c_RNI126N4_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10043\,
            in2 => \N__10766\,
            in3 => \N__9509\,
            lcout => \ALU.mult_AdderTree2_bigtree_840\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_10_1\,
            carryout => \ALU.regsA_result_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_11_THRU_LUT4_0_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9506\,
            lcout => \ALU.regsA_result_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXstate_fast_RNIP6NA1_3_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__15662\,
            in1 => \N__15883\,
            in2 => \N__15785\,
            in3 => \N__16188\,
            lcout => \TXstate_fast_RNIP6NA1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_10_l_ofx_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__14875\,
            in1 => \N__12649\,
            in2 => \N__14157\,
            in3 => \N__10292\,
            lcout => \ALU.regsA_result_axb_10_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_3_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11264\,
            in1 => \N__9482\,
            in2 => \_gnd_net_\,
            in3 => \N__9470\,
            lcout => res_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXbuffer_3_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__15911\,
            in1 => \N__15678\,
            in2 => \N__9461\,
            in3 => \N__9446\,
            lcout => \TXbufferZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16115\,
            ce => \N__9385\,
            sr => \_gnd_net_\
        );

    \TXbuffer_1_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__9427\,
            in1 => \N__15677\,
            in2 => \N__9410\,
            in3 => \N__15913\,
            lcout => \TXbufferZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16115\,
            ce => \N__9385\,
            sr => \_gnd_net_\
        );

    \TXbuffer_4_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__15912\,
            in1 => \N__15679\,
            in2 => \N__9398\,
            in3 => \N__11153\,
            lcout => \TXbufferZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16115\,
            ce => \N__9385\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_11_l_ofx_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__9581\,
            in1 => \N__12648\,
            in2 => \N__10276\,
            in3 => \N__14841\,
            lcout => \ALU.regsA_result_axb_11_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_11_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10417\,
            lcout => \bZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16080\,
            ce => \N__14199\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_10_ma_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__10258\,
            in1 => \N__14840\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_10_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_11_l_ofx_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__10262\,
            in1 => \N__12444\,
            in2 => \N__14162\,
            in3 => \N__13533\,
            lcout => \ALU.regsA_result_axb_11_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_13_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__15189\,
            in1 => \N__10271\,
            in2 => \N__9593\,
            in3 => \N__10852\,
            lcout => \ALU.regsA_result_axb_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_12_l_ofx_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12443\,
            in1 => \N__13512\,
            in2 => \N__10286\,
            in3 => \N__9577\,
            lcout => \ALU.regsA_result_axb_12_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_10_l_ofx_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__12379\,
            in1 => \N__12442\,
            in2 => \N__13536\,
            in3 => \N__14149\,
            lcout => \ALU.regsA_result_axb_10_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_2_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11107\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16084\,
            ce => \N__15275\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_11_ma_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14148\,
            in2 => \_gnd_net_\,
            in3 => \N__13463\,
            lcout => \ALU.regsA_result_cry_11_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_2_rep1_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11108\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \a_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16084\,
            ce => \N__15275\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_2_l_ofx_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__11946\,
            in1 => \N__11746\,
            in2 => \N__13537\,
            in3 => \N__9769\,
            lcout => \ALU.regsA_result_axb_2_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_3_l_ofx_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__13464\,
            in1 => \N__11797\,
            in2 => \N__9789\,
            in3 => \N__13285\,
            lcout => \ALU.regsA_result_axb_3_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_4_l_ofx_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13286\,
            in1 => \N__11644\,
            in2 => \N__13538\,
            in3 => \N__9773\,
            lcout => \ALU.regsA_result_axb_4_l_ofx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_5_l_ofx_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__13465\,
            in1 => \N__11645\,
            in2 => \N__9790\,
            in3 => \N__15024\,
            lcout => \ALU.regsA_result_axb_5_l_ofx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_1_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__13726\,
            in1 => \N__13439\,
            in2 => \N__9671\,
            in3 => \N__11945\,
            lcout => \ALU.mult_AdderTree2_bigtree_564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_fast_2_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11105\,
            lcout => \a_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16091\,
            ce => \N__15249\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__13727\,
            in1 => \N__13440\,
            in2 => \N__11993\,
            in3 => \N__9667\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_3_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10420\,
            lcout => \aZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16091\,
            ce => \N__15249\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_1_0_c_RNO_0_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13642\,
            in2 => \_gnd_net_\,
            in3 => \N__13435\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_2_ma_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13436\,
            in1 => \N__11944\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_2_ma_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_3_ma_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11749\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13437\,
            lcout => \ALU.regsA_result_cry_3_ma_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_4_ma_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13438\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13287\,
            lcout => \ALU.regsA_result_cry_4_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNIUA504_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__13906\,
            in1 => \N__13869\,
            in2 => \_gnd_net_\,
            in3 => \N__13670\,
            lcout => \ALU.mult_AdderTree2_bigtree_831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_0_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14503\,
            lcout => \bZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16096\,
            ce => \N__11396\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__9830\,
            in1 => \N__9791\,
            in2 => \_gnd_net_\,
            in3 => \N__13669\,
            lcout => \ALU.regsA_result_cry_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_4_ma_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14998\,
            in2 => \_gnd_net_\,
            in3 => \N__14820\,
            lcout => \ALU.regsA_result_cry_4_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_5_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12282\,
            lcout => \bZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16096\,
            ce => \N__11396\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_6_ma_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14999\,
            lcout => \ALU.regsA_result_cry_6_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_6_l_ofx_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__12806\,
            in1 => \N__14832\,
            in2 => \N__13068\,
            in3 => \N__12607\,
            lcout => \ALU.regsA_result_axb_6_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_6_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14307\,
            lcout => \bZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16102\,
            ce => \N__11387\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_5_ma_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14831\,
            lcout => \ALU.regsA_result_cry_5_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_6_l_ofx_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15001\,
            in1 => \N__15188\,
            in2 => \N__13067\,
            in3 => \N__10833\,
            lcout => \ALU.regsA_result_axb_6_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_6_l_ofx_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12454\,
            in1 => \N__13039\,
            in2 => \N__13521\,
            in3 => \N__15000\,
            lcout => \ALU.regsA_result_axb_6_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_7_ma_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13488\,
            in2 => \N__13069\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_7_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_7_l_ofx_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12455\,
            in1 => \N__13043\,
            in2 => \N__13522\,
            in3 => \N__12805\,
            lcout => \ALU.regsA_result_axb_7_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_7_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12115\,
            lcout => \bZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16104\,
            ce => \N__11395\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_6_ma_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14847\,
            lcout => \ALU.regsA_result_cry_6_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_ma_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12803\,
            in2 => \_gnd_net_\,
            in3 => \N__15180\,
            lcout => \ALU.regsA_result_cry_8_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_7_l_ofx_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15181\,
            in1 => \N__13054\,
            in2 => \N__10847\,
            in3 => \N__12831\,
            lcout => \ALU.regsA_result_axb_7_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_8_ma_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12802\,
            in2 => \_gnd_net_\,
            in3 => \N__13495\,
            lcout => \ALU.regsA_result_cry_8_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_8_l_ofx_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15182\,
            in1 => \N__12832\,
            in2 => \N__10848\,
            in3 => \N__13171\,
            lcout => \ALU.regsA_result_axb_8_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_7_l_ofx_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13055\,
            in1 => \N__13867\,
            in2 => \N__12968\,
            in3 => \N__12804\,
            lcout => \ALU.regsA_result_axb_7_l_ofx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10370\,
            in2 => \N__10700\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \ALU.regsA_result_cry_1_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNI5R443_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10358\,
            in2 => \N__10724\,
            in3 => \N__9983\,
            lcout => \ALU.mult_AdderTree2_bigtree_600\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_7\,
            carryout => \ALU.regsA_result_cry_2_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_0_c_RNI92BO2_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12143\,
            in2 => \N__10346\,
            in3 => \N__9971\,
            lcout => \ALU.mult_AdderTree2_bigtree_601\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_9\,
            carryout => \ALU.regsA_result_cry_3_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_0_c_RNI0ARQ2_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10889\,
            in2 => \N__10682\,
            in3 => \N__9959\,
            lcout => \ALU.mult_AdderTree2_bigtree_602\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_9\,
            carryout => \ALU.regsA_result_cry_4_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_0_c_RNI4H1V2_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10883\,
            in2 => \N__10910\,
            in3 => \N__9947\,
            lcout => \ALU.mult_AdderTree2_bigtree_603\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_8\,
            carryout => \ALU.regsA_result_cry_5_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_0_c_RNI8O733_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10877\,
            in2 => \N__10142\,
            in3 => \N__10121\,
            lcout => \ALU.mult_AdderTree2_bigtree_604\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_8\,
            carryout => \ALU.regsA_result_cry_6_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_0_c_RNICVDN2_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10715\,
            in2 => \N__10118\,
            in3 => \N__10100\,
            lcout => \ALU.mult_AdderTree2_bigtree_605\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_7\,
            carryout => \ALU.regsA_result_cry_7_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_0_c_RNIG6KR2_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10097\,
            in2 => \N__10088\,
            in3 => \N__10067\,
            lcout => \ALU.mult_AdderTree2_bigtree_606\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_7_6\,
            carryout => \ALU.regsA_result_cry_8_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_8_0_c_RNIKDQV2_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10736\,
            in2 => \N__10775\,
            in3 => \N__10055\,
            lcout => \ALU.mult_AdderTree2_bigtree_607\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \ALU.regsA_result_cry_9_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_0_c_RNIVAML2_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10217\,
            in2 => \N__10001\,
            in3 => \N__10046\,
            lcout => \ALU.mult_AdderTree2_bigtree_608\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_9_4\,
            carryout => \ALU.regsA_result_cry_10_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_0_c_RNIONSH1_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10298\,
            in2 => \N__10226\,
            in3 => \N__10037\,
            lcout => \ALU.mult_AdderTree2_bigtree_609\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_10_3\,
            carryout => \ALU.regsA_result_cry_11_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_6_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10709\,
            in1 => \N__10745\,
            in2 => \N__10034\,
            in3 => \N__10019\,
            lcout => \ALU.regsA_result_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_10_l_ofx_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__12355\,
            in1 => \N__10828\,
            in2 => \N__15205\,
            in3 => \N__14127\,
            lcout => \ALU.regsA_result_axb_10_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_11_ma_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__14128\,
            in1 => \_gnd_net_\,
            in2 => \N__15206\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_11_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_11_l_ofx_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__15199\,
            in1 => \N__10829\,
            in2 => \N__10291\,
            in3 => \N__14129\,
            lcout => \ALU.regsA_result_axb_11_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_10_ma_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12354\,
            lcout => \ALU.regsA_result_cry_10_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_1_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10196\,
            in1 => \N__15424\,
            in2 => \_gnd_net_\,
            in3 => \N__10211\,
            lcout => \FTDI.TXshiftZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15425\,
            in1 => \N__10148\,
            in2 => \_gnd_net_\,
            in3 => \N__10205\,
            lcout => \FTDI.TXshiftZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_6_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__15429\,
            in2 => \_gnd_net_\,
            in3 => \N__10190\,
            lcout => \FTDI.TXshiftZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_4_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15427\,
            in1 => \N__10304\,
            in2 => \_gnd_net_\,
            in3 => \N__10181\,
            lcout => \FTDI.TXshiftZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_0_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10175\,
            in1 => \N__15423\,
            in2 => \_gnd_net_\,
            in3 => \N__10169\,
            lcout => \FTDI.TXshiftZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_3_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10160\,
            in1 => \N__10154\,
            in2 => \_gnd_net_\,
            in3 => \N__15426\,
            lcout => \FTDI.TXshiftZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_5_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15428\,
            in1 => \N__10319\,
            in2 => \_gnd_net_\,
            in3 => \N__10313\,
            lcout => \FTDI.TXshiftZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_1C_net\,
            ce => \N__12713\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_2_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10418\,
            lcout => \RXbuffer_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_2C_net\,
            ce => \N__10993\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_4_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12271\,
            lcout => \RXbuffer_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_2C_net\,
            ce => \N__10993\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_3_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10942\,
            lcout => \RXbuffer_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_2C_net\,
            ce => \N__10993\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_7_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11024\,
            lcout => \RXbuffer_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_2C_net\,
            ce => \N__10993\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_5_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14296\,
            lcout => \RXbuffer_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_5C_net\,
            ce => \N__10997\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_0_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11320\,
            lcout => \RXbuffer_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_5C_net\,
            ce => \N__10997\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_6_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12103\,
            lcout => \RXbuffer_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_5C_net\,
            ce => \N__10997\,
            sr => \_gnd_net_\
        );

    \FTDI.RXbuffer_1_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11084\,
            lcout => \RXbuffer_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXbuffer_5C_net\,
            ce => \N__10997\,
            sr => \_gnd_net_\
        );

    \b_1_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11314\,
            lcout => \bZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16081\,
            ce => \N__11374\,
            sr => \_gnd_net_\
        );

    \b_2_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11094\,
            lcout => \bZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16081\,
            ce => \N__11374\,
            sr => \_gnd_net_\
        );

    \b_3_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10419\,
            lcout => \bZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16081\,
            ce => \N__11374\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_1_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__13671\,
            in1 => \N__15159\,
            in2 => \N__11948\,
            in3 => \N__10505\,
            lcout => \ALU.mult_AdderTree2_bigtree_599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_fast_4_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10943\,
            lcout => \a_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16085\,
            ce => \N__15264\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__13674\,
            in1 => \N__10491\,
            in2 => \N__11947\,
            in3 => \N__15161\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_2_l_ofx_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__15160\,
            in1 => \N__11904\,
            in2 => \N__10503\,
            in3 => \N__11747\,
            lcout => \ALU.regsA_result_axb_2_l_ofx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_3_l_ofx_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__11748\,
            in1 => \N__10495\,
            in2 => \N__15190\,
            in3 => \N__13252\,
            lcout => \ALU.regsA_result_axb_3_l_ofx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_3_m1_forloop_1_1_regsA_result_cry_0_c_RNO_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__10471\,
            in1 => \_gnd_net_\,
            in2 => \N__10504\,
            in3 => \N__13672\,
            lcout => \ALU.regsA_result_cry_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_RNO_1_4_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__13673\,
            in1 => \N__10499\,
            in2 => \_gnd_net_\,
            in3 => \N__10470\,
            lcout => \ALU.mult_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_5_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12286\,
            lcout => \aZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16085\,
            ce => \N__15264\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_1_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__12940\,
            in1 => \N__13643\,
            in2 => \N__13873\,
            in3 => \N__11967\,
            lcout => \ALU.mult_AdderTree2_bigtree_634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_6_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \aZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16092\,
            ce => \N__15285\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__12948\,
            in1 => \N__13644\,
            in2 => \N__11994\,
            in3 => \N__13828\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_2_l_ofx_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__11968\,
            in1 => \N__12941\,
            in2 => \N__13864\,
            in3 => \N__11781\,
            lcout => \ALU.regsA_result_axb_2_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_3_l_ofx_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__11782\,
            in1 => \N__13297\,
            in2 => \N__12962\,
            in3 => \N__13832\,
            lcout => \ALU.regsA_result_axb_3_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_4_l_ofx_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__13298\,
            in1 => \N__12945\,
            in2 => \N__13865\,
            in3 => \N__11646\,
            lcout => \ALU.regsA_result_axb_4_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_5_l_ofx_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__12946\,
            in1 => \N__13836\,
            in2 => \N__11662\,
            in3 => \N__14987\,
            lcout => \ALU.regsA_result_axb_5_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_6_l_ofx_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14988\,
            in1 => \N__12947\,
            in2 => \N__13866\,
            in3 => \N__13044\,
            lcout => \ALU.regsA_result_axb_6_l_ofx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10691\,
            in2 => \N__10673\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \ALU.regsA_result_cry_1_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNIVOCL2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11840\,
            in2 => \N__10664\,
            in3 => \N__10643\,
            lcout => \ALU.mult_AdderTree2_bigtree_635\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_1_9\,
            carryout => \ALU.regsA_result_cry_2_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_0_c_RNI30JP2_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11678\,
            in2 => \N__10640\,
            in3 => \N__10619\,
            lcout => \ALU.mult_AdderTree2_bigtree_636\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_2_11\,
            carryout => \ALU.regsA_result_cry_3_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_0_c_RNI77PT2_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10616\,
            in2 => \N__11672\,
            in3 => \N__10598\,
            lcout => \ALU.mult_AdderTree2_bigtree_637\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_3_11\,
            carryout => \ALU.regsA_result_cry_4_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_0_c_RNIBEV13_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11522\,
            in2 => \N__10595\,
            in3 => \N__10574\,
            lcout => \ALU.mult_AdderTree2_bigtree_638\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_4_10\,
            carryout => \ALU.regsA_result_cry_5_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_0_c_RNIFL5M2_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12659\,
            in2 => \N__10571\,
            in3 => \N__10550\,
            lcout => \ALU.mult_AdderTree2_bigtree_639\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_5_10\,
            carryout => \ALU.regsA_result_cry_6_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_0_c_RNIJSBQ2_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12974\,
            in2 => \N__10547\,
            in3 => \N__10526\,
            lcout => \ALU.mult_AdderTree2_bigtree_640\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_6_9\,
            carryout => \ALU.regsA_result_cry_7_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_0_c_RNIN3IU2_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12389\,
            in2 => \N__12761\,
            in3 => \N__10508\,
            lcout => \ALU.mult_AdderTree2_bigtree_641\,
            ltout => OPEN,
            carryin => \ALU.regsA_result_cry_7_8\,
            carryout => \ALU.regsA_result_cry_8_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_0_c_RNIRAO23_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13097\,
            in2 => \N__12296\,
            in3 => \N__10751\,
            lcout => \ALU.mult_AdderTree2_bigtree_642\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \ALU.regsA_result_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.regsA_result_cry_9_THRU_LUT4_0_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10748\,
            lcout => \ALU.regsA_result_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_9_ma_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13153\,
            in2 => \_gnd_net_\,
            in3 => \N__15134\,
            lcout => \ALU.regsA_result_cry_9_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_2_ma_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11970\,
            lcout => \ALU.regsA_result_cry_2_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_7_ma_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13045\,
            in1 => \N__15135\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_7_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.overflow_RNO_12_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__12371\,
            in1 => \N__13868\,
            in2 => \N__14153\,
            in3 => \N__12939\,
            lcout => \ALU.regsA_result_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_1_0_c_RNO_0_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13676\,
            in1 => \N__15132\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_1_0_c_RNO_0_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13675\,
            in2 => \_gnd_net_\,
            in3 => \N__12938\,
            lcout => \ALU.regsA_result_cry_1_0_c_RNO_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_4_l_ofx_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13346\,
            in1 => \N__11651\,
            in2 => \N__15179\,
            in3 => \N__10822\,
            lcout => \ALU.regsA_result_axb_4_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_4_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10956\,
            lcout => \aZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16105\,
            ce => \N__15296\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_5_l_ofx_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__10823\,
            in2 => \N__11663\,
            in3 => \N__15017\,
            lcout => \ALU.regsA_result_axb_5_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_4_l_ofx_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11653\,
            in1 => \_gnd_net_\,
            in2 => \N__10843\,
            in3 => \N__14426\,
            lcout => \ALU.addsub_axb_4_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_4_ma_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13296\,
            in1 => \N__15136\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_4_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_5_ma_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__15137\,
            in1 => \N__11652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_5_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_6_ma_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15138\,
            lcout => \ALU.regsA_result_cry_6_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_9_l_ofx_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__14130\,
            in1 => \N__14874\,
            in2 => \N__12652\,
            in3 => \N__12353\,
            lcout => \ALU.regsA_result_axb_9_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_9_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11331\,
            lcout => \bZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16107\,
            ce => \N__14224\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_axb_9_l_ofx_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__15195\,
            in1 => \N__12352\,
            in2 => \N__13184\,
            in3 => \N__10827\,
            lcout => \ALU.regsA_result_axb_9_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_10_ma_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12351\,
            in1 => \N__13534\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_10_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_10_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11099\,
            lcout => \bZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16107\,
            ce => \N__14224\,
            sr => \_gnd_net_\
        );

    \FTDI.TXshift_7_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15422\,
            in2 => \_gnd_net_\,
            in3 => \N__11039\,
            lcout => \FTDI.TXshiftZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.TXshift_7C_net\,
            ce => \N__12712\,
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNIV5TH_0_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11510\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13951\,
            lcout => \FTDI.N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNO_0_3_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110001"
        )
    port map (
            in0 => \N__11451\,
            in1 => \N__11023\,
            in2 => \N__11495\,
            in3 => \N__11417\,
            lcout => OPEN,
            ltout => \FTDI.m13_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_3_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101010000"
        )
    port map (
            in0 => \N__11511\,
            in1 => \N__13956\,
            in2 => \N__11000\,
            in3 => \N__11490\,
            lcout => \FTDI.RXstateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXstate_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_1_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__11489\,
            in1 => \N__11418\,
            in2 => \N__13958\,
            in3 => \N__11513\,
            lcout => \FTDI.RXstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXstate_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_RNI29TH_2_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13952\,
            in2 => \_gnd_net_\,
            in3 => \N__11488\,
            lcout => \FTDI.N_201_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNI67DS1_0_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11449\,
            in1 => \N__11415\,
            in2 => \N__11494\,
            in3 => \N__11509\,
            lcout => \FTDI.gap8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_RNO_0_0_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111110"
        )
    port map (
            in0 => \N__11416\,
            in1 => \N__11450\,
            in2 => \N__13957\,
            in3 => \N__11484\,
            lcout => OPEN,
            ltout => \FTDI.N_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_0_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110001000"
        )
    port map (
            in0 => \N__11491\,
            in1 => \N__13950\,
            in2 => \N__11516\,
            in3 => \N__11512\,
            lcout => \FTDI.RXstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXstate_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXstate_2_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__11420\,
            in1 => \N__11431\,
            in2 => \N__11456\,
            in3 => \N__11493\,
            lcout => \FTDI.RXstateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXstate_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXready_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11492\,
            in1 => \N__11452\,
            in2 => \N__11432\,
            in3 => \N__11419\,
            lcout => \RXready\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.RXstate_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXready_RNIICV7_1_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__15605\,
            in1 => \N__15881\,
            in2 => \N__15783\,
            in3 => \N__15498\,
            lcout => \RXready_RNIICV7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXready_RNIICV7_0_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15584\,
            in1 => \N__15880\,
            in2 => \N__15782\,
            in3 => \N__15499\,
            lcout => \RXready_RNIICV7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \op_1_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__15500\,
            in1 => \N__11321\,
            in2 => \N__15962\,
            in3 => \N__11203\,
            lcout => \opZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.res_4_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11202\,
            in1 => \N__11174\,
            in2 => \_gnd_net_\,
            in3 => \N__11159\,
            lcout => res_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_7_regsA_result_cry_2_ma_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14603\,
            in2 => \_gnd_net_\,
            in3 => \N__11940\,
            lcout => \ALU.regsA_result_cry_2_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_13_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12281\,
            lcout => \aZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16079\,
            ce => \N__12213\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_1_ma_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11729\,
            in2 => \_gnd_net_\,
            in3 => \N__14740\,
            lcout => \ALU.regsA_result_cry_1_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_3_regsA_result_cry_3_ma_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15099\,
            lcout => \ALU.regsA_result_cry_3_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_2_ma_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13264\,
            in2 => \_gnd_net_\,
            in3 => \N__14741\,
            lcout => \ALU.regsA_result_cry_2_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_7_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12114\,
            lcout => \aZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16082\,
            ce => \N__15274\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_2_ma_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__11969\,
            in1 => \N__12926\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_2_ma_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_3_ma_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12927\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11783\,
            lcout => \ALU.regsA_result_cry_3_ma_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_4_ma_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13299\,
            in1 => \N__12928\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_4_ma_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_5_ma_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11650\,
            lcout => \ALU.regsA_result_cry_5_ma_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_6_ma_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__15005\,
            in1 => \N__12930\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_6_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_axb_8_l_ofx_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13152\,
            in1 => \N__14753\,
            in2 => \N__12653\,
            in3 => \N__12370\,
            lcout => \ALU.regsA_result_axb_8_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_8_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14516\,
            lcout => \bZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16087\,
            ce => \N__14219\,
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_7_ma_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13148\,
            in1 => \N__14752\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_7_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_8_l_ofx_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13515\,
            in1 => \N__12456\,
            in2 => \N__12857\,
            in3 => \N__13149\,
            lcout => \ALU.regsA_result_axb_8_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_cry_9_ma_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__13151\,
            in1 => \N__13514\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_9_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_2_regsA_result_axb_9_l_ofx_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13155\,
            in1 => \N__12457\,
            in2 => \N__13535\,
            in3 => \N__12368\,
            lcout => \ALU.regsA_result_axb_9_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_8_l_ofx_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13150\,
            in1 => \N__12934\,
            in2 => \N__13878\,
            in3 => \N__12856\,
            lcout => \ALU.regsA_result_axb_8_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_axb_9_l_ofx_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13156\,
            in1 => \N__12369\,
            in2 => \N__12961\,
            in3 => \N__13863\,
            lcout => \ALU.regsA_result_axb_9_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_6_l_ofx_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13080\,
            in1 => \_gnd_net_\,
            in2 => \N__13880\,
            in3 => \N__14372\,
            lcout => \ALU.addsub_axb_6_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_2_m1_forloop_1_2_regsA_result_cry_2_c_RNO_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__13913\,
            in1 => \N__13874\,
            in2 => \_gnd_net_\,
            in3 => \N__13748\,
            lcout => \ALU.regsA_result_cry_2_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_3_l_ofx_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14371\,
            in1 => \N__13520\,
            in2 => \_gnd_net_\,
            in3 => \N__13338\,
            lcout => \ALU.addsub_axb_3_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_9_ma_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13154\,
            in2 => \_gnd_net_\,
            in3 => \N__12951\,
            lcout => \ALU.regsA_result_cry_9_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_7_ma_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12949\,
            in2 => \_gnd_net_\,
            in3 => \N__13079\,
            lcout => \ALU.regsA_result_cry_7_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_4_regsA_result_cry_8_ma_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12950\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12830\,
            lcout => \ALU.regsA_result_cry_8_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.baudAcc_RNID8HD2_2_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__16186\,
            in1 => \N__12752\,
            in2 => \N__15435\,
            in3 => \N__12682\,
            lcout => \FTDI.un1_TXstate_0_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TXstart_esr_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__15849\,
            in1 => \N__15768\,
            in2 => \N__15650\,
            in3 => \N__16185\,
            lcout => \TXstartZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16098\,
            ce => \N__12671\,
            sr => \N__15961\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_9_ma_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14112\,
            in1 => \N__14821\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.regsA_result_cry_9_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_2_c_inv_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__14063\,
            in1 => \N__15454\,
            in2 => \_gnd_net_\,
            in3 => \N__14027\,
            lcout => \FTDI.un3_TX_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_1_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__13981\,
            in1 => \N__13969\,
            in2 => \_gnd_net_\,
            in3 => \N__13993\,
            lcout => \FTDI.gapZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_0_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13968\,
            in2 => \_gnd_net_\,
            in3 => \N__13992\,
            lcout => \FTDI.gapZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.gap_2_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__13994\,
            in1 => \N__13982\,
            in2 => \N__13973\,
            in3 => \_gnd_net_\,
            lcout => \FTDI.gapZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVFTDI.gap_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXready_RNIICV7_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15606\,
            in1 => \N__15882\,
            in2 => \N__15784\,
            in3 => \N__15501\,
            lcout => \RXready_RNIICV7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_10_2_0__m7_x1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101010"
        )
    port map (
            in0 => \N__15573\,
            in1 => \N__15853\,
            in2 => \N__15760\,
            in3 => \N__15502\,
            lcout => m7_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.RXready_RNIICV7_2_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15504\,
            in1 => \N__15735\,
            in2 => \N__15879\,
            in3 => \N__15572\,
            lcout => \RXready_RNIICV7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_10_2_0__m7_x0_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010101010"
        )
    port map (
            in0 => \N__15574\,
            in1 => \N__15854\,
            in2 => \N__15761\,
            in3 => \N__15503\,
            lcout => OPEN,
            ltout => \m7_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_1_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15305\,
            in2 => \N__15299\,
            in3 => \N__16196\,
            lcout => \testStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \a_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14510\,
            lcout => \aZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16093\,
            ce => \N__15273\,
            sr => \_gnd_net_\
        );

    \testState_RNIJBO_1_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15601\,
            in2 => \_gnd_net_\,
            in3 => \N__15872\,
            lcout => OPEN,
            ltout => \testState30_testState30_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_2_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101011101010"
        )
    port map (
            in0 => \N__15731\,
            in1 => \N__15518\,
            in2 => \N__15209\,
            in3 => \N__16195\,
            lcout => \testStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_5_l_ofx_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__15191\,
            in1 => \N__14368\,
            in2 => \_gnd_net_\,
            in3 => \N__15036\,
            lcout => \ALU.addsub_axb_5_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_AdderTree2_forloop2_1_m1_forloop_1_1_regsA_result_cry_13_ma_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14243\,
            in2 => \_gnd_net_\,
            in3 => \N__14754\,
            lcout => \ALU.regsA_result_cry_13_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_axb_13_l_ofx_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__14622\,
            in1 => \N__14579\,
            in2 => \_gnd_net_\,
            in3 => \N__14369\,
            lcout => \ALU.addsub_axb_13_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \op_0_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__15954\,
            in1 => \N__15517\,
            in2 => \N__14515\,
            in3 => \N__14370\,
            lcout => \opZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_14_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14317\,
            lcout => \bZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16103\,
            ce => \N__14215\,
            sr => \_gnd_net_\
        );

    \testState_10_2_0__i3_mux_i_x0_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110110101010"
        )
    port map (
            in0 => \N__15828\,
            in1 => \N__15734\,
            in2 => \N__15646\,
            in3 => \N__15516\,
            lcout => OPEN,
            ltout => \i3_mux_i_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_0_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15461\,
            in2 => \N__16199\,
            in3 => \N__16187\,
            lcout => \testStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_RNIUI41_2_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15732\,
            in1 => \N__15612\,
            in2 => \_gnd_net_\,
            in3 => \N__15826\,
            lcout => \testState27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \testState_10_2_0__i3_mux_i_x1_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100010"
        )
    port map (
            in0 => \N__15827\,
            in1 => \N__15733\,
            in2 => \N__15645\,
            in3 => \N__15515\,
            lcout => i3_mux_i_x1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_2_c_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15455\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \FTDI.un3_TX_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_3_c_inv_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15443\,
            in2 => \_gnd_net_\,
            in3 => \N__15437\,
            lcout => \FTDI.un3_TX_axb_3\,
            ltout => OPEN,
            carryin => \FTDI.un3_TX_cry_2\,
            carryout => \FTDI.un3_TX_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__15436\,
            in1 => \N__15341\,
            in2 => \_gnd_net_\,
            in3 => \N__15329\,
            lcout => \FTDI_TX_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
