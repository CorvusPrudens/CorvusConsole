// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Aug 15 2020 12:51:41

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    TX,
    GPIO11,
    CLK,
    RX,
    GPIO9,
    GPIO3);

    output TX;
    output GPIO11;
    input CLK;
    input RX;
    output GPIO9;
    output GPIO3;

    wire N__57007;
    wire N__57006;
    wire N__57005;
    wire N__56996;
    wire N__56995;
    wire N__56994;
    wire N__56987;
    wire N__56986;
    wire N__56985;
    wire N__56978;
    wire N__56977;
    wire N__56976;
    wire N__56969;
    wire N__56968;
    wire N__56967;
    wire N__56950;
    wire N__56949;
    wire N__56948;
    wire N__56947;
    wire N__56946;
    wire N__56945;
    wire N__56942;
    wire N__56937;
    wire N__56932;
    wire N__56929;
    wire N__56920;
    wire N__56917;
    wire N__56914;
    wire N__56911;
    wire N__56908;
    wire N__56905;
    wire N__56904;
    wire N__56901;
    wire N__56900;
    wire N__56897;
    wire N__56896;
    wire N__56895;
    wire N__56894;
    wire N__56891;
    wire N__56888;
    wire N__56885;
    wire N__56882;
    wire N__56877;
    wire N__56866;
    wire N__56865;
    wire N__56864;
    wire N__56863;
    wire N__56862;
    wire N__56861;
    wire N__56858;
    wire N__56851;
    wire N__56846;
    wire N__56839;
    wire N__56838;
    wire N__56837;
    wire N__56836;
    wire N__56835;
    wire N__56834;
    wire N__56833;
    wire N__56832;
    wire N__56831;
    wire N__56826;
    wire N__56817;
    wire N__56816;
    wire N__56811;
    wire N__56810;
    wire N__56807;
    wire N__56804;
    wire N__56801;
    wire N__56800;
    wire N__56799;
    wire N__56798;
    wire N__56797;
    wire N__56796;
    wire N__56795;
    wire N__56792;
    wire N__56789;
    wire N__56786;
    wire N__56781;
    wire N__56778;
    wire N__56773;
    wire N__56768;
    wire N__56763;
    wire N__56760;
    wire N__56743;
    wire N__56742;
    wire N__56741;
    wire N__56740;
    wire N__56739;
    wire N__56738;
    wire N__56737;
    wire N__56732;
    wire N__56727;
    wire N__56720;
    wire N__56713;
    wire N__56710;
    wire N__56707;
    wire N__56704;
    wire N__56703;
    wire N__56702;
    wire N__56701;
    wire N__56696;
    wire N__56695;
    wire N__56692;
    wire N__56689;
    wire N__56686;
    wire N__56681;
    wire N__56674;
    wire N__56673;
    wire N__56670;
    wire N__56669;
    wire N__56666;
    wire N__56661;
    wire N__56656;
    wire N__56655;
    wire N__56652;
    wire N__56649;
    wire N__56644;
    wire N__56641;
    wire N__56640;
    wire N__56635;
    wire N__56632;
    wire N__56629;
    wire N__56626;
    wire N__56623;
    wire N__56620;
    wire N__56617;
    wire N__56614;
    wire N__56611;
    wire N__56608;
    wire N__56605;
    wire N__56602;
    wire N__56599;
    wire N__56596;
    wire N__56593;
    wire N__56590;
    wire N__56587;
    wire N__56586;
    wire N__56583;
    wire N__56580;
    wire N__56579;
    wire N__56578;
    wire N__56573;
    wire N__56570;
    wire N__56567;
    wire N__56564;
    wire N__56561;
    wire N__56558;
    wire N__56555;
    wire N__56550;
    wire N__56545;
    wire N__56542;
    wire N__56539;
    wire N__56536;
    wire N__56533;
    wire N__56530;
    wire N__56527;
    wire N__56524;
    wire N__56521;
    wire N__56518;
    wire N__56515;
    wire N__56512;
    wire N__56509;
    wire N__56508;
    wire N__56507;
    wire N__56506;
    wire N__56505;
    wire N__56504;
    wire N__56501;
    wire N__56498;
    wire N__56495;
    wire N__56492;
    wire N__56489;
    wire N__56488;
    wire N__56485;
    wire N__56482;
    wire N__56481;
    wire N__56478;
    wire N__56477;
    wire N__56476;
    wire N__56475;
    wire N__56472;
    wire N__56469;
    wire N__56466;
    wire N__56463;
    wire N__56460;
    wire N__56457;
    wire N__56454;
    wire N__56451;
    wire N__56448;
    wire N__56445;
    wire N__56442;
    wire N__56437;
    wire N__56434;
    wire N__56431;
    wire N__56426;
    wire N__56423;
    wire N__56420;
    wire N__56417;
    wire N__56414;
    wire N__56413;
    wire N__56410;
    wire N__56399;
    wire N__56398;
    wire N__56397;
    wire N__56394;
    wire N__56389;
    wire N__56386;
    wire N__56381;
    wire N__56378;
    wire N__56375;
    wire N__56372;
    wire N__56369;
    wire N__56366;
    wire N__56363;
    wire N__56360;
    wire N__56357;
    wire N__56354;
    wire N__56351;
    wire N__56348;
    wire N__56343;
    wire N__56334;
    wire N__56331;
    wire N__56326;
    wire N__56323;
    wire N__56322;
    wire N__56319;
    wire N__56316;
    wire N__56311;
    wire N__56308;
    wire N__56305;
    wire N__56304;
    wire N__56303;
    wire N__56302;
    wire N__56301;
    wire N__56300;
    wire N__56299;
    wire N__56298;
    wire N__56297;
    wire N__56296;
    wire N__56295;
    wire N__56294;
    wire N__56293;
    wire N__56292;
    wire N__56291;
    wire N__56290;
    wire N__56289;
    wire N__56288;
    wire N__56287;
    wire N__56286;
    wire N__56285;
    wire N__56284;
    wire N__56283;
    wire N__56282;
    wire N__56281;
    wire N__56280;
    wire N__56279;
    wire N__56278;
    wire N__56277;
    wire N__56276;
    wire N__56275;
    wire N__56274;
    wire N__56273;
    wire N__56272;
    wire N__56271;
    wire N__56270;
    wire N__56269;
    wire N__56268;
    wire N__56267;
    wire N__56266;
    wire N__56265;
    wire N__56264;
    wire N__56263;
    wire N__56262;
    wire N__56261;
    wire N__56260;
    wire N__56259;
    wire N__56258;
    wire N__56257;
    wire N__56256;
    wire N__56255;
    wire N__56254;
    wire N__56253;
    wire N__56252;
    wire N__56251;
    wire N__56250;
    wire N__56249;
    wire N__56248;
    wire N__56247;
    wire N__56246;
    wire N__56245;
    wire N__56244;
    wire N__56243;
    wire N__56242;
    wire N__56241;
    wire N__56240;
    wire N__56239;
    wire N__56238;
    wire N__56237;
    wire N__56236;
    wire N__56235;
    wire N__56234;
    wire N__56233;
    wire N__56232;
    wire N__56231;
    wire N__56230;
    wire N__56229;
    wire N__56228;
    wire N__56227;
    wire N__56226;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56058;
    wire N__56057;
    wire N__56056;
    wire N__56055;
    wire N__56054;
    wire N__56053;
    wire N__56052;
    wire N__56051;
    wire N__56050;
    wire N__56049;
    wire N__56048;
    wire N__56047;
    wire N__56046;
    wire N__56045;
    wire N__56044;
    wire N__56043;
    wire N__56042;
    wire N__56041;
    wire N__56040;
    wire N__56039;
    wire N__56038;
    wire N__56037;
    wire N__56036;
    wire N__55987;
    wire N__55984;
    wire N__55981;
    wire N__55978;
    wire N__55975;
    wire N__55972;
    wire N__55969;
    wire N__55968;
    wire N__55965;
    wire N__55962;
    wire N__55961;
    wire N__55960;
    wire N__55959;
    wire N__55958;
    wire N__55957;
    wire N__55956;
    wire N__55955;
    wire N__55952;
    wire N__55951;
    wire N__55950;
    wire N__55947;
    wire N__55946;
    wire N__55943;
    wire N__55942;
    wire N__55941;
    wire N__55940;
    wire N__55939;
    wire N__55934;
    wire N__55933;
    wire N__55932;
    wire N__55931;
    wire N__55930;
    wire N__55929;
    wire N__55928;
    wire N__55927;
    wire N__55924;
    wire N__55921;
    wire N__55920;
    wire N__55919;
    wire N__55916;
    wire N__55913;
    wire N__55910;
    wire N__55905;
    wire N__55904;
    wire N__55903;
    wire N__55902;
    wire N__55901;
    wire N__55900;
    wire N__55899;
    wire N__55896;
    wire N__55893;
    wire N__55888;
    wire N__55885;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55871;
    wire N__55862;
    wire N__55861;
    wire N__55858;
    wire N__55853;
    wire N__55848;
    wire N__55847;
    wire N__55842;
    wire N__55841;
    wire N__55840;
    wire N__55839;
    wire N__55834;
    wire N__55831;
    wire N__55826;
    wire N__55819;
    wire N__55818;
    wire N__55817;
    wire N__55814;
    wire N__55809;
    wire N__55808;
    wire N__55807;
    wire N__55806;
    wire N__55805;
    wire N__55802;
    wire N__55801;
    wire N__55800;
    wire N__55799;
    wire N__55798;
    wire N__55787;
    wire N__55784;
    wire N__55777;
    wire N__55776;
    wire N__55773;
    wire N__55772;
    wire N__55769;
    wire N__55766;
    wire N__55763;
    wire N__55760;
    wire N__55759;
    wire N__55754;
    wire N__55749;
    wire N__55744;
    wire N__55741;
    wire N__55738;
    wire N__55737;
    wire N__55736;
    wire N__55731;
    wire N__55730;
    wire N__55729;
    wire N__55724;
    wire N__55723;
    wire N__55722;
    wire N__55719;
    wire N__55716;
    wire N__55709;
    wire N__55706;
    wire N__55701;
    wire N__55694;
    wire N__55693;
    wire N__55690;
    wire N__55685;
    wire N__55682;
    wire N__55679;
    wire N__55676;
    wire N__55671;
    wire N__55666;
    wire N__55663;
    wire N__55660;
    wire N__55659;
    wire N__55656;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55642;
    wire N__55641;
    wire N__55640;
    wire N__55631;
    wire N__55626;
    wire N__55623;
    wire N__55618;
    wire N__55609;
    wire N__55604;
    wire N__55601;
    wire N__55598;
    wire N__55589;
    wire N__55586;
    wire N__55585;
    wire N__55582;
    wire N__55579;
    wire N__55574;
    wire N__55567;
    wire N__55564;
    wire N__55555;
    wire N__55552;
    wire N__55537;
    wire N__55536;
    wire N__55535;
    wire N__55534;
    wire N__55533;
    wire N__55530;
    wire N__55529;
    wire N__55528;
    wire N__55527;
    wire N__55524;
    wire N__55523;
    wire N__55522;
    wire N__55521;
    wire N__55518;
    wire N__55517;
    wire N__55514;
    wire N__55513;
    wire N__55510;
    wire N__55507;
    wire N__55506;
    wire N__55503;
    wire N__55500;
    wire N__55497;
    wire N__55492;
    wire N__55491;
    wire N__55490;
    wire N__55489;
    wire N__55488;
    wire N__55485;
    wire N__55482;
    wire N__55481;
    wire N__55480;
    wire N__55477;
    wire N__55476;
    wire N__55473;
    wire N__55468;
    wire N__55465;
    wire N__55462;
    wire N__55459;
    wire N__55458;
    wire N__55449;
    wire N__55448;
    wire N__55447;
    wire N__55446;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55434;
    wire N__55431;
    wire N__55428;
    wire N__55423;
    wire N__55420;
    wire N__55417;
    wire N__55414;
    wire N__55411;
    wire N__55404;
    wire N__55401;
    wire N__55400;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55388;
    wire N__55383;
    wire N__55382;
    wire N__55381;
    wire N__55378;
    wire N__55375;
    wire N__55366;
    wire N__55359;
    wire N__55356;
    wire N__55353;
    wire N__55348;
    wire N__55345;
    wire N__55342;
    wire N__55337;
    wire N__55334;
    wire N__55331;
    wire N__55328;
    wire N__55325;
    wire N__55322;
    wire N__55319;
    wire N__55316;
    wire N__55311;
    wire N__55306;
    wire N__55303;
    wire N__55282;
    wire N__55281;
    wire N__55280;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55272;
    wire N__55269;
    wire N__55268;
    wire N__55265;
    wire N__55264;
    wire N__55263;
    wire N__55262;
    wire N__55261;
    wire N__55260;
    wire N__55259;
    wire N__55256;
    wire N__55253;
    wire N__55250;
    wire N__55247;
    wire N__55244;
    wire N__55241;
    wire N__55238;
    wire N__55235;
    wire N__55234;
    wire N__55231;
    wire N__55230;
    wire N__55227;
    wire N__55224;
    wire N__55223;
    wire N__55222;
    wire N__55221;
    wire N__55220;
    wire N__55217;
    wire N__55216;
    wire N__55205;
    wire N__55202;
    wire N__55199;
    wire N__55196;
    wire N__55193;
    wire N__55192;
    wire N__55189;
    wire N__55186;
    wire N__55185;
    wire N__55182;
    wire N__55179;
    wire N__55176;
    wire N__55173;
    wire N__55172;
    wire N__55169;
    wire N__55168;
    wire N__55167;
    wire N__55166;
    wire N__55163;
    wire N__55162;
    wire N__55159;
    wire N__55156;
    wire N__55153;
    wire N__55150;
    wire N__55143;
    wire N__55142;
    wire N__55139;
    wire N__55138;
    wire N__55133;
    wire N__55130;
    wire N__55123;
    wire N__55120;
    wire N__55117;
    wire N__55114;
    wire N__55111;
    wire N__55108;
    wire N__55105;
    wire N__55102;
    wire N__55099;
    wire N__55098;
    wire N__55095;
    wire N__55092;
    wire N__55085;
    wire N__55082;
    wire N__55079;
    wire N__55076;
    wire N__55073;
    wire N__55072;
    wire N__55071;
    wire N__55068;
    wire N__55065;
    wire N__55062;
    wire N__55057;
    wire N__55048;
    wire N__55045;
    wire N__55042;
    wire N__55035;
    wire N__55030;
    wire N__55027;
    wire N__55024;
    wire N__55021;
    wire N__55018;
    wire N__55015;
    wire N__55008;
    wire N__55003;
    wire N__54998;
    wire N__54991;
    wire N__54976;
    wire N__54973;
    wire N__54972;
    wire N__54969;
    wire N__54966;
    wire N__54961;
    wire N__54960;
    wire N__54959;
    wire N__54958;
    wire N__54957;
    wire N__54956;
    wire N__54955;
    wire N__54940;
    wire N__54937;
    wire N__54936;
    wire N__54933;
    wire N__54930;
    wire N__54925;
    wire N__54924;
    wire N__54923;
    wire N__54922;
    wire N__54921;
    wire N__54920;
    wire N__54919;
    wire N__54916;
    wire N__54915;
    wire N__54914;
    wire N__54911;
    wire N__54908;
    wire N__54907;
    wire N__54906;
    wire N__54905;
    wire N__54902;
    wire N__54901;
    wire N__54900;
    wire N__54899;
    wire N__54898;
    wire N__54895;
    wire N__54894;
    wire N__54891;
    wire N__54890;
    wire N__54889;
    wire N__54888;
    wire N__54887;
    wire N__54886;
    wire N__54885;
    wire N__54884;
    wire N__54881;
    wire N__54878;
    wire N__54871;
    wire N__54864;
    wire N__54861;
    wire N__54860;
    wire N__54859;
    wire N__54858;
    wire N__54855;
    wire N__54850;
    wire N__54843;
    wire N__54838;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54834;
    wire N__54833;
    wire N__54830;
    wire N__54829;
    wire N__54828;
    wire N__54827;
    wire N__54824;
    wire N__54823;
    wire N__54822;
    wire N__54821;
    wire N__54818;
    wire N__54817;
    wire N__54814;
    wire N__54813;
    wire N__54812;
    wire N__54811;
    wire N__54810;
    wire N__54807;
    wire N__54806;
    wire N__54805;
    wire N__54804;
    wire N__54803;
    wire N__54802;
    wire N__54801;
    wire N__54800;
    wire N__54797;
    wire N__54796;
    wire N__54795;
    wire N__54792;
    wire N__54791;
    wire N__54790;
    wire N__54789;
    wire N__54788;
    wire N__54787;
    wire N__54786;
    wire N__54785;
    wire N__54784;
    wire N__54783;
    wire N__54782;
    wire N__54781;
    wire N__54780;
    wire N__54779;
    wire N__54778;
    wire N__54777;
    wire N__54770;
    wire N__54765;
    wire N__54760;
    wire N__54757;
    wire N__54754;
    wire N__54749;
    wire N__54746;
    wire N__54739;
    wire N__54734;
    wire N__54731;
    wire N__54728;
    wire N__54725;
    wire N__54720;
    wire N__54719;
    wire N__54718;
    wire N__54715;
    wire N__54708;
    wire N__54703;
    wire N__54702;
    wire N__54701;
    wire N__54698;
    wire N__54697;
    wire N__54694;
    wire N__54691;
    wire N__54686;
    wire N__54681;
    wire N__54672;
    wire N__54669;
    wire N__54664;
    wire N__54659;
    wire N__54658;
    wire N__54655;
    wire N__54652;
    wire N__54651;
    wire N__54648;
    wire N__54645;
    wire N__54642;
    wire N__54641;
    wire N__54640;
    wire N__54639;
    wire N__54638;
    wire N__54633;
    wire N__54632;
    wire N__54631;
    wire N__54630;
    wire N__54629;
    wire N__54628;
    wire N__54627;
    wire N__54626;
    wire N__54625;
    wire N__54622;
    wire N__54619;
    wire N__54618;
    wire N__54617;
    wire N__54616;
    wire N__54615;
    wire N__54612;
    wire N__54611;
    wire N__54608;
    wire N__54607;
    wire N__54606;
    wire N__54605;
    wire N__54604;
    wire N__54603;
    wire N__54600;
    wire N__54597;
    wire N__54596;
    wire N__54595;
    wire N__54594;
    wire N__54593;
    wire N__54592;
    wire N__54591;
    wire N__54590;
    wire N__54587;
    wire N__54586;
    wire N__54585;
    wire N__54584;
    wire N__54583;
    wire N__54582;
    wire N__54581;
    wire N__54580;
    wire N__54577;
    wire N__54568;
    wire N__54563;
    wire N__54558;
    wire N__54557;
    wire N__54556;
    wire N__54555;
    wire N__54554;
    wire N__54553;
    wire N__54552;
    wire N__54547;
    wire N__54540;
    wire N__54533;
    wire N__54528;
    wire N__54521;
    wire N__54520;
    wire N__54517;
    wire N__54512;
    wire N__54509;
    wire N__54504;
    wire N__54501;
    wire N__54496;
    wire N__54489;
    wire N__54484;
    wire N__54479;
    wire N__54478;
    wire N__54475;
    wire N__54470;
    wire N__54467;
    wire N__54464;
    wire N__54461;
    wire N__54448;
    wire N__54447;
    wire N__54442;
    wire N__54439;
    wire N__54432;
    wire N__54429;
    wire N__54426;
    wire N__54423;
    wire N__54420;
    wire N__54417;
    wire N__54414;
    wire N__54409;
    wire N__54406;
    wire N__54403;
    wire N__54396;
    wire N__54393;
    wire N__54384;
    wire N__54383;
    wire N__54376;
    wire N__54373;
    wire N__54370;
    wire N__54365;
    wire N__54362;
    wire N__54359;
    wire N__54352;
    wire N__54349;
    wire N__54346;
    wire N__54343;
    wire N__54338;
    wire N__54335;
    wire N__54328;
    wire N__54325;
    wire N__54322;
    wire N__54319;
    wire N__54316;
    wire N__54301;
    wire N__54298;
    wire N__54295;
    wire N__54290;
    wire N__54287;
    wire N__54280;
    wire N__54277;
    wire N__54274;
    wire N__54269;
    wire N__54260;
    wire N__54257;
    wire N__54250;
    wire N__54247;
    wire N__54244;
    wire N__54239;
    wire N__54236;
    wire N__54233;
    wire N__54230;
    wire N__54219;
    wire N__54216;
    wire N__54215;
    wire N__54212;
    wire N__54209;
    wire N__54204;
    wire N__54193;
    wire N__54188;
    wire N__54185;
    wire N__54178;
    wire N__54167;
    wire N__54164;
    wire N__54155;
    wire N__54152;
    wire N__54145;
    wire N__54142;
    wire N__54133;
    wire N__54130;
    wire N__54129;
    wire N__54128;
    wire N__54125;
    wire N__54120;
    wire N__54111;
    wire N__54108;
    wire N__54105;
    wire N__54102;
    wire N__54099;
    wire N__54096;
    wire N__54091;
    wire N__54086;
    wire N__54081;
    wire N__54070;
    wire N__54069;
    wire N__54066;
    wire N__54063;
    wire N__54062;
    wire N__54061;
    wire N__54060;
    wire N__54059;
    wire N__54058;
    wire N__54057;
    wire N__54056;
    wire N__54055;
    wire N__54054;
    wire N__54053;
    wire N__54052;
    wire N__54051;
    wire N__54050;
    wire N__54049;
    wire N__54048;
    wire N__54047;
    wire N__54042;
    wire N__54041;
    wire N__54040;
    wire N__54039;
    wire N__54038;
    wire N__54037;
    wire N__54036;
    wire N__54033;
    wire N__54032;
    wire N__54029;
    wire N__54028;
    wire N__54027;
    wire N__54026;
    wire N__54025;
    wire N__54024;
    wire N__54023;
    wire N__54022;
    wire N__54021;
    wire N__54020;
    wire N__54017;
    wire N__54014;
    wire N__54009;
    wire N__54006;
    wire N__54003;
    wire N__54002;
    wire N__54001;
    wire N__54000;
    wire N__53999;
    wire N__53998;
    wire N__53997;
    wire N__53996;
    wire N__53987;
    wire N__53986;
    wire N__53985;
    wire N__53980;
    wire N__53977;
    wire N__53976;
    wire N__53975;
    wire N__53974;
    wire N__53973;
    wire N__53972;
    wire N__53971;
    wire N__53970;
    wire N__53969;
    wire N__53968;
    wire N__53967;
    wire N__53966;
    wire N__53965;
    wire N__53964;
    wire N__53963;
    wire N__53962;
    wire N__53961;
    wire N__53960;
    wire N__53959;
    wire N__53958;
    wire N__53957;
    wire N__53956;
    wire N__53955;
    wire N__53952;
    wire N__53951;
    wire N__53950;
    wire N__53949;
    wire N__53948;
    wire N__53947;
    wire N__53946;
    wire N__53945;
    wire N__53942;
    wire N__53939;
    wire N__53930;
    wire N__53929;
    wire N__53928;
    wire N__53927;
    wire N__53926;
    wire N__53925;
    wire N__53924;
    wire N__53923;
    wire N__53920;
    wire N__53917;
    wire N__53914;
    wire N__53913;
    wire N__53912;
    wire N__53911;
    wire N__53908;
    wire N__53901;
    wire N__53900;
    wire N__53899;
    wire N__53898;
    wire N__53897;
    wire N__53896;
    wire N__53895;
    wire N__53894;
    wire N__53893;
    wire N__53890;
    wire N__53887;
    wire N__53886;
    wire N__53885;
    wire N__53880;
    wire N__53875;
    wire N__53874;
    wire N__53873;
    wire N__53872;
    wire N__53871;
    wire N__53864;
    wire N__53861;
    wire N__53858;
    wire N__53857;
    wire N__53856;
    wire N__53853;
    wire N__53848;
    wire N__53843;
    wire N__53838;
    wire N__53835;
    wire N__53832;
    wire N__53829;
    wire N__53826;
    wire N__53823;
    wire N__53816;
    wire N__53813;
    wire N__53812;
    wire N__53811;
    wire N__53808;
    wire N__53807;
    wire N__53806;
    wire N__53805;
    wire N__53804;
    wire N__53799;
    wire N__53792;
    wire N__53783;
    wire N__53782;
    wire N__53781;
    wire N__53780;
    wire N__53779;
    wire N__53778;
    wire N__53771;
    wire N__53766;
    wire N__53763;
    wire N__53760;
    wire N__53759;
    wire N__53758;
    wire N__53757;
    wire N__53754;
    wire N__53753;
    wire N__53748;
    wire N__53743;
    wire N__53742;
    wire N__53735;
    wire N__53732;
    wire N__53725;
    wire N__53718;
    wire N__53709;
    wire N__53702;
    wire N__53695;
    wire N__53690;
    wire N__53687;
    wire N__53686;
    wire N__53685;
    wire N__53682;
    wire N__53681;
    wire N__53680;
    wire N__53677;
    wire N__53676;
    wire N__53675;
    wire N__53672;
    wire N__53669;
    wire N__53662;
    wire N__53657;
    wire N__53652;
    wire N__53647;
    wire N__53646;
    wire N__53645;
    wire N__53644;
    wire N__53641;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53625;
    wire N__53620;
    wire N__53613;
    wire N__53610;
    wire N__53607;
    wire N__53594;
    wire N__53591;
    wire N__53590;
    wire N__53587;
    wire N__53584;
    wire N__53579;
    wire N__53576;
    wire N__53573;
    wire N__53570;
    wire N__53565;
    wire N__53562;
    wire N__53559;
    wire N__53552;
    wire N__53543;
    wire N__53540;
    wire N__53535;
    wire N__53532;
    wire N__53529;
    wire N__53526;
    wire N__53523;
    wire N__53520;
    wire N__53517;
    wire N__53516;
    wire N__53513;
    wire N__53510;
    wire N__53505;
    wire N__53500;
    wire N__53495;
    wire N__53486;
    wire N__53483;
    wire N__53480;
    wire N__53475;
    wire N__53466;
    wire N__53461;
    wire N__53454;
    wire N__53447;
    wire N__53442;
    wire N__53435;
    wire N__53430;
    wire N__53425;
    wire N__53422;
    wire N__53421;
    wire N__53418;
    wire N__53415;
    wire N__53412;
    wire N__53401;
    wire N__53396;
    wire N__53387;
    wire N__53380;
    wire N__53377;
    wire N__53374;
    wire N__53365;
    wire N__53358;
    wire N__53357;
    wire N__53356;
    wire N__53351;
    wire N__53342;
    wire N__53335;
    wire N__53330;
    wire N__53327;
    wire N__53320;
    wire N__53317;
    wire N__53310;
    wire N__53305;
    wire N__53302;
    wire N__53299;
    wire N__53294;
    wire N__53289;
    wire N__53282;
    wire N__53275;
    wire N__53268;
    wire N__53257;
    wire N__53256;
    wire N__53255;
    wire N__53254;
    wire N__53251;
    wire N__53250;
    wire N__53247;
    wire N__53244;
    wire N__53243;
    wire N__53242;
    wire N__53241;
    wire N__53240;
    wire N__53239;
    wire N__53238;
    wire N__53237;
    wire N__53236;
    wire N__53233;
    wire N__53232;
    wire N__53231;
    wire N__53230;
    wire N__53229;
    wire N__53228;
    wire N__53225;
    wire N__53224;
    wire N__53223;
    wire N__53222;
    wire N__53221;
    wire N__53220;
    wire N__53219;
    wire N__53218;
    wire N__53217;
    wire N__53216;
    wire N__53215;
    wire N__53214;
    wire N__53213;
    wire N__53212;
    wire N__53209;
    wire N__53208;
    wire N__53207;
    wire N__53206;
    wire N__53205;
    wire N__53200;
    wire N__53197;
    wire N__53196;
    wire N__53195;
    wire N__53194;
    wire N__53193;
    wire N__53190;
    wire N__53187;
    wire N__53184;
    wire N__53183;
    wire N__53182;
    wire N__53181;
    wire N__53180;
    wire N__53177;
    wire N__53176;
    wire N__53175;
    wire N__53170;
    wire N__53169;
    wire N__53168;
    wire N__53167;
    wire N__53166;
    wire N__53165;
    wire N__53164;
    wire N__53163;
    wire N__53162;
    wire N__53161;
    wire N__53160;
    wire N__53159;
    wire N__53158;
    wire N__53155;
    wire N__53154;
    wire N__53153;
    wire N__53152;
    wire N__53149;
    wire N__53146;
    wire N__53145;
    wire N__53144;
    wire N__53143;
    wire N__53140;
    wire N__53139;
    wire N__53136;
    wire N__53135;
    wire N__53134;
    wire N__53131;
    wire N__53130;
    wire N__53129;
    wire N__53126;
    wire N__53123;
    wire N__53122;
    wire N__53121;
    wire N__53120;
    wire N__53119;
    wire N__53118;
    wire N__53115;
    wire N__53114;
    wire N__53111;
    wire N__53108;
    wire N__53105;
    wire N__53104;
    wire N__53103;
    wire N__53102;
    wire N__53099;
    wire N__53098;
    wire N__53095;
    wire N__53092;
    wire N__53091;
    wire N__53090;
    wire N__53087;
    wire N__53084;
    wire N__53081;
    wire N__53080;
    wire N__53077;
    wire N__53074;
    wire N__53069;
    wire N__53068;
    wire N__53065;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53052;
    wire N__53045;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53018;
    wire N__53015;
    wire N__53014;
    wire N__53011;
    wire N__53008;
    wire N__53005;
    wire N__53004;
    wire N__53003;
    wire N__53000;
    wire N__52997;
    wire N__52996;
    wire N__52993;
    wire N__52992;
    wire N__52989;
    wire N__52986;
    wire N__52985;
    wire N__52984;
    wire N__52983;
    wire N__52982;
    wire N__52979;
    wire N__52976;
    wire N__52973;
    wire N__52972;
    wire N__52971;
    wire N__52970;
    wire N__52967;
    wire N__52964;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52954;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52941;
    wire N__52940;
    wire N__52939;
    wire N__52938;
    wire N__52937;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52925;
    wire N__52922;
    wire N__52915;
    wire N__52912;
    wire N__52909;
    wire N__52906;
    wire N__52903;
    wire N__52900;
    wire N__52897;
    wire N__52894;
    wire N__52893;
    wire N__52890;
    wire N__52887;
    wire N__52884;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52876;
    wire N__52873;
    wire N__52870;
    wire N__52867;
    wire N__52864;
    wire N__52861;
    wire N__52858;
    wire N__52855;
    wire N__52848;
    wire N__52841;
    wire N__52838;
    wire N__52833;
    wire N__52830;
    wire N__52827;
    wire N__52824;
    wire N__52821;
    wire N__52820;
    wire N__52819;
    wire N__52816;
    wire N__52811;
    wire N__52808;
    wire N__52803;
    wire N__52800;
    wire N__52793;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52775;
    wire N__52766;
    wire N__52759;
    wire N__52742;
    wire N__52741;
    wire N__52738;
    wire N__52735;
    wire N__52732;
    wire N__52729;
    wire N__52726;
    wire N__52723;
    wire N__52720;
    wire N__52719;
    wire N__52718;
    wire N__52713;
    wire N__52710;
    wire N__52703;
    wire N__52700;
    wire N__52697;
    wire N__52694;
    wire N__52691;
    wire N__52688;
    wire N__52683;
    wire N__52674;
    wire N__52669;
    wire N__52664;
    wire N__52657;
    wire N__52654;
    wire N__52647;
    wire N__52640;
    wire N__52633;
    wire N__52630;
    wire N__52625;
    wire N__52620;
    wire N__52617;
    wire N__52610;
    wire N__52605;
    wire N__52602;
    wire N__52599;
    wire N__52598;
    wire N__52593;
    wire N__52586;
    wire N__52581;
    wire N__52574;
    wire N__52567;
    wire N__52564;
    wire N__52561;
    wire N__52558;
    wire N__52555;
    wire N__52550;
    wire N__52545;
    wire N__52544;
    wire N__52541;
    wire N__52538;
    wire N__52537;
    wire N__52534;
    wire N__52531;
    wire N__52526;
    wire N__52523;
    wire N__52520;
    wire N__52517;
    wire N__52512;
    wire N__52509;
    wire N__52498;
    wire N__52491;
    wire N__52486;
    wire N__52483;
    wire N__52474;
    wire N__52469;
    wire N__52466;
    wire N__52463;
    wire N__52456;
    wire N__52449;
    wire N__52448;
    wire N__52447;
    wire N__52444;
    wire N__52437;
    wire N__52434;
    wire N__52429;
    wire N__52426;
    wire N__52419;
    wire N__52416;
    wire N__52401;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52385;
    wire N__52382;
    wire N__52379;
    wire N__52376;
    wire N__52371;
    wire N__52360;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52344;
    wire N__52327;
    wire N__52326;
    wire N__52325;
    wire N__52324;
    wire N__52323;
    wire N__52322;
    wire N__52321;
    wire N__52320;
    wire N__52317;
    wire N__52314;
    wire N__52311;
    wire N__52310;
    wire N__52309;
    wire N__52308;
    wire N__52303;
    wire N__52302;
    wire N__52301;
    wire N__52300;
    wire N__52299;
    wire N__52294;
    wire N__52293;
    wire N__52290;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52278;
    wire N__52277;
    wire N__52276;
    wire N__52275;
    wire N__52272;
    wire N__52269;
    wire N__52266;
    wire N__52263;
    wire N__52260;
    wire N__52257;
    wire N__52256;
    wire N__52255;
    wire N__52254;
    wire N__52253;
    wire N__52250;
    wire N__52247;
    wire N__52244;
    wire N__52241;
    wire N__52232;
    wire N__52229;
    wire N__52228;
    wire N__52223;
    wire N__52222;
    wire N__52221;
    wire N__52218;
    wire N__52215;
    wire N__52212;
    wire N__52205;
    wire N__52200;
    wire N__52199;
    wire N__52198;
    wire N__52195;
    wire N__52192;
    wire N__52189;
    wire N__52184;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52152;
    wire N__52151;
    wire N__52144;
    wire N__52143;
    wire N__52140;
    wire N__52139;
    wire N__52136;
    wire N__52131;
    wire N__52128;
    wire N__52123;
    wire N__52122;
    wire N__52121;
    wire N__52118;
    wire N__52111;
    wire N__52108;
    wire N__52105;
    wire N__52104;
    wire N__52103;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52084;
    wire N__52079;
    wire N__52070;
    wire N__52063;
    wire N__52048;
    wire N__52045;
    wire N__52042;
    wire N__52039;
    wire N__52036;
    wire N__52035;
    wire N__52034;
    wire N__52033;
    wire N__52030;
    wire N__52029;
    wire N__52028;
    wire N__52025;
    wire N__52024;
    wire N__52021;
    wire N__52018;
    wire N__52015;
    wire N__52012;
    wire N__52009;
    wire N__52004;
    wire N__52003;
    wire N__52002;
    wire N__52001;
    wire N__52000;
    wire N__51997;
    wire N__51992;
    wire N__51989;
    wire N__51988;
    wire N__51987;
    wire N__51984;
    wire N__51983;
    wire N__51980;
    wire N__51979;
    wire N__51976;
    wire N__51975;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51959;
    wire N__51958;
    wire N__51953;
    wire N__51950;
    wire N__51947;
    wire N__51944;
    wire N__51941;
    wire N__51940;
    wire N__51939;
    wire N__51936;
    wire N__51933;
    wire N__51928;
    wire N__51923;
    wire N__51920;
    wire N__51919;
    wire N__51918;
    wire N__51917;
    wire N__51914;
    wire N__51909;
    wire N__51908;
    wire N__51905;
    wire N__51902;
    wire N__51899;
    wire N__51896;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51878;
    wire N__51875;
    wire N__51870;
    wire N__51867;
    wire N__51856;
    wire N__51841;
    wire N__51840;
    wire N__51839;
    wire N__51838;
    wire N__51837;
    wire N__51836;
    wire N__51833;
    wire N__51832;
    wire N__51831;
    wire N__51830;
    wire N__51829;
    wire N__51828;
    wire N__51827;
    wire N__51826;
    wire N__51825;
    wire N__51822;
    wire N__51819;
    wire N__51816;
    wire N__51815;
    wire N__51812;
    wire N__51811;
    wire N__51810;
    wire N__51809;
    wire N__51808;
    wire N__51807;
    wire N__51806;
    wire N__51805;
    wire N__51804;
    wire N__51801;
    wire N__51798;
    wire N__51797;
    wire N__51796;
    wire N__51795;
    wire N__51794;
    wire N__51791;
    wire N__51788;
    wire N__51781;
    wire N__51776;
    wire N__51773;
    wire N__51770;
    wire N__51767;
    wire N__51762;
    wire N__51759;
    wire N__51756;
    wire N__51751;
    wire N__51748;
    wire N__51747;
    wire N__51744;
    wire N__51743;
    wire N__51742;
    wire N__51739;
    wire N__51736;
    wire N__51733;
    wire N__51732;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51720;
    wire N__51717;
    wire N__51716;
    wire N__51713;
    wire N__51702;
    wire N__51699;
    wire N__51696;
    wire N__51691;
    wire N__51688;
    wire N__51683;
    wire N__51680;
    wire N__51677;
    wire N__51672;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51660;
    wire N__51653;
    wire N__51652;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51638;
    wire N__51631;
    wire N__51626;
    wire N__51623;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51594;
    wire N__51587;
    wire N__51582;
    wire N__51575;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51541;
    wire N__51538;
    wire N__51537;
    wire N__51534;
    wire N__51533;
    wire N__51532;
    wire N__51531;
    wire N__51530;
    wire N__51529;
    wire N__51528;
    wire N__51527;
    wire N__51524;
    wire N__51523;
    wire N__51522;
    wire N__51521;
    wire N__51520;
    wire N__51519;
    wire N__51518;
    wire N__51515;
    wire N__51514;
    wire N__51513;
    wire N__51510;
    wire N__51509;
    wire N__51508;
    wire N__51507;
    wire N__51504;
    wire N__51501;
    wire N__51500;
    wire N__51499;
    wire N__51498;
    wire N__51495;
    wire N__51492;
    wire N__51491;
    wire N__51488;
    wire N__51485;
    wire N__51484;
    wire N__51483;
    wire N__51482;
    wire N__51479;
    wire N__51476;
    wire N__51475;
    wire N__51474;
    wire N__51473;
    wire N__51472;
    wire N__51469;
    wire N__51466;
    wire N__51465;
    wire N__51462;
    wire N__51457;
    wire N__51454;
    wire N__51447;
    wire N__51446;
    wire N__51443;
    wire N__51442;
    wire N__51441;
    wire N__51438;
    wire N__51435;
    wire N__51430;
    wire N__51427;
    wire N__51424;
    wire N__51423;
    wire N__51420;
    wire N__51415;
    wire N__51414;
    wire N__51411;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51392;
    wire N__51389;
    wire N__51386;
    wire N__51381;
    wire N__51378;
    wire N__51371;
    wire N__51368;
    wire N__51363;
    wire N__51360;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51350;
    wire N__51347;
    wire N__51342;
    wire N__51337;
    wire N__51334;
    wire N__51329;
    wire N__51326;
    wire N__51323;
    wire N__51320;
    wire N__51315;
    wire N__51312;
    wire N__51305;
    wire N__51304;
    wire N__51303;
    wire N__51302;
    wire N__51301;
    wire N__51300;
    wire N__51297;
    wire N__51296;
    wire N__51291;
    wire N__51286;
    wire N__51281;
    wire N__51276;
    wire N__51269;
    wire N__51268;
    wire N__51265;
    wire N__51258;
    wire N__51247;
    wire N__51246;
    wire N__51245;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51231;
    wire N__51228;
    wire N__51225;
    wire N__51224;
    wire N__51223;
    wire N__51222;
    wire N__51221;
    wire N__51218;
    wire N__51213;
    wire N__51212;
    wire N__51205;
    wire N__51202;
    wire N__51199;
    wire N__51196;
    wire N__51193;
    wire N__51190;
    wire N__51185;
    wire N__51182;
    wire N__51179;
    wire N__51172;
    wire N__51167;
    wire N__51164;
    wire N__51159;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51143;
    wire N__51136;
    wire N__51123;
    wire N__51106;
    wire N__51105;
    wire N__51104;
    wire N__51103;
    wire N__51102;
    wire N__51101;
    wire N__51100;
    wire N__51099;
    wire N__51098;
    wire N__51093;
    wire N__51090;
    wire N__51089;
    wire N__51088;
    wire N__51087;
    wire N__51084;
    wire N__51081;
    wire N__51080;
    wire N__51075;
    wire N__51074;
    wire N__51071;
    wire N__51068;
    wire N__51065;
    wire N__51062;
    wire N__51059;
    wire N__51058;
    wire N__51055;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51047;
    wire N__51044;
    wire N__51041;
    wire N__51040;
    wire N__51039;
    wire N__51038;
    wire N__51037;
    wire N__51034;
    wire N__51033;
    wire N__51032;
    wire N__51029;
    wire N__51028;
    wire N__51027;
    wire N__51026;
    wire N__51025;
    wire N__51024;
    wire N__51021;
    wire N__51016;
    wire N__51011;
    wire N__51004;
    wire N__51003;
    wire N__51002;
    wire N__51001;
    wire N__51000;
    wire N__50999;
    wire N__50996;
    wire N__50995;
    wire N__50994;
    wire N__50993;
    wire N__50992;
    wire N__50989;
    wire N__50986;
    wire N__50985;
    wire N__50984;
    wire N__50979;
    wire N__50974;
    wire N__50971;
    wire N__50968;
    wire N__50965;
    wire N__50962;
    wire N__50961;
    wire N__50958;
    wire N__50955;
    wire N__50952;
    wire N__50949;
    wire N__50942;
    wire N__50933;
    wire N__50932;
    wire N__50931;
    wire N__50926;
    wire N__50921;
    wire N__50918;
    wire N__50915;
    wire N__50912;
    wire N__50909;
    wire N__50904;
    wire N__50899;
    wire N__50894;
    wire N__50889;
    wire N__50882;
    wire N__50879;
    wire N__50878;
    wire N__50875;
    wire N__50874;
    wire N__50873;
    wire N__50860;
    wire N__50857;
    wire N__50856;
    wire N__50853;
    wire N__50850;
    wire N__50845;
    wire N__50834;
    wire N__50825;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50810;
    wire N__50803;
    wire N__50800;
    wire N__50795;
    wire N__50792;
    wire N__50773;
    wire N__50772;
    wire N__50769;
    wire N__50766;
    wire N__50765;
    wire N__50762;
    wire N__50759;
    wire N__50756;
    wire N__50753;
    wire N__50752;
    wire N__50749;
    wire N__50744;
    wire N__50741;
    wire N__50740;
    wire N__50737;
    wire N__50734;
    wire N__50731;
    wire N__50728;
    wire N__50719;
    wire N__50716;
    wire N__50713;
    wire N__50710;
    wire N__50707;
    wire N__50706;
    wire N__50705;
    wire N__50702;
    wire N__50701;
    wire N__50700;
    wire N__50697;
    wire N__50694;
    wire N__50691;
    wire N__50686;
    wire N__50683;
    wire N__50680;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50670;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50654;
    wire N__50651;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50637;
    wire N__50634;
    wire N__50623;
    wire N__50622;
    wire N__50621;
    wire N__50618;
    wire N__50615;
    wire N__50612;
    wire N__50611;
    wire N__50610;
    wire N__50607;
    wire N__50604;
    wire N__50601;
    wire N__50596;
    wire N__50593;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50573;
    wire N__50568;
    wire N__50565;
    wire N__50560;
    wire N__50557;
    wire N__50554;
    wire N__50551;
    wire N__50548;
    wire N__50547;
    wire N__50544;
    wire N__50541;
    wire N__50538;
    wire N__50533;
    wire N__50530;
    wire N__50527;
    wire N__50524;
    wire N__50521;
    wire N__50518;
    wire N__50515;
    wire N__50512;
    wire N__50509;
    wire N__50506;
    wire N__50503;
    wire N__50500;
    wire N__50499;
    wire N__50498;
    wire N__50497;
    wire N__50494;
    wire N__50493;
    wire N__50490;
    wire N__50489;
    wire N__50486;
    wire N__50485;
    wire N__50484;
    wire N__50467;
    wire N__50466;
    wire N__50463;
    wire N__50462;
    wire N__50461;
    wire N__50458;
    wire N__50455;
    wire N__50450;
    wire N__50443;
    wire N__50442;
    wire N__50441;
    wire N__50440;
    wire N__50439;
    wire N__50438;
    wire N__50437;
    wire N__50436;
    wire N__50419;
    wire N__50416;
    wire N__50413;
    wire N__50412;
    wire N__50411;
    wire N__50408;
    wire N__50403;
    wire N__50398;
    wire N__50395;
    wire N__50392;
    wire N__50389;
    wire N__50386;
    wire N__50383;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50350;
    wire N__50347;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50308;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50269;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50232;
    wire N__50229;
    wire N__50226;
    wire N__50223;
    wire N__50220;
    wire N__50217;
    wire N__50214;
    wire N__50211;
    wire N__50208;
    wire N__50203;
    wire N__50200;
    wire N__50199;
    wire N__50196;
    wire N__50193;
    wire N__50192;
    wire N__50189;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50175;
    wire N__50172;
    wire N__50171;
    wire N__50168;
    wire N__50163;
    wire N__50160;
    wire N__50159;
    wire N__50156;
    wire N__50153;
    wire N__50150;
    wire N__50145;
    wire N__50142;
    wire N__50137;
    wire N__50136;
    wire N__50129;
    wire N__50126;
    wire N__50123;
    wire N__50120;
    wire N__50115;
    wire N__50110;
    wire N__50107;
    wire N__50104;
    wire N__50103;
    wire N__50100;
    wire N__50097;
    wire N__50094;
    wire N__50091;
    wire N__50088;
    wire N__50085;
    wire N__50082;
    wire N__50079;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50065;
    wire N__50062;
    wire N__50061;
    wire N__50056;
    wire N__50053;
    wire N__50052;
    wire N__50049;
    wire N__50046;
    wire N__50041;
    wire N__50038;
    wire N__50035;
    wire N__50032;
    wire N__50031;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50011;
    wire N__50008;
    wire N__50005;
    wire N__50002;
    wire N__49999;
    wire N__49996;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49978;
    wire N__49975;
    wire N__49974;
    wire N__49971;
    wire N__49970;
    wire N__49969;
    wire N__49968;
    wire N__49967;
    wire N__49964;
    wire N__49961;
    wire N__49958;
    wire N__49955;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49941;
    wire N__49940;
    wire N__49939;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49933;
    wire N__49932;
    wire N__49929;
    wire N__49926;
    wire N__49925;
    wire N__49922;
    wire N__49919;
    wire N__49916;
    wire N__49911;
    wire N__49906;
    wire N__49903;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49881;
    wire N__49874;
    wire N__49871;
    wire N__49868;
    wire N__49865;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49853;
    wire N__49850;
    wire N__49847;
    wire N__49842;
    wire N__49837;
    wire N__49832;
    wire N__49829;
    wire N__49816;
    wire N__49813;
    wire N__49810;
    wire N__49807;
    wire N__49804;
    wire N__49803;
    wire N__49802;
    wire N__49801;
    wire N__49800;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49792;
    wire N__49791;
    wire N__49788;
    wire N__49787;
    wire N__49784;
    wire N__49781;
    wire N__49778;
    wire N__49761;
    wire N__49756;
    wire N__49753;
    wire N__49750;
    wire N__49747;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49739;
    wire N__49734;
    wire N__49733;
    wire N__49732;
    wire N__49731;
    wire N__49730;
    wire N__49727;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49719;
    wire N__49718;
    wire N__49717;
    wire N__49716;
    wire N__49713;
    wire N__49710;
    wire N__49707;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49686;
    wire N__49685;
    wire N__49682;
    wire N__49679;
    wire N__49676;
    wire N__49673;
    wire N__49670;
    wire N__49667;
    wire N__49664;
    wire N__49661;
    wire N__49658;
    wire N__49655;
    wire N__49652;
    wire N__49649;
    wire N__49646;
    wire N__49643;
    wire N__49640;
    wire N__49637;
    wire N__49634;
    wire N__49631;
    wire N__49626;
    wire N__49619;
    wire N__49616;
    wire N__49609;
    wire N__49606;
    wire N__49603;
    wire N__49600;
    wire N__49597;
    wire N__49594;
    wire N__49591;
    wire N__49588;
    wire N__49583;
    wire N__49580;
    wire N__49577;
    wire N__49574;
    wire N__49569;
    wire N__49566;
    wire N__49561;
    wire N__49558;
    wire N__49549;
    wire N__49546;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49534;
    wire N__49531;
    wire N__49528;
    wire N__49525;
    wire N__49522;
    wire N__49519;
    wire N__49516;
    wire N__49513;
    wire N__49512;
    wire N__49509;
    wire N__49506;
    wire N__49501;
    wire N__49498;
    wire N__49495;
    wire N__49492;
    wire N__49489;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49468;
    wire N__49465;
    wire N__49462;
    wire N__49459;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49441;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49426;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49417;
    wire N__49416;
    wire N__49413;
    wire N__49412;
    wire N__49409;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49398;
    wire N__49397;
    wire N__49394;
    wire N__49393;
    wire N__49390;
    wire N__49387;
    wire N__49384;
    wire N__49381;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49367;
    wire N__49366;
    wire N__49365;
    wire N__49364;
    wire N__49363;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49357;
    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49351;
    wire N__49350;
    wire N__49349;
    wire N__49348;
    wire N__49345;
    wire N__49342;
    wire N__49341;
    wire N__49338;
    wire N__49335;
    wire N__49326;
    wire N__49325;
    wire N__49324;
    wire N__49319;
    wire N__49316;
    wire N__49309;
    wire N__49306;
    wire N__49303;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49289;
    wire N__49288;
    wire N__49283;
    wire N__49278;
    wire N__49277;
    wire N__49274;
    wire N__49271;
    wire N__49268;
    wire N__49265;
    wire N__49260;
    wire N__49255;
    wire N__49254;
    wire N__49253;
    wire N__49250;
    wire N__49247;
    wire N__49242;
    wire N__49239;
    wire N__49238;
    wire N__49237;
    wire N__49236;
    wire N__49227;
    wire N__49224;
    wire N__49219;
    wire N__49216;
    wire N__49213;
    wire N__49202;
    wire N__49197;
    wire N__49192;
    wire N__49187;
    wire N__49184;
    wire N__49179;
    wire N__49170;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49140;
    wire N__49137;
    wire N__49136;
    wire N__49133;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49115;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49083;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49073;
    wire N__49070;
    wire N__49067;
    wire N__49064;
    wire N__49061;
    wire N__49058;
    wire N__49055;
    wire N__49054;
    wire N__49049;
    wire N__49046;
    wire N__49043;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49017;
    wire N__49016;
    wire N__49015;
    wire N__49014;
    wire N__49013;
    wire N__49012;
    wire N__49009;
    wire N__49008;
    wire N__49005;
    wire N__49004;
    wire N__49003;
    wire N__49002;
    wire N__49001;
    wire N__49000;
    wire N__48999;
    wire N__48998;
    wire N__48995;
    wire N__48990;
    wire N__48989;
    wire N__48988;
    wire N__48987;
    wire N__48984;
    wire N__48983;
    wire N__48980;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48968;
    wire N__48965;
    wire N__48962;
    wire N__48959;
    wire N__48956;
    wire N__48955;
    wire N__48950;
    wire N__48949;
    wire N__48946;
    wire N__48945;
    wire N__48944;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48936;
    wire N__48935;
    wire N__48934;
    wire N__48933;
    wire N__48932;
    wire N__48929;
    wire N__48928;
    wire N__48927;
    wire N__48926;
    wire N__48923;
    wire N__48922;
    wire N__48921;
    wire N__48920;
    wire N__48917;
    wire N__48916;
    wire N__48915;
    wire N__48914;
    wire N__48913;
    wire N__48912;
    wire N__48911;
    wire N__48910;
    wire N__48909;
    wire N__48908;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48894;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48870;
    wire N__48867;
    wire N__48860;
    wire N__48855;
    wire N__48846;
    wire N__48839;
    wire N__48834;
    wire N__48831;
    wire N__48830;
    wire N__48827;
    wire N__48822;
    wire N__48819;
    wire N__48816;
    wire N__48809;
    wire N__48802;
    wire N__48799;
    wire N__48794;
    wire N__48793;
    wire N__48792;
    wire N__48785;
    wire N__48782;
    wire N__48779;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48763;
    wire N__48762;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48750;
    wire N__48747;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48727;
    wire N__48724;
    wire N__48719;
    wire N__48716;
    wire N__48713;
    wire N__48708;
    wire N__48699;
    wire N__48690;
    wire N__48687;
    wire N__48674;
    wire N__48655;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48649;
    wire N__48648;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48621;
    wire N__48618;
    wire N__48617;
    wire N__48616;
    wire N__48615;
    wire N__48614;
    wire N__48613;
    wire N__48612;
    wire N__48611;
    wire N__48610;
    wire N__48609;
    wire N__48608;
    wire N__48605;
    wire N__48602;
    wire N__48597;
    wire N__48594;
    wire N__48587;
    wire N__48582;
    wire N__48577;
    wire N__48576;
    wire N__48575;
    wire N__48572;
    wire N__48571;
    wire N__48570;
    wire N__48569;
    wire N__48568;
    wire N__48567;
    wire N__48564;
    wire N__48561;
    wire N__48554;
    wire N__48553;
    wire N__48550;
    wire N__48545;
    wire N__48536;
    wire N__48531;
    wire N__48528;
    wire N__48521;
    wire N__48516;
    wire N__48515;
    wire N__48514;
    wire N__48513;
    wire N__48512;
    wire N__48511;
    wire N__48510;
    wire N__48509;
    wire N__48506;
    wire N__48505;
    wire N__48500;
    wire N__48497;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48479;
    wire N__48474;
    wire N__48473;
    wire N__48472;
    wire N__48469;
    wire N__48464;
    wire N__48461;
    wire N__48458;
    wire N__48455;
    wire N__48452;
    wire N__48443;
    wire N__48436;
    wire N__48431;
    wire N__48426;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48399;
    wire N__48396;
    wire N__48395;
    wire N__48392;
    wire N__48391;
    wire N__48390;
    wire N__48387;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48366;
    wire N__48365;
    wire N__48364;
    wire N__48363;
    wire N__48362;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48351;
    wire N__48348;
    wire N__48343;
    wire N__48342;
    wire N__48339;
    wire N__48336;
    wire N__48335;
    wire N__48330;
    wire N__48327;
    wire N__48324;
    wire N__48323;
    wire N__48320;
    wire N__48315;
    wire N__48308;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48296;
    wire N__48293;
    wire N__48292;
    wire N__48291;
    wire N__48290;
    wire N__48289;
    wire N__48288;
    wire N__48285;
    wire N__48282;
    wire N__48279;
    wire N__48274;
    wire N__48271;
    wire N__48264;
    wire N__48261;
    wire N__48258;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48235;
    wire N__48230;
    wire N__48225;
    wire N__48222;
    wire N__48217;
    wire N__48206;
    wire N__48195;
    wire N__48190;
    wire N__48185;
    wire N__48180;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48137;
    wire N__48136;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48094;
    wire N__48091;
    wire N__48088;
    wire N__48085;
    wire N__48082;
    wire N__48079;
    wire N__48078;
    wire N__48077;
    wire N__48076;
    wire N__48073;
    wire N__48070;
    wire N__48065;
    wire N__48062;
    wire N__48061;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48031;
    wire N__48026;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48012;
    wire N__48009;
    wire N__48004;
    wire N__48001;
    wire N__47998;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47986;
    wire N__47983;
    wire N__47980;
    wire N__47977;
    wire N__47976;
    wire N__47973;
    wire N__47970;
    wire N__47969;
    wire N__47966;
    wire N__47963;
    wire N__47960;
    wire N__47959;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47947;
    wire N__47938;
    wire N__47935;
    wire N__47932;
    wire N__47929;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47895;
    wire N__47892;
    wire N__47889;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47875;
    wire N__47872;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47859;
    wire N__47856;
    wire N__47853;
    wire N__47850;
    wire N__47847;
    wire N__47842;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47791;
    wire N__47788;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47764;
    wire N__47763;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47743;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47724;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47712;
    wire N__47709;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47691;
    wire N__47690;
    wire N__47687;
    wire N__47686;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47671;
    wire N__47668;
    wire N__47665;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47645;
    wire N__47642;
    wire N__47639;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47593;
    wire N__47588;
    wire N__47581;
    wire N__47578;
    wire N__47577;
    wire N__47576;
    wire N__47573;
    wire N__47570;
    wire N__47569;
    wire N__47566;
    wire N__47561;
    wire N__47560;
    wire N__47559;
    wire N__47556;
    wire N__47553;
    wire N__47550;
    wire N__47547;
    wire N__47544;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47482;
    wire N__47479;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47474;
    wire N__47473;
    wire N__47472;
    wire N__47471;
    wire N__47470;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47458;
    wire N__47457;
    wire N__47456;
    wire N__47455;
    wire N__47452;
    wire N__47449;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47426;
    wire N__47425;
    wire N__47424;
    wire N__47423;
    wire N__47420;
    wire N__47417;
    wire N__47414;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47398;
    wire N__47395;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47377;
    wire N__47374;
    wire N__47369;
    wire N__47366;
    wire N__47361;
    wire N__47358;
    wire N__47353;
    wire N__47352;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47342;
    wire N__47335;
    wire N__47330;
    wire N__47325;
    wire N__47322;
    wire N__47317;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47287;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47266;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47233;
    wire N__47230;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47209;
    wire N__47206;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47196;
    wire N__47195;
    wire N__47194;
    wire N__47191;
    wire N__47186;
    wire N__47185;
    wire N__47184;
    wire N__47183;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47166;
    wire N__47163;
    wire N__47160;
    wire N__47153;
    wire N__47150;
    wire N__47149;
    wire N__47148;
    wire N__47145;
    wire N__47140;
    wire N__47139;
    wire N__47136;
    wire N__47133;
    wire N__47128;
    wire N__47125;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47112;
    wire N__47107;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47081;
    wire N__47076;
    wire N__47071;
    wire N__47070;
    wire N__47067;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47056;
    wire N__47053;
    wire N__47052;
    wire N__47051;
    wire N__47050;
    wire N__47047;
    wire N__47046;
    wire N__47045;
    wire N__47042;
    wire N__47041;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47033;
    wire N__47032;
    wire N__47031;
    wire N__47030;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47011;
    wire N__47010;
    wire N__47009;
    wire N__47008;
    wire N__47007;
    wire N__47004;
    wire N__47003;
    wire N__47002;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46992;
    wire N__46989;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46977;
    wire N__46974;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46959;
    wire N__46956;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46933;
    wire N__46930;
    wire N__46925;
    wire N__46922;
    wire N__46919;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46891;
    wire N__46886;
    wire N__46883;
    wire N__46870;
    wire N__46867;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46833;
    wire N__46832;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46811;
    wire N__46808;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46802;
    wire N__46799;
    wire N__46798;
    wire N__46797;
    wire N__46796;
    wire N__46795;
    wire N__46794;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46782;
    wire N__46781;
    wire N__46780;
    wire N__46779;
    wire N__46778;
    wire N__46777;
    wire N__46776;
    wire N__46775;
    wire N__46772;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46754;
    wire N__46751;
    wire N__46750;
    wire N__46749;
    wire N__46748;
    wire N__46747;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46723;
    wire N__46714;
    wire N__46711;
    wire N__46710;
    wire N__46705;
    wire N__46702;
    wire N__46699;
    wire N__46694;
    wire N__46693;
    wire N__46690;
    wire N__46687;
    wire N__46684;
    wire N__46681;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46673;
    wire N__46672;
    wire N__46671;
    wire N__46670;
    wire N__46663;
    wire N__46660;
    wire N__46655;
    wire N__46652;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46631;
    wire N__46626;
    wire N__46621;
    wire N__46618;
    wire N__46615;
    wire N__46612;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46598;
    wire N__46595;
    wire N__46586;
    wire N__46575;
    wire N__46572;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46522;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46502;
    wire N__46497;
    wire N__46494;
    wire N__46493;
    wire N__46488;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46461;
    wire N__46460;
    wire N__46457;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46433;
    wire N__46432;
    wire N__46431;
    wire N__46426;
    wire N__46423;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46412;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46400;
    wire N__46397;
    wire N__46392;
    wire N__46387;
    wire N__46384;
    wire N__46383;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46375;
    wire N__46372;
    wire N__46367;
    wire N__46364;
    wire N__46363;
    wire N__46360;
    wire N__46355;
    wire N__46352;
    wire N__46349;
    wire N__46348;
    wire N__46345;
    wire N__46340;
    wire N__46337;
    wire N__46336;
    wire N__46335;
    wire N__46334;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46317;
    wire N__46316;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46308;
    wire N__46307;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46276;
    wire N__46269;
    wire N__46264;
    wire N__46261;
    wire N__46256;
    wire N__46245;
    wire N__46228;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46220;
    wire N__46219;
    wire N__46218;
    wire N__46217;
    wire N__46216;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46204;
    wire N__46201;
    wire N__46200;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46188;
    wire N__46183;
    wire N__46182;
    wire N__46181;
    wire N__46180;
    wire N__46179;
    wire N__46178;
    wire N__46177;
    wire N__46174;
    wire N__46173;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46162;
    wire N__46161;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46153;
    wire N__46152;
    wire N__46151;
    wire N__46148;
    wire N__46143;
    wire N__46140;
    wire N__46139;
    wire N__46136;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46120;
    wire N__46115;
    wire N__46112;
    wire N__46109;
    wire N__46104;
    wire N__46103;
    wire N__46100;
    wire N__46097;
    wire N__46094;
    wire N__46091;
    wire N__46086;
    wire N__46081;
    wire N__46080;
    wire N__46075;
    wire N__46074;
    wire N__46073;
    wire N__46070;
    wire N__46063;
    wire N__46056;
    wire N__46055;
    wire N__46052;
    wire N__46047;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46016;
    wire N__46013;
    wire N__46010;
    wire N__46009;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45989;
    wire N__45988;
    wire N__45983;
    wire N__45980;
    wire N__45971;
    wire N__45966;
    wire N__45957;
    wire N__45954;
    wire N__45947;
    wire N__45944;
    wire N__45941;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45901;
    wire N__45898;
    wire N__45895;
    wire N__45892;
    wire N__45889;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45846;
    wire N__45843;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45805;
    wire N__45802;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45766;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45748;
    wire N__45745;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45700;
    wire N__45697;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45687;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45673;
    wire N__45670;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45658;
    wire N__45655;
    wire N__45650;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45636;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45595;
    wire N__45592;
    wire N__45589;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45568;
    wire N__45565;
    wire N__45562;
    wire N__45559;
    wire N__45556;
    wire N__45553;
    wire N__45550;
    wire N__45547;
    wire N__45544;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45513;
    wire N__45512;
    wire N__45511;
    wire N__45510;
    wire N__45507;
    wire N__45506;
    wire N__45505;
    wire N__45504;
    wire N__45501;
    wire N__45500;
    wire N__45497;
    wire N__45496;
    wire N__45495;
    wire N__45494;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45484;
    wire N__45483;
    wire N__45480;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45463;
    wire N__45462;
    wire N__45461;
    wire N__45458;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45440;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45426;
    wire N__45419;
    wire N__45418;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45406;
    wire N__45405;
    wire N__45404;
    wire N__45401;
    wire N__45398;
    wire N__45395;
    wire N__45392;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45384;
    wire N__45383;
    wire N__45380;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45362;
    wire N__45361;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45349;
    wire N__45346;
    wire N__45341;
    wire N__45334;
    wire N__45331;
    wire N__45328;
    wire N__45325;
    wire N__45322;
    wire N__45317;
    wire N__45312;
    wire N__45305;
    wire N__45300;
    wire N__45297;
    wire N__45288;
    wire N__45285;
    wire N__45262;
    wire N__45261;
    wire N__45260;
    wire N__45259;
    wire N__45258;
    wire N__45257;
    wire N__45254;
    wire N__45251;
    wire N__45250;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45237;
    wire N__45234;
    wire N__45233;
    wire N__45232;
    wire N__45231;
    wire N__45230;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45222;
    wire N__45219;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45207;
    wire N__45206;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45196;
    wire N__45195;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45189;
    wire N__45188;
    wire N__45185;
    wire N__45182;
    wire N__45181;
    wire N__45180;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45167;
    wire N__45164;
    wire N__45159;
    wire N__45156;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45142;
    wire N__45137;
    wire N__45134;
    wire N__45129;
    wire N__45128;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45107;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45089;
    wire N__45086;
    wire N__45081;
    wire N__45078;
    wire N__45073;
    wire N__45070;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45047;
    wire N__45042;
    wire N__45035;
    wire N__45028;
    wire N__45013;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45005;
    wire N__45002;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44917;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44889;
    wire N__44888;
    wire N__44885;
    wire N__44882;
    wire N__44879;
    wire N__44872;
    wire N__44869;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44844;
    wire N__44843;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44827;
    wire N__44824;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44814;
    wire N__44811;
    wire N__44806;
    wire N__44805;
    wire N__44802;
    wire N__44801;
    wire N__44798;
    wire N__44797;
    wire N__44794;
    wire N__44791;
    wire N__44790;
    wire N__44789;
    wire N__44788;
    wire N__44785;
    wire N__44784;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44766;
    wire N__44765;
    wire N__44764;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44750;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44723;
    wire N__44720;
    wire N__44719;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44705;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44678;
    wire N__44677;
    wire N__44676;
    wire N__44675;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44656;
    wire N__44645;
    wire N__44640;
    wire N__44631;
    wire N__44628;
    wire N__44611;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44603;
    wire N__44602;
    wire N__44601;
    wire N__44600;
    wire N__44597;
    wire N__44596;
    wire N__44595;
    wire N__44594;
    wire N__44593;
    wire N__44590;
    wire N__44589;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44553;
    wire N__44552;
    wire N__44551;
    wire N__44550;
    wire N__44549;
    wire N__44546;
    wire N__44545;
    wire N__44544;
    wire N__44543;
    wire N__44542;
    wire N__44539;
    wire N__44538;
    wire N__44537;
    wire N__44532;
    wire N__44531;
    wire N__44530;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44519;
    wire N__44518;
    wire N__44509;
    wire N__44506;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44490;
    wire N__44489;
    wire N__44488;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44478;
    wire N__44473;
    wire N__44470;
    wire N__44465;
    wire N__44462;
    wire N__44455;
    wire N__44450;
    wire N__44449;
    wire N__44448;
    wire N__44447;
    wire N__44446;
    wire N__44441;
    wire N__44436;
    wire N__44435;
    wire N__44430;
    wire N__44423;
    wire N__44406;
    wire N__44403;
    wire N__44394;
    wire N__44389;
    wire N__44386;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44361;
    wire N__44360;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44352;
    wire N__44351;
    wire N__44350;
    wire N__44349;
    wire N__44348;
    wire N__44347;
    wire N__44346;
    wire N__44345;
    wire N__44344;
    wire N__44343;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44335;
    wire N__44332;
    wire N__44329;
    wire N__44322;
    wire N__44319;
    wire N__44314;
    wire N__44313;
    wire N__44310;
    wire N__44309;
    wire N__44308;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44276;
    wire N__44275;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44260;
    wire N__44253;
    wire N__44252;
    wire N__44251;
    wire N__44250;
    wire N__44249;
    wire N__44248;
    wire N__44241;
    wire N__44234;
    wire N__44227;
    wire N__44222;
    wire N__44215;
    wire N__44210;
    wire N__44203;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44169;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44159;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44141;
    wire N__44136;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44095;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44056;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44041;
    wire N__44038;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44014;
    wire N__44013;
    wire N__44010;
    wire N__44009;
    wire N__44008;
    wire N__44005;
    wire N__44002;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43985;
    wire N__43982;
    wire N__43977;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43962;
    wire N__43961;
    wire N__43958;
    wire N__43955;
    wire N__43954;
    wire N__43951;
    wire N__43950;
    wire N__43949;
    wire N__43948;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43937;
    wire N__43936;
    wire N__43933;
    wire N__43932;
    wire N__43931;
    wire N__43930;
    wire N__43929;
    wire N__43928;
    wire N__43921;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43915;
    wire N__43914;
    wire N__43909;
    wire N__43904;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43898;
    wire N__43897;
    wire N__43896;
    wire N__43893;
    wire N__43888;
    wire N__43887;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43877;
    wire N__43874;
    wire N__43871;
    wire N__43868;
    wire N__43863;
    wire N__43862;
    wire N__43861;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43837;
    wire N__43834;
    wire N__43829;
    wire N__43824;
    wire N__43823;
    wire N__43822;
    wire N__43821;
    wire N__43820;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43812;
    wire N__43809;
    wire N__43804;
    wire N__43799;
    wire N__43794;
    wire N__43789;
    wire N__43782;
    wire N__43777;
    wire N__43774;
    wire N__43767;
    wire N__43760;
    wire N__43751;
    wire N__43744;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43686;
    wire N__43683;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43668;
    wire N__43667;
    wire N__43666;
    wire N__43665;
    wire N__43664;
    wire N__43661;
    wire N__43658;
    wire N__43657;
    wire N__43656;
    wire N__43655;
    wire N__43652;
    wire N__43651;
    wire N__43650;
    wire N__43649;
    wire N__43648;
    wire N__43645;
    wire N__43644;
    wire N__43643;
    wire N__43640;
    wire N__43639;
    wire N__43638;
    wire N__43637;
    wire N__43636;
    wire N__43635;
    wire N__43632;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43608;
    wire N__43607;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43590;
    wire N__43589;
    wire N__43586;
    wire N__43581;
    wire N__43576;
    wire N__43571;
    wire N__43570;
    wire N__43567;
    wire N__43562;
    wire N__43559;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43522;
    wire N__43521;
    wire N__43520;
    wire N__43517;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43495;
    wire N__43492;
    wire N__43487;
    wire N__43484;
    wire N__43473;
    wire N__43468;
    wire N__43463;
    wire N__43460;
    wire N__43449;
    wire N__43438;
    wire N__43437;
    wire N__43436;
    wire N__43435;
    wire N__43432;
    wire N__43431;
    wire N__43430;
    wire N__43429;
    wire N__43426;
    wire N__43425;
    wire N__43424;
    wire N__43421;
    wire N__43420;
    wire N__43417;
    wire N__43416;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43408;
    wire N__43405;
    wire N__43404;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43395;
    wire N__43394;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43380;
    wire N__43379;
    wire N__43378;
    wire N__43377;
    wire N__43376;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43355;
    wire N__43352;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43333;
    wire N__43330;
    wire N__43325;
    wire N__43320;
    wire N__43315;
    wire N__43310;
    wire N__43309;
    wire N__43308;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43284;
    wire N__43283;
    wire N__43282;
    wire N__43281;
    wire N__43280;
    wire N__43279;
    wire N__43276;
    wire N__43269;
    wire N__43266;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43247;
    wire N__43242;
    wire N__43239;
    wire N__43228;
    wire N__43221;
    wire N__43218;
    wire N__43213;
    wire N__43202;
    wire N__43199;
    wire N__43194;
    wire N__43189;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43128;
    wire N__43127;
    wire N__43124;
    wire N__43123;
    wire N__43118;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43092;
    wire N__43089;
    wire N__43086;
    wire N__43079;
    wire N__43076;
    wire N__43071;
    wire N__43066;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43055;
    wire N__43054;
    wire N__43049;
    wire N__43046;
    wire N__43043;
    wire N__43038;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43011;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42993;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42915;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42897;
    wire N__42896;
    wire N__42893;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42867;
    wire N__42866;
    wire N__42863;
    wire N__42862;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42851;
    wire N__42850;
    wire N__42849;
    wire N__42848;
    wire N__42845;
    wire N__42844;
    wire N__42843;
    wire N__42842;
    wire N__42839;
    wire N__42838;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42827;
    wire N__42826;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42818;
    wire N__42817;
    wire N__42816;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42804;
    wire N__42801;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42782;
    wire N__42779;
    wire N__42774;
    wire N__42771;
    wire N__42766;
    wire N__42759;
    wire N__42756;
    wire N__42755;
    wire N__42754;
    wire N__42753;
    wire N__42752;
    wire N__42747;
    wire N__42744;
    wire N__42739;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42727;
    wire N__42726;
    wire N__42725;
    wire N__42724;
    wire N__42723;
    wire N__42720;
    wire N__42715;
    wire N__42712;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42691;
    wire N__42686;
    wire N__42683;
    wire N__42678;
    wire N__42675;
    wire N__42670;
    wire N__42663;
    wire N__42660;
    wire N__42655;
    wire N__42650;
    wire N__42645;
    wire N__42642;
    wire N__42635;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42562;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42550;
    wire N__42547;
    wire N__42544;
    wire N__42541;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42469;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42454;
    wire N__42451;
    wire N__42448;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42440;
    wire N__42437;
    wire N__42434;
    wire N__42431;
    wire N__42430;
    wire N__42427;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42399;
    wire N__42396;
    wire N__42395;
    wire N__42392;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42374;
    wire N__42369;
    wire N__42366;
    wire N__42361;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42343;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42322;
    wire N__42321;
    wire N__42318;
    wire N__42317;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42305;
    wire N__42298;
    wire N__42295;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42283;
    wire N__42280;
    wire N__42279;
    wire N__42274;
    wire N__42271;
    wire N__42268;
    wire N__42267;
    wire N__42266;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42231;
    wire N__42226;
    wire N__42223;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42208;
    wire N__42205;
    wire N__42204;
    wire N__42203;
    wire N__42200;
    wire N__42199;
    wire N__42194;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42156;
    wire N__42155;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42147;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42139;
    wire N__42136;
    wire N__42133;
    wire N__42130;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42073;
    wire N__42070;
    wire N__42061;
    wire N__42058;
    wire N__42057;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42043;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41968;
    wire N__41965;
    wire N__41962;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41952;
    wire N__41951;
    wire N__41948;
    wire N__41943;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41933;
    wire N__41928;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41884;
    wire N__41881;
    wire N__41878;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41824;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41727;
    wire N__41726;
    wire N__41723;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41707;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41687;
    wire N__41686;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41674;
    wire N__41671;
    wire N__41662;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41650;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41629;
    wire N__41626;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41607;
    wire N__41602;
    wire N__41599;
    wire N__41596;
    wire N__41593;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41571;
    wire N__41570;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41562;
    wire N__41561;
    wire N__41558;
    wire N__41557;
    wire N__41556;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41548;
    wire N__41545;
    wire N__41544;
    wire N__41543;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41520;
    wire N__41517;
    wire N__41512;
    wire N__41505;
    wire N__41504;
    wire N__41503;
    wire N__41502;
    wire N__41501;
    wire N__41500;
    wire N__41499;
    wire N__41498;
    wire N__41493;
    wire N__41490;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41468;
    wire N__41465;
    wire N__41464;
    wire N__41449;
    wire N__41446;
    wire N__41445;
    wire N__41442;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41408;
    wire N__41405;
    wire N__41400;
    wire N__41395;
    wire N__41390;
    wire N__41387;
    wire N__41368;
    wire N__41367;
    wire N__41366;
    wire N__41365;
    wire N__41364;
    wire N__41363;
    wire N__41362;
    wire N__41359;
    wire N__41358;
    wire N__41357;
    wire N__41356;
    wire N__41355;
    wire N__41354;
    wire N__41353;
    wire N__41352;
    wire N__41351;
    wire N__41350;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41329;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41317;
    wire N__41316;
    wire N__41315;
    wire N__41314;
    wire N__41311;
    wire N__41306;
    wire N__41303;
    wire N__41302;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41294;
    wire N__41293;
    wire N__41290;
    wire N__41285;
    wire N__41282;
    wire N__41277;
    wire N__41276;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41248;
    wire N__41243;
    wire N__41240;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41180;
    wire N__41173;
    wire N__41170;
    wire N__41167;
    wire N__41162;
    wire N__41155;
    wire N__41150;
    wire N__41145;
    wire N__41140;
    wire N__41135;
    wire N__41132;
    wire N__41119;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41091;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41025;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40992;
    wire N__40991;
    wire N__40990;
    wire N__40989;
    wire N__40988;
    wire N__40987;
    wire N__40986;
    wire N__40983;
    wire N__40982;
    wire N__40981;
    wire N__40974;
    wire N__40971;
    wire N__40970;
    wire N__40969;
    wire N__40968;
    wire N__40967;
    wire N__40966;
    wire N__40965;
    wire N__40964;
    wire N__40963;
    wire N__40962;
    wire N__40961;
    wire N__40960;
    wire N__40959;
    wire N__40958;
    wire N__40957;
    wire N__40956;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40932;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40912;
    wire N__40911;
    wire N__40908;
    wire N__40901;
    wire N__40898;
    wire N__40893;
    wire N__40892;
    wire N__40889;
    wire N__40886;
    wire N__40883;
    wire N__40878;
    wire N__40877;
    wire N__40876;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40862;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40829;
    wire N__40824;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40806;
    wire N__40793;
    wire N__40788;
    wire N__40785;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40732;
    wire N__40731;
    wire N__40730;
    wire N__40727;
    wire N__40722;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40704;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40694;
    wire N__40691;
    wire N__40688;
    wire N__40687;
    wire N__40684;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40607;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40587;
    wire N__40584;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40533;
    wire N__40532;
    wire N__40531;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40523;
    wire N__40522;
    wire N__40521;
    wire N__40520;
    wire N__40519;
    wire N__40518;
    wire N__40513;
    wire N__40512;
    wire N__40511;
    wire N__40510;
    wire N__40509;
    wire N__40508;
    wire N__40505;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40489;
    wire N__40488;
    wire N__40487;
    wire N__40486;
    wire N__40485;
    wire N__40482;
    wire N__40477;
    wire N__40474;
    wire N__40469;
    wire N__40466;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40434;
    wire N__40433;
    wire N__40432;
    wire N__40431;
    wire N__40430;
    wire N__40429;
    wire N__40428;
    wire N__40425;
    wire N__40420;
    wire N__40415;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40394;
    wire N__40391;
    wire N__40386;
    wire N__40381;
    wire N__40376;
    wire N__40371;
    wire N__40366;
    wire N__40361;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40289;
    wire N__40288;
    wire N__40287;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40275;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40244;
    wire N__40243;
    wire N__40240;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40182;
    wire N__40177;
    wire N__40176;
    wire N__40175;
    wire N__40174;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40160;
    wire N__40159;
    wire N__40158;
    wire N__40157;
    wire N__40156;
    wire N__40155;
    wire N__40154;
    wire N__40151;
    wire N__40146;
    wire N__40143;
    wire N__40142;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40120;
    wire N__40115;
    wire N__40114;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40106;
    wire N__40103;
    wire N__40098;
    wire N__40097;
    wire N__40092;
    wire N__40087;
    wire N__40086;
    wire N__40085;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40055;
    wire N__40054;
    wire N__40049;
    wire N__40046;
    wire N__40039;
    wire N__40036;
    wire N__40025;
    wire N__40022;
    wire N__40009;
    wire N__40008;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39994;
    wire N__39993;
    wire N__39992;
    wire N__39989;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39981;
    wire N__39974;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39946;
    wire N__39943;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39910;
    wire N__39907;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39876;
    wire N__39875;
    wire N__39874;
    wire N__39873;
    wire N__39872;
    wire N__39867;
    wire N__39864;
    wire N__39863;
    wire N__39862;
    wire N__39861;
    wire N__39860;
    wire N__39859;
    wire N__39854;
    wire N__39851;
    wire N__39850;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39838;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39830;
    wire N__39827;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39814;
    wire N__39813;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39783;
    wire N__39780;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39747;
    wire N__39744;
    wire N__39739;
    wire N__39732;
    wire N__39727;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39700;
    wire N__39697;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39618;
    wire N__39617;
    wire N__39616;
    wire N__39613;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39597;
    wire N__39594;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39525;
    wire N__39524;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39494;
    wire N__39493;
    wire N__39490;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39439;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39431;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39403;
    wire N__39402;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39391;
    wire N__39388;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39317;
    wire N__39312;
    wire N__39309;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39202;
    wire N__39201;
    wire N__39200;
    wire N__39197;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39169;
    wire N__39168;
    wire N__39167;
    wire N__39164;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39132;
    wire N__39129;
    wire N__39128;
    wire N__39125;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39091;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39083;
    wire N__39082;
    wire N__39079;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39052;
    wire N__39047;
    wire N__39044;
    wire N__39043;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39010;
    wire N__39001;
    wire N__39000;
    wire N__38999;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38874;
    wire N__38873;
    wire N__38872;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38855;
    wire N__38850;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38828;
    wire N__38827;
    wire N__38824;
    wire N__38819;
    wire N__38816;
    wire N__38815;
    wire N__38808;
    wire N__38805;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38747;
    wire N__38742;
    wire N__38741;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38727;
    wire N__38724;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38712;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38683;
    wire N__38682;
    wire N__38681;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38632;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38548;
    wire N__38545;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38520;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38467;
    wire N__38464;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38452;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38344;
    wire N__38341;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38258;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38222;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38205;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38186;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38076;
    wire N__38075;
    wire N__38072;
    wire N__38067;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38052;
    wire N__38051;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38039;
    wire N__38032;
    wire N__38031;
    wire N__38030;
    wire N__38029;
    wire N__38028;
    wire N__38027;
    wire N__38026;
    wire N__38025;
    wire N__38022;
    wire N__38021;
    wire N__38020;
    wire N__38019;
    wire N__38018;
    wire N__38017;
    wire N__38016;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38008;
    wire N__38007;
    wire N__38002;
    wire N__37995;
    wire N__37994;
    wire N__37993;
    wire N__37992;
    wire N__37989;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37977;
    wire N__37974;
    wire N__37973;
    wire N__37970;
    wire N__37969;
    wire N__37968;
    wire N__37967;
    wire N__37966;
    wire N__37965;
    wire N__37964;
    wire N__37961;
    wire N__37960;
    wire N__37955;
    wire N__37950;
    wire N__37945;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37908;
    wire N__37903;
    wire N__37900;
    wire N__37899;
    wire N__37898;
    wire N__37897;
    wire N__37896;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37888;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37875;
    wire N__37870;
    wire N__37867;
    wire N__37860;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37842;
    wire N__37837;
    wire N__37832;
    wire N__37831;
    wire N__37830;
    wire N__37829;
    wire N__37828;
    wire N__37827;
    wire N__37826;
    wire N__37823;
    wire N__37814;
    wire N__37811;
    wire N__37804;
    wire N__37799;
    wire N__37794;
    wire N__37789;
    wire N__37784;
    wire N__37775;
    wire N__37756;
    wire N__37753;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37735;
    wire N__37734;
    wire N__37731;
    wire N__37730;
    wire N__37727;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37709;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37693;
    wire N__37690;
    wire N__37689;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37637;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37576;
    wire N__37573;
    wire N__37568;
    wire N__37565;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37438;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37212;
    wire N__37211;
    wire N__37210;
    wire N__37209;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37189;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37138;
    wire N__37129;
    wire N__37126;
    wire N__37125;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37089;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36918;
    wire N__36917;
    wire N__36914;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36784;
    wire N__36783;
    wire N__36782;
    wire N__36779;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36771;
    wire N__36770;
    wire N__36769;
    wire N__36768;
    wire N__36767;
    wire N__36766;
    wire N__36765;
    wire N__36764;
    wire N__36763;
    wire N__36760;
    wire N__36759;
    wire N__36756;
    wire N__36755;
    wire N__36754;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36689;
    wire N__36686;
    wire N__36685;
    wire N__36682;
    wire N__36681;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36664;
    wire N__36661;
    wire N__36656;
    wire N__36651;
    wire N__36648;
    wire N__36645;
    wire N__36640;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36585;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36564;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36534;
    wire N__36531;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36515;
    wire N__36508;
    wire N__36505;
    wire N__36500;
    wire N__36487;
    wire N__36486;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36440;
    wire N__36439;
    wire N__36434;
    wire N__36429;
    wire N__36426;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36252;
    wire N__36249;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36147;
    wire N__36142;
    wire N__36141;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36101;
    wire N__36100;
    wire N__36097;
    wire N__36094;
    wire N__36091;
    wire N__36088;
    wire N__36081;
    wire N__36078;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36014;
    wire N__36013;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35834;
    wire N__35833;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35772;
    wire N__35769;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35752;
    wire N__35749;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35637;
    wire N__35636;
    wire N__35633;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35615;
    wire N__35608;
    wire N__35605;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35595;
    wire N__35594;
    wire N__35593;
    wire N__35592;
    wire N__35589;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35581;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35577;
    wire N__35574;
    wire N__35573;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35567;
    wire N__35566;
    wire N__35563;
    wire N__35562;
    wire N__35559;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35541;
    wire N__35540;
    wire N__35539;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35507;
    wire N__35502;
    wire N__35501;
    wire N__35500;
    wire N__35497;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35483;
    wire N__35478;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35460;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35425;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35411;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35393;
    wire N__35392;
    wire N__35389;
    wire N__35388;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35374;
    wire N__35373;
    wire N__35368;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35348;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35313;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35297;
    wire N__35296;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35274;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35115;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35053;
    wire N__35050;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35042;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35026;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35018;
    wire N__35013;
    wire N__35010;
    wire N__35009;
    wire N__35004;
    wire N__35001;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34942;
    wire N__34941;
    wire N__34936;
    wire N__34933;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34854;
    wire N__34853;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34699;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34579;
    wire N__34576;
    wire N__34571;
    wire N__34568;
    wire N__34563;
    wire N__34560;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34405;
    wire N__34402;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34374;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34338;
    wire N__34333;
    wire N__34330;
    wire N__34329;
    wire N__34326;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34305;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34290;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34263;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34089;
    wire N__34084;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34038;
    wire N__34033;
    wire N__34032;
    wire N__34031;
    wire N__34028;
    wire N__34027;
    wire N__34026;
    wire N__34023;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34015;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33983;
    wire N__33978;
    wire N__33969;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33753;
    wire N__33748;
    wire N__33745;
    wire N__33744;
    wire N__33739;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33717;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33699;
    wire N__33696;
    wire N__33691;
    wire N__33688;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33664;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33586;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33468;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33442;
    wire N__33439;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33411;
    wire N__33408;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33388;
    wire N__33385;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33352;
    wire N__33349;
    wire N__33348;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33304;
    wire N__33303;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33285;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33237;
    wire N__33234;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33205;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33161;
    wire N__33156;
    wire N__33153;
    wire N__33142;
    wire N__33141;
    wire N__33140;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33132;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33114;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33057;
    wire N__33056;
    wire N__33053;
    wire N__33048;
    wire N__33045;
    wire N__33040;
    wire N__33037;
    wire N__33036;
    wire N__33031;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32955;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32940;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32888;
    wire N__32887;
    wire N__32884;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32864;
    wire N__32863;
    wire N__32862;
    wire N__32861;
    wire N__32856;
    wire N__32853;
    wire N__32842;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32834;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32817;
    wire N__32816;
    wire N__32815;
    wire N__32812;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32788;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32768;
    wire N__32763;
    wire N__32752;
    wire N__32749;
    wire N__32748;
    wire N__32745;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32719;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32692;
    wire N__32691;
    wire N__32686;
    wire N__32685;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32677;
    wire N__32676;
    wire N__32675;
    wire N__32672;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32660;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32624;
    wire N__32621;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32605;
    wire N__32602;
    wire N__32593;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32575;
    wire N__32574;
    wire N__32571;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32549;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32526;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32487;
    wire N__32476;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32465;
    wire N__32464;
    wire N__32461;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32453;
    wire N__32448;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32407;
    wire N__32402;
    wire N__32397;
    wire N__32394;
    wire N__32389;
    wire N__32384;
    wire N__32377;
    wire N__32376;
    wire N__32375;
    wire N__32374;
    wire N__32373;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32350;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32295;
    wire N__32290;
    wire N__32283;
    wire N__32278;
    wire N__32277;
    wire N__32276;
    wire N__32273;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32265;
    wire N__32264;
    wire N__32263;
    wire N__32262;
    wire N__32261;
    wire N__32258;
    wire N__32257;
    wire N__32254;
    wire N__32249;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32238;
    wire N__32237;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32229;
    wire N__32228;
    wire N__32225;
    wire N__32224;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32206;
    wire N__32203;
    wire N__32202;
    wire N__32201;
    wire N__32200;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32186;
    wire N__32185;
    wire N__32182;
    wire N__32179;
    wire N__32178;
    wire N__32175;
    wire N__32174;
    wire N__32173;
    wire N__32170;
    wire N__32163;
    wire N__32162;
    wire N__32161;
    wire N__32156;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32133;
    wire N__32130;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32110;
    wire N__32107;
    wire N__32106;
    wire N__32103;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32091;
    wire N__32086;
    wire N__32083;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32055;
    wire N__32050;
    wire N__32045;
    wire N__32044;
    wire N__32043;
    wire N__32042;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32026;
    wire N__32023;
    wire N__32014;
    wire N__32011;
    wire N__32004;
    wire N__31997;
    wire N__31994;
    wire N__31987;
    wire N__31982;
    wire N__31977;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31924;
    wire N__31923;
    wire N__31922;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31911;
    wire N__31908;
    wire N__31903;
    wire N__31902;
    wire N__31901;
    wire N__31898;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31863;
    wire N__31858;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31840;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31834;
    wire N__31833;
    wire N__31830;
    wire N__31829;
    wire N__31828;
    wire N__31825;
    wire N__31824;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31793;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31760;
    wire N__31755;
    wire N__31752;
    wire N__31741;
    wire N__31740;
    wire N__31739;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31731;
    wire N__31726;
    wire N__31723;
    wire N__31722;
    wire N__31721;
    wire N__31720;
    wire N__31719;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31666;
    wire N__31665;
    wire N__31664;
    wire N__31661;
    wire N__31656;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31648;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31633;
    wire N__31632;
    wire N__31631;
    wire N__31630;
    wire N__31627;
    wire N__31622;
    wire N__31619;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31564;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31399;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31135;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31086;
    wire N__31085;
    wire N__31084;
    wire N__31081;
    wire N__31072;
    wire N__31069;
    wire N__31068;
    wire N__31067;
    wire N__31066;
    wire N__31063;
    wire N__31062;
    wire N__31061;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31033;
    wire N__31028;
    wire N__31025;
    wire N__31012;
    wire N__31011;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30979;
    wire N__30978;
    wire N__30977;
    wire N__30976;
    wire N__30975;
    wire N__30974;
    wire N__30973;
    wire N__30972;
    wire N__30971;
    wire N__30970;
    wire N__30965;
    wire N__30958;
    wire N__30947;
    wire N__30944;
    wire N__30937;
    wire N__30936;
    wire N__30931;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30927;
    wire N__30926;
    wire N__30925;
    wire N__30924;
    wire N__30921;
    wire N__30916;
    wire N__30915;
    wire N__30914;
    wire N__30913;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30890;
    wire N__30889;
    wire N__30888;
    wire N__30887;
    wire N__30886;
    wire N__30885;
    wire N__30880;
    wire N__30875;
    wire N__30872;
    wire N__30867;
    wire N__30862;
    wire N__30857;
    wire N__30852;
    wire N__30845;
    wire N__30842;
    wire N__30833;
    wire N__30828;
    wire N__30817;
    wire N__30814;
    wire N__30813;
    wire N__30812;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30774;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30741;
    wire N__30740;
    wire N__30737;
    wire N__30732;
    wire N__30727;
    wire N__30724;
    wire N__30723;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30715;
    wire N__30712;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30671;
    wire N__30664;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30625;
    wire N__30622;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30614;
    wire N__30613;
    wire N__30610;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30567;
    wire N__30564;
    wire N__30563;
    wire N__30560;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30554;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30543;
    wire N__30542;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30515;
    wire N__30506;
    wire N__30503;
    wire N__30498;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30480;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30451;
    wire N__30448;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30434;
    wire N__30429;
    wire N__30426;
    wire N__30421;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30415;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30398;
    wire N__30397;
    wire N__30396;
    wire N__30395;
    wire N__30394;
    wire N__30389;
    wire N__30388;
    wire N__30387;
    wire N__30386;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30364;
    wire N__30361;
    wire N__30360;
    wire N__30359;
    wire N__30356;
    wire N__30355;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30340;
    wire N__30337;
    wire N__30336;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30310;
    wire N__30309;
    wire N__30306;
    wire N__30305;
    wire N__30304;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30292;
    wire N__30285;
    wire N__30282;
    wire N__30281;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30269;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30240;
    wire N__30237;
    wire N__30230;
    wire N__30225;
    wire N__30220;
    wire N__30215;
    wire N__30210;
    wire N__30209;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30193;
    wire N__30190;
    wire N__30183;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30145;
    wire N__30138;
    wire N__30135;
    wire N__30118;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30090;
    wire N__30085;
    wire N__30084;
    wire N__30083;
    wire N__30082;
    wire N__30081;
    wire N__30080;
    wire N__30079;
    wire N__30074;
    wire N__30069;
    wire N__30068;
    wire N__30067;
    wire N__30066;
    wire N__30065;
    wire N__30064;
    wire N__30063;
    wire N__30062;
    wire N__30061;
    wire N__30060;
    wire N__30059;
    wire N__30058;
    wire N__30055;
    wire N__30054;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30048;
    wire N__30047;
    wire N__30046;
    wire N__30045;
    wire N__30044;
    wire N__30043;
    wire N__30042;
    wire N__30041;
    wire N__30040;
    wire N__30039;
    wire N__30038;
    wire N__30037;
    wire N__30036;
    wire N__30033;
    wire N__30028;
    wire N__30021;
    wire N__30012;
    wire N__30005;
    wire N__29998;
    wire N__29991;
    wire N__29990;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29986;
    wire N__29985;
    wire N__29982;
    wire N__29977;
    wire N__29976;
    wire N__29975;
    wire N__29974;
    wire N__29973;
    wire N__29972;
    wire N__29971;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29962;
    wire N__29953;
    wire N__29944;
    wire N__29935;
    wire N__29934;
    wire N__29933;
    wire N__29932;
    wire N__29931;
    wire N__29930;
    wire N__29929;
    wire N__29924;
    wire N__29921;
    wire N__29914;
    wire N__29911;
    wire N__29904;
    wire N__29903;
    wire N__29900;
    wire N__29895;
    wire N__29888;
    wire N__29887;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29876;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29860;
    wire N__29859;
    wire N__29856;
    wire N__29845;
    wire N__29844;
    wire N__29843;
    wire N__29842;
    wire N__29839;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29811;
    wire N__29806;
    wire N__29797;
    wire N__29792;
    wire N__29789;
    wire N__29784;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29763;
    wire N__29756;
    wire N__29747;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29671;
    wire N__29670;
    wire N__29669;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29517;
    wire N__29516;
    wire N__29515;
    wire N__29514;
    wire N__29509;
    wire N__29508;
    wire N__29507;
    wire N__29504;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29489;
    wire N__29488;
    wire N__29487;
    wire N__29486;
    wire N__29483;
    wire N__29482;
    wire N__29481;
    wire N__29476;
    wire N__29471;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29451;
    wire N__29440;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29407;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29364;
    wire N__29361;
    wire N__29360;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29339;
    wire N__29332;
    wire N__29331;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29289;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29274;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29227;
    wire N__29226;
    wire N__29221;
    wire N__29220;
    wire N__29219;
    wire N__29216;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29208;
    wire N__29207;
    wire N__29206;
    wire N__29203;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29161;
    wire N__29160;
    wire N__29157;
    wire N__29156;
    wire N__29151;
    wire N__29146;
    wire N__29141;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29119;
    wire N__29112;
    wire N__29101;
    wire N__29100;
    wire N__29097;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29081;
    wire N__29080;
    wire N__29079;
    wire N__29078;
    wire N__29077;
    wire N__29076;
    wire N__29073;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29048;
    wire N__29045;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29026;
    wire N__29021;
    wire N__29014;
    wire N__29013;
    wire N__29010;
    wire N__29009;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28978;
    wire N__28971;
    wire N__28968;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28935;
    wire N__28930;
    wire N__28925;
    wire N__28918;
    wire N__28917;
    wire N__28916;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28893;
    wire N__28892;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28869;
    wire N__28868;
    wire N__28865;
    wire N__28860;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28839;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28791;
    wire N__28790;
    wire N__28789;
    wire N__28788;
    wire N__28785;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28781;
    wire N__28772;
    wire N__28769;
    wire N__28760;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28705;
    wire N__28702;
    wire N__28701;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28663;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28536;
    wire N__28535;
    wire N__28528;
    wire N__28525;
    wire N__28524;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28446;
    wire N__28443;
    wire N__28442;
    wire N__28441;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28427;
    wire N__28424;
    wire N__28423;
    wire N__28420;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28402;
    wire N__28397;
    wire N__28392;
    wire N__28387;
    wire N__28384;
    wire N__28375;
    wire N__28374;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28311;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28295;
    wire N__28294;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28259;
    wire N__28246;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28191;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28153;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28123;
    wire N__28122;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28090;
    wire N__28089;
    wire N__28088;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28060;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28046;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28017;
    wire N__28016;
    wire N__28013;
    wire N__28008;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27937;
    wire N__27936;
    wire N__27933;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27882;
    wire N__27879;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27843;
    wire N__27842;
    wire N__27839;
    wire N__27834;
    wire N__27829;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27821;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27753;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27745;
    wire N__27742;
    wire N__27741;
    wire N__27740;
    wire N__27735;
    wire N__27734;
    wire N__27729;
    wire N__27724;
    wire N__27721;
    wire N__27720;
    wire N__27717;
    wire N__27710;
    wire N__27707;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27681;
    wire N__27680;
    wire N__27677;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27567;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27342;
    wire N__27341;
    wire N__27338;
    wire N__27333;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27280;
    wire N__27279;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27142;
    wire N__27139;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27127;
    wire N__27124;
    wire N__27123;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27075;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27055;
    wire N__27052;
    wire N__27051;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26976;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26937;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26878;
    wire N__26875;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26860;
    wire N__26859;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26853;
    wire N__26852;
    wire N__26851;
    wire N__26850;
    wire N__26847;
    wire N__26846;
    wire N__26845;
    wire N__26844;
    wire N__26841;
    wire N__26834;
    wire N__26833;
    wire N__26832;
    wire N__26829;
    wire N__26828;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26816;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26799;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26783;
    wire N__26780;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26762;
    wire N__26757;
    wire N__26752;
    wire N__26747;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26724;
    wire N__26719;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26688;
    wire N__26683;
    wire N__26680;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26632;
    wire N__26629;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26614;
    wire N__26611;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26599;
    wire N__26598;
    wire N__26593;
    wire N__26590;
    wire N__26589;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26557;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26545;
    wire N__26544;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26532;
    wire N__26531;
    wire N__26528;
    wire N__26523;
    wire N__26518;
    wire N__26515;
    wire N__26514;
    wire N__26513;
    wire N__26512;
    wire N__26509;
    wire N__26508;
    wire N__26505;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26466;
    wire N__26463;
    wire N__26458;
    wire N__26449;
    wire N__26448;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26436;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26395;
    wire N__26390;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26305;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26280;
    wire N__26279;
    wire N__26278;
    wire N__26277;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26242;
    wire N__26241;
    wire N__26232;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26212;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26198;
    wire N__26193;
    wire N__26190;
    wire N__26185;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26176;
    wire N__26173;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26149;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26119;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26083;
    wire N__26080;
    wire N__26079;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26050;
    wire N__26049;
    wire N__26046;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26029;
    wire N__26026;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__25998;
    wire N__25993;
    wire N__25990;
    wire N__25989;
    wire N__25988;
    wire N__25987;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25976;
    wire N__25973;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25927;
    wire N__25926;
    wire N__25923;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25891;
    wire N__25888;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25844;
    wire N__25839;
    wire N__25836;
    wire N__25831;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25798;
    wire N__25797;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25776;
    wire N__25773;
    wire N__25768;
    wire N__25765;
    wire N__25764;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25706;
    wire N__25701;
    wire N__25698;
    wire N__25693;
    wire N__25692;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25684;
    wire N__25683;
    wire N__25682;
    wire N__25681;
    wire N__25680;
    wire N__25679;
    wire N__25678;
    wire N__25665;
    wire N__25664;
    wire N__25663;
    wire N__25662;
    wire N__25657;
    wire N__25652;
    wire N__25651;
    wire N__25650;
    wire N__25649;
    wire N__25648;
    wire N__25647;
    wire N__25644;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25620;
    wire N__25615;
    wire N__25610;
    wire N__25603;
    wire N__25602;
    wire N__25601;
    wire N__25600;
    wire N__25599;
    wire N__25598;
    wire N__25597;
    wire N__25596;
    wire N__25591;
    wire N__25586;
    wire N__25581;
    wire N__25580;
    wire N__25579;
    wire N__25578;
    wire N__25577;
    wire N__25576;
    wire N__25575;
    wire N__25572;
    wire N__25571;
    wire N__25570;
    wire N__25569;
    wire N__25566;
    wire N__25565;
    wire N__25564;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25541;
    wire N__25538;
    wire N__25531;
    wire N__25522;
    wire N__25519;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25479;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25453;
    wire N__25452;
    wire N__25449;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25431;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25412;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25365;
    wire N__25360;
    wire N__25357;
    wire N__25356;
    wire N__25353;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25329;
    wire N__25326;
    wire N__25321;
    wire N__25318;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25288;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25257;
    wire N__25254;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25236;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25171;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25138;
    wire N__25137;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25102;
    wire N__25101;
    wire N__25100;
    wire N__25099;
    wire N__25098;
    wire N__25097;
    wire N__25096;
    wire N__25093;
    wire N__25080;
    wire N__25079;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25075;
    wire N__25074;
    wire N__25073;
    wire N__25068;
    wire N__25067;
    wire N__25066;
    wire N__25061;
    wire N__25052;
    wire N__25051;
    wire N__25048;
    wire N__25047;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25032;
    wire N__25023;
    wire N__25012;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25004;
    wire N__25003;
    wire N__25002;
    wire N__25001;
    wire N__25000;
    wire N__24999;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24984;
    wire N__24975;
    wire N__24972;
    wire N__24961;
    wire N__24958;
    wire N__24957;
    wire N__24954;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24925;
    wire N__24924;
    wire N__24923;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24908;
    wire N__24907;
    wire N__24906;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24882;
    wire N__24879;
    wire N__24874;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24816;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24799;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24780;
    wire N__24777;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24735;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24717;
    wire N__24712;
    wire N__24711;
    wire N__24710;
    wire N__24707;
    wire N__24706;
    wire N__24705;
    wire N__24702;
    wire N__24701;
    wire N__24700;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24688;
    wire N__24685;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24664;
    wire N__24655;
    wire N__24654;
    wire N__24653;
    wire N__24650;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24642;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24631;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24582;
    wire N__24581;
    wire N__24578;
    wire N__24573;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24547;
    wire N__24544;
    wire N__24543;
    wire N__24540;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24393;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24337;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24329;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24264;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24249;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24205;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24183;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24128;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24106;
    wire N__24103;
    wire N__24102;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24079;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24057;
    wire N__24054;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24036;
    wire N__24033;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23965;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23917;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23775;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23757;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23745;
    wire N__23742;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23715;
    wire N__23710;
    wire N__23707;
    wire N__23706;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23679;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23658;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23622;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23595;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23548;
    wire N__23547;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23467;
    wire N__23464;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23406;
    wire N__23405;
    wire N__23404;
    wire N__23401;
    wire N__23394;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23379;
    wire N__23378;
    wire N__23375;
    wire N__23370;
    wire N__23367;
    wire N__23362;
    wire N__23361;
    wire N__23358;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23283;
    wire N__23282;
    wire N__23279;
    wire N__23274;
    wire N__23271;
    wire N__23266;
    wire N__23263;
    wire N__23262;
    wire N__23257;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23225;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23207;
    wire N__23202;
    wire N__23197;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23163;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23106;
    wire N__23103;
    wire N__23102;
    wire N__23101;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23063;
    wire N__23060;
    wire N__23053;
    wire N__23050;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23038;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22935;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22914;
    wire N__22909;
    wire N__22906;
    wire N__22905;
    wire N__22904;
    wire N__22901;
    wire N__22896;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22872;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22846;
    wire N__22843;
    wire N__22842;
    wire N__22841;
    wire N__22838;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22815;
    wire N__22814;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22680;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22614;
    wire N__22611;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22572;
    wire N__22569;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22534;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22526;
    wire N__22521;
    wire N__22516;
    wire N__22513;
    wire N__22512;
    wire N__22511;
    wire N__22508;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22482;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22424;
    wire N__22419;
    wire N__22416;
    wire N__22411;
    wire N__22408;
    wire N__22407;
    wire N__22406;
    wire N__22403;
    wire N__22398;
    wire N__22393;
    wire N__22390;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22366;
    wire N__22363;
    wire N__22362;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22250;
    wire N__22245;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22227;
    wire N__22226;
    wire N__22225;
    wire N__22224;
    wire N__22221;
    wire N__22212;
    wire N__22207;
    wire N__22206;
    wire N__22205;
    wire N__22202;
    wire N__22197;
    wire N__22194;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22158;
    wire N__22157;
    wire N__22154;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22122;
    wire N__22117;
    wire N__22114;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22092;
    wire N__22091;
    wire N__22088;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22041;
    wire N__22036;
    wire N__22033;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21999;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21976;
    wire N__21971;
    wire N__21970;
    wire N__21969;
    wire N__21968;
    wire N__21965;
    wire N__21964;
    wire N__21963;
    wire N__21960;
    wire N__21947;
    wire N__21944;
    wire N__21943;
    wire N__21936;
    wire N__21935;
    wire N__21934;
    wire N__21929;
    wire N__21926;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21907;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21873;
    wire N__21872;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21860;
    wire N__21857;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21763;
    wire N__21760;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21745;
    wire N__21742;
    wire N__21741;
    wire N__21736;
    wire N__21735;
    wire N__21734;
    wire N__21731;
    wire N__21726;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21691;
    wire N__21688;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21673;
    wire N__21672;
    wire N__21669;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21549;
    wire N__21548;
    wire N__21543;
    wire N__21540;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21243;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21228;
    wire N__21225;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21198;
    wire N__21195;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21166;
    wire N__21163;
    wire N__21162;
    wire N__21161;
    wire N__21154;
    wire N__21151;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21143;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21093;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21064;
    wire N__21063;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21017;
    wire N__21010;
    wire N__21009;
    wire N__21008;
    wire N__21003;
    wire N__21002;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20990;
    wire N__20983;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20971;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20959;
    wire N__20956;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20944;
    wire N__20941;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20911;
    wire N__20908;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20896;
    wire N__20893;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20885;
    wire N__20882;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20866;
    wire N__20865;
    wire N__20860;
    wire N__20857;
    wire N__20856;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20839;
    wire N__20838;
    wire N__20833;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20821;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20773;
    wire N__20770;
    wire N__20769;
    wire N__20768;
    wire N__20765;
    wire N__20760;
    wire N__20757;
    wire N__20752;
    wire N__20749;
    wire N__20748;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20730;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20707;
    wire N__20704;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20692;
    wire N__20689;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20681;
    wire N__20676;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20664;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20640;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20580;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20568;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20556;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20410;
    wire N__20407;
    wire N__20406;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20286;
    wire N__20285;
    wire N__20282;
    wire N__20277;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20247;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20232;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20220;
    wire N__20215;
    wire N__20212;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20167;
    wire N__20166;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20088;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20076;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20002;
    wire N__19999;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19978;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19944;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19929;
    wire N__19924;
    wire N__19921;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19909;
    wire N__19908;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19884;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19855;
    wire N__19854;
    wire N__19851;
    wire N__19850;
    wire N__19847;
    wire N__19842;
    wire N__19837;
    wire N__19834;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19819;
    wire N__19816;
    wire N__19815;
    wire N__19814;
    wire N__19813;
    wire N__19810;
    wire N__19803;
    wire N__19798;
    wire N__19797;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19785;
    wire N__19784;
    wire N__19783;
    wire N__19778;
    wire N__19773;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19759;
    wire N__19756;
    wire N__19755;
    wire N__19754;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19719;
    wire N__19714;
    wire N__19711;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19699;
    wire N__19698;
    wire N__19697;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19668;
    wire N__19665;
    wire N__19664;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19642;
    wire N__19641;
    wire N__19640;
    wire N__19639;
    wire N__19636;
    wire N__19631;
    wire N__19628;
    wire N__19621;
    wire N__19620;
    wire N__19615;
    wire N__19612;
    wire N__19611;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19572;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19280;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19212;
    wire N__19207;
    wire N__19204;
    wire N__19203;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19116;
    wire N__19115;
    wire N__19110;
    wire N__19107;
    wire N__19102;
    wire N__19099;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19056;
    wire N__19051;
    wire GNDG0;
    wire VCCG0;
    wire \ALU.N_675_0_0_cascade_ ;
    wire \ALU.N_703_0_0_0_cascade_ ;
    wire \ALU.N_681_0_0_0 ;
    wire \ALU.g0_0_2_cascade_ ;
    wire \ALU.N_699_0 ;
    wire \ALU.madd_167_cascade_ ;
    wire \ALU.madd_167 ;
    wire \ALU.g0_2 ;
    wire \ALU.a5_b_4_cascade_ ;
    wire \ALU.madd_139 ;
    wire \ALU.a2_b_8_cascade_ ;
    wire \ALU.madd_181_cascade_ ;
    wire \ALU.a3_b_8 ;
    wire \ALU.a3_b_8_cascade_ ;
    wire \ALU.madd_181 ;
    wire \ALU.madd_234_cascade_ ;
    wire \ALU.a7_b_8_cascade_ ;
    wire \ALU.madd_490_3 ;
    wire \ALU.madd_171_0_tz_cascade_ ;
    wire \ALU.madd_97 ;
    wire \ALU.madd_171_x_cascade_ ;
    wire \ALU.madd_171_0_tz ;
    wire \ALU.madd_171_cascade_ ;
    wire \ALU.madd_315_0_tz_cascade_ ;
    wire \ALU.madd_214 ;
    wire \ALU.madd_311_cascade_ ;
    wire \ALU.madd_268 ;
    wire \ALU.madd_268_cascade_ ;
    wire \ALU.madd_311 ;
    wire \ALU.madd_316 ;
    wire \ALU.a8_b_5 ;
    wire \ALU.a1_b_13_cascade_ ;
    wire \ALU.madd_388_cascade_ ;
    wire \ALU.madd_403_cascade_ ;
    wire \ALU.a1_b_13 ;
    wire \ALU.madd_403_0_cascade_ ;
    wire \ALU.a_6_ns_1_2_cascade_ ;
    wire TXbuffer_18_13_ns_1_2_cascade_;
    wire TXbuffer_18_6_ns_1_2_cascade_;
    wire TXbuffer_RNO_6Z0Z_2_cascade_;
    wire \ALU.madd_417 ;
    wire \ALU.madd_490_1_0_cascade_ ;
    wire \ALU.madd_378_0 ;
    wire \ALU.madd_388 ;
    wire \ALU.madd_402_cascade_ ;
    wire \ALU.madd_330 ;
    wire \ALU.madd_490_21 ;
    wire \ALU.madd_397 ;
    wire \ALU.a6_b_9_cascade_ ;
    wire \ALU.madd_490_10_cascade_ ;
    wire \ALU.madd_490_7_cascade_ ;
    wire \ALU.madd_490_11 ;
    wire \ALU.a2_b_13 ;
    wire TXbuffer_18_13_ns_1_0_cascade_;
    wire TXbuffer_RNO_5Z0Z_4_cascade_;
    wire TXbuffer_18_15_ns_1_4_cascade_;
    wire TXbuffer_RNO_1Z0Z_0;
    wire TXbuffer_18_15_ns_1_0_cascade_;
    wire TXbuffer_18_10_ns_1_3_cascade_;
    wire TXbuffer_RNO_0Z0Z_3_cascade_;
    wire TXbuffer_18_10_ns_1_4_cascade_;
    wire TXbuffer_RNO_0Z0Z_4;
    wire TXbuffer_RNO_1Z0Z_3;
    wire bfn_1_15_0_;
    wire clkdiv_cry_0;
    wire clkdiv_cry_1;
    wire clkdiv_cry_2;
    wire clkdiv_cry_3;
    wire clkdiv_cry_4;
    wire clkdiv_cry_5;
    wire clkdiv_cry_6;
    wire clkdiv_cry_7;
    wire clkdivZ0Z_8;
    wire bfn_1_16_0_;
    wire clkdivZ0Z_9;
    wire clkdiv_cry_8;
    wire clkdivZ0Z_10;
    wire clkdiv_cry_9;
    wire clkdivZ0Z_11;
    wire clkdiv_cry_10;
    wire clkdivZ0Z_12;
    wire clkdiv_cry_11;
    wire clkdivZ0Z_13;
    wire clkdiv_cry_12;
    wire clkdivZ0Z_14;
    wire clkdiv_cry_13;
    wire clkdivZ0Z_15;
    wire clkdiv_cry_14;
    wire clkdiv_cry_15;
    wire clkdivZ0Z_16;
    wire bfn_1_17_0_;
    wire clkdivZ0Z_17;
    wire clkdiv_cry_16;
    wire clkdivZ0Z_18;
    wire clkdiv_cry_17;
    wire clkdivZ0Z_19;
    wire clkdiv_cry_18;
    wire clkdivZ0Z_20;
    wire clkdiv_cry_19;
    wire clkdivZ0Z_21;
    wire clkdiv_cry_20;
    wire clkdivZ0Z_22;
    wire clkdiv_cry_21;
    wire clkdiv_cry_22;
    wire GPIO3_c;
    wire \ALU.madd_154_cascade_ ;
    wire \ALU.N_703_1_cascade_ ;
    wire \ALU.g0_cascade_ ;
    wire \ALU.madd_206 ;
    wire \ALU.madd_334_cascade_ ;
    wire \ALU.N_724_0_0_0 ;
    wire \ALU.madd_192_0 ;
    wire \ALU.madd_144 ;
    wire \ALU.g0_1 ;
    wire \ALU.N_695_0 ;
    wire \ALU.g0_4 ;
    wire \ALU.madd_197 ;
    wire \ALU.madd_112 ;
    wire \ALU.madd_191 ;
    wire \ALU.madd_234 ;
    wire \ALU.madd_112_cascade_ ;
    wire \ALU.madd_196_0 ;
    wire \ALU.madd_187 ;
    wire \ALU.madd_154 ;
    wire \ALU.madd_134 ;
    wire \ALU.g2_0_1 ;
    wire \ALU.madd_182_0 ;
    wire \ALU.a3_b_7 ;
    wire \ALU.a2_b_8 ;
    wire \ALU.madd_177 ;
    wire \ALU.madd_229 ;
    wire \ALU.madd_243_cascade_ ;
    wire \ALU.madd_219_0 ;
    wire \ALU.madd_181_0 ;
    wire \ALU.madd_315_0 ;
    wire \ALU.madd_320 ;
    wire \ALU.madd_393_cascade_ ;
    wire \ALU.madd_412 ;
    wire \ALU.madd_308_0_tz_0 ;
    wire \ALU.madd_299 ;
    wire \ALU.madd_209 ;
    wire \ALU.madd_243 ;
    wire \ALU.a0_b_13_cascade_ ;
    wire \ALU.madd_356 ;
    wire \ALU.madd_303_0 ;
    wire \ALU.madd_356_cascade_ ;
    wire \ALU.madd_175 ;
    wire \ALU.madd_388_0 ;
    wire \ALU.madd_393 ;
    wire \ALU.madd_340 ;
    wire \ALU.madd_355_cascade_ ;
    wire \ALU.madd_418 ;
    wire \ALU.madd_413_0 ;
    wire \ALU.madd_418_cascade_ ;
    wire \ALU.madd_293 ;
    wire \ALU.madd_336_0 ;
    wire \ALU.madd_351 ;
    wire \ALU.madd_346 ;
    wire \ALU.madd_172 ;
    wire \ALU.madd_346_cascade_ ;
    wire \ALU.madd_298_0 ;
    wire \ALU.madd_360 ;
    wire \ALU.madd_190 ;
    wire \ALU.madd_330_0_tz ;
    wire \ALU.madd_326 ;
    wire \ALU.madd_326_cascade_ ;
    wire \ALU.madd_350_0 ;
    wire \ALU.madd_355 ;
    wire \ALU.madd_408 ;
    wire \ALU.madd_350_0_cascade_ ;
    wire \ALU.madd_422 ;
    wire \ALU.a7_b_7_cascade_ ;
    wire \ALU.madd_383 ;
    wire \ALU.b_9_cascade_ ;
    wire \ALU.madd_326_0 ;
    wire \ALU.a5_b_9_cascade_ ;
    wire \ALU.a6_b_8 ;
    wire \ALU.a5_b_9 ;
    wire \ALU.a6_b_8_cascade_ ;
    wire \ALU.madd_378 ;
    wire \ALU.b_i_3_cascade_ ;
    wire \ALU.a3_b_11 ;
    wire \ALU.madd_382 ;
    wire \ALU.a4_b_10 ;
    wire \ALU.a11_b_3_cascade_ ;
    wire \ALU.madd_373 ;
    wire \ALU.a11_b_3 ;
    wire \ALU.madd_392 ;
    wire \ALU.madd_490_16 ;
    wire \ALU.madd_490_15_cascade_ ;
    wire \ALU.madd_490_19 ;
    wire \ALU.madd_339 ;
    wire \ALU.madd_340_0 ;
    wire \ALU.madd_490_1 ;
    wire \ALU.madd_490_9 ;
    wire \ALU.madd_490_0_cascade_ ;
    wire \ALU.madd_490_13 ;
    wire \ALU.madd_490_14 ;
    wire \ALU.r2_RNIFR6TZ0Z_15_cascade_ ;
    wire \ALU.b_15_cascade_ ;
    wire TXbuffer_18_13_ns_1_3;
    wire \ALU.r1_RNIAFSRZ0Z_15 ;
    wire \ALU.r5_RNIJBVTZ0Z_15_cascade_ ;
    wire \ALU.b_7_ns_1_15 ;
    wire \ALU.a_15_cascade_ ;
    wire \ALU.lshift_3_ns_1_15_cascade_ ;
    wire \ALU.b_6_ns_1_13_cascade_ ;
    wire \ALU.r6_RNIC9GA2Z0Z_13_cascade_ ;
    wire \ALU.b_13_cascade_ ;
    wire TXbuffer_18_13_ns_1_4_cascade_;
    wire TXbuffer_RNO_1Z0Z_4;
    wire \ALU.N_661_0 ;
    wire \ALU.madd_155_cascade_ ;
    wire \ALU.madd_109_0_tz_cascade_ ;
    wire \ALU.madd_109_cascade_ ;
    wire \ALU.N_687_0 ;
    wire \ALU.madd_159_N_2L1 ;
    wire \ALU.madd_159 ;
    wire \ALU.madd_150 ;
    wire \ALU.madd_155 ;
    wire \ALU.a7_b_1_cascade_ ;
    wire \ALU.a6_b_2 ;
    wire \ALU.a6_b_2_cascade_ ;
    wire \ALU.a7_b_1 ;
    wire \ALU.madd_99_cascade_ ;
    wire \ALU.madd_149 ;
    wire \ALU.madd_99 ;
    wire \ALU.madd_145 ;
    wire \ALU.madd_244 ;
    wire \ALU.madd_201 ;
    wire \ALU.madd_239 ;
    wire \ALU.a3_b_9_cascade_ ;
    wire \ALU.a3_b_9 ;
    wire \ALU.a4_b_8 ;
    wire \ALU.a4_b_8_cascade_ ;
    wire \ALU.madd_269 ;
    wire \ALU.madd_274 ;
    wire \ALU.madd_269_cascade_ ;
    wire \ALU.madd_289 ;
    wire \ALU.madd_185_1_cascade_ ;
    wire \ALU.madd_106 ;
    wire \ALU.g0_2_N_2L1_cascade_ ;
    wire \ALU.madd_186_0 ;
    wire \ALU.madd_228 ;
    wire \ALU.madd_338 ;
    wire \ALU.madd_337 ;
    wire \ALU.a0_b_13 ;
    wire \ALU.madd_335_0 ;
    wire \ALU.madd_233 ;
    wire \ALU.madd_238 ;
    wire \ALU.madd_294 ;
    wire \ALU.madd_304 ;
    wire \ALU.madd_253 ;
    wire \ALU.madd_341 ;
    wire \ALU.madd_336 ;
    wire \ALU.madd_335 ;
    wire \ALU.madd_283 ;
    wire \ALU.madd_124_0 ;
    wire \ALU.madd_218_0_tz ;
    wire \ALU.madd_218_cascade_ ;
    wire \ALU.madd_346_1 ;
    wire \ALU.a2_b_10 ;
    wire \ALU.a0_b_12_cascade_ ;
    wire \ALU.madd_279_0 ;
    wire \ALU.madd_331_0 ;
    wire \ALU.a0_b_12 ;
    wire \ALU.madd_218 ;
    wire \ALU.madd_202 ;
    wire \ALU.a12_b_0_cascade_ ;
    wire \ALU.madd_263 ;
    wire \ALU.madd_264_cascade_ ;
    wire \ALU.madd_288 ;
    wire \ALU.a12_b_0 ;
    wire \ALU.a10_b_2 ;
    wire \ALU.madd_259 ;
    wire \ALU.a7_b_5 ;
    wire \ALU.madd_259_cascade_ ;
    wire \ALU.madd_284_0 ;
    wire \ALU.b_3_ns_1_9_cascade_ ;
    wire \ALU.r4_RNIM58R1Z0Z_9 ;
    wire \ALU.b_3_ns_1_10_cascade_ ;
    wire \ALU.b_3_ns_1_11_cascade_ ;
    wire \ALU.r5_RNIQGFS1Z0Z_11_cascade_ ;
    wire \ALU.b_6_ns_1_10_cascade_ ;
    wire \ALU.b_6_ns_1_11_cascade_ ;
    wire \ALU.r6_RNI2H0U1Z0Z_11 ;
    wire \ALU.b_6_ns_1_9_cascade_ ;
    wire \ALU.r6_RNIUT042Z0Z_9 ;
    wire \ALU.r5_RNIH9VTZ0Z_14 ;
    wire \ALU.r1_RNI8DSRZ0Z_14_cascade_ ;
    wire \ALU.r2_RNIDP6TZ0Z_14 ;
    wire \ALU.b_7_ns_1_14_cascade_ ;
    wire \ALU.r6_RNILPNUZ0Z_14 ;
    wire \ALU.b_14_cascade_ ;
    wire bfn_3_11_0_;
    wire \ALU.r0_12_prm_8_11_s1_cy ;
    wire \ALU.r0_12_prm_7_11_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_11_s1 ;
    wire \ALU.r0_12_prm_7_11_s1 ;
    wire \ALU.r0_12_prm_5_11_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_11_s1 ;
    wire \ALU.r0_12_prm_5_11_s1 ;
    wire \ALU.r0_12_prm_4_11_s1 ;
    wire \ALU.r0_12_prm_3_11_s1 ;
    wire \ALU.r0_12_prm_2_11_s1 ;
    wire \ALU.r0_12_prm_1_11_s1_c_RNOZ0 ;
    wire bfn_3_12_0_;
    wire \ALU.r0_12_s1_11 ;
    wire \ALU.b_3_ns_1_12_cascade_ ;
    wire \ALU.b_6_ns_1_12_cascade_ ;
    wire \ALU.r6_RNI85GA2Z0Z_12 ;
    wire \ALU.r5_RNI05V82Z0Z_12 ;
    wire \ALU.r6_RNI85GA2Z0Z_12_cascade_ ;
    wire \ALU.b_3_ns_1_13_cascade_ ;
    wire \ALU.r5_RNI49V82Z0Z_13 ;
    wire \ALU.a_6_ns_1_15_cascade_ ;
    wire \ALU.r6_RNIH8772Z0Z_15 ;
    wire \ALU.r6_RNINRNUZ0Z_15 ;
    wire TXbuffer_18_6_ns_1_0_cascade_;
    wire TXbuffer_RNO_6Z0Z_0;
    wire TXbuffer_18_13_ns_1_7;
    wire bfn_3_15_0_;
    wire \ALU.r0_12_prm_8_11_s0_cy ;
    wire \ALU.r5_RNIE0AK8_0Z0Z_11 ;
    wire \ALU.r0_12_prm_8_11_s0 ;
    wire \ALU.r0_12_prm_7_11_s0 ;
    wire \ALU.r5_RNIE0AK8_1Z0Z_11 ;
    wire \ALU.r0_12_prm_6_11_s0 ;
    wire \ALU.a_i_11 ;
    wire \ALU.r0_12_prm_5_11_s0 ;
    wire \ALU.r0_12_prm_3_11_s0_sf ;
    wire \ALU.r0_12_prm_4_11_s0 ;
    wire \ALU.r0_12_prm_3_11_s0 ;
    wire \ALU.r0_12_prm_2_11_s0 ;
    wire bfn_3_16_0_;
    wire \ALU.r0_12_s0_11 ;
    wire \ALU.r0_12_s0_11_THRU_CO ;
    wire \ALU.g1_7_cascade_ ;
    wire \ALU.a4_b_0_0_5 ;
    wire \ALU.N_663_0_cascade_ ;
    wire \ALU.madd_109 ;
    wire \ALU.N_683_0_0_0 ;
    wire \ALU.madd_43_0_cascade_ ;
    wire \ALU.madd_77_0_tz ;
    wire \ALU.madd_278 ;
    wire \ALU.madd_273 ;
    wire \ALU.madd_345 ;
    wire \ALU.madd_159_N_3L3 ;
    wire \ALU.madd_61 ;
    wire \ALU.madd_140_0 ;
    wire \ALU.madd_140_0_cascade_ ;
    wire \ALU.madd_155_1 ;
    wire \ALU.madd_144_0_tz ;
    wire \ALU.a4_b_5 ;
    wire \ALU.g0_6_1 ;
    wire \ALU.r6_RNIUC0U1Z0Z_10 ;
    wire \ALU.r5_RNIMCFS1Z0Z_10 ;
    wire \ALU.a0_b_10 ;
    wire \ALU.a5_b_8_cascade_ ;
    wire \ALU.madd_325 ;
    wire \ALU.b_7_cascade_ ;
    wire \ALU.a5_b_7 ;
    wire \ALU.a5_b_5_cascade_ ;
    wire \ALU.madd_176 ;
    wire \ALU.a5_b_8 ;
    wire \ALU.a6_b_7 ;
    wire \ALU.madd_321 ;
    wire \ALU.b_6_ns_1_6_cascade_ ;
    wire \ALU.r6_RNIIH042Z0Z_6_cascade_ ;
    wire \ALU.b_6_cascade_ ;
    wire \ALU.g0_2_N_3L3 ;
    wire bZ0Z_2;
    wire \ALU.b_3_ns_1_6_cascade_ ;
    wire \ALU.r4_RNIAP7R1Z0Z_6 ;
    wire \ALU.a0_b_14 ;
    wire \ALU.g2_0 ;
    wire \ALU.g0_2_N_4L5 ;
    wire \ALU.madd_134_0_tz ;
    wire \ALU.madd_130_0 ;
    wire \ALU.madd_130 ;
    wire \ALU.madd_171_sx ;
    wire \ALU.madd_213 ;
    wire \ALU.a9_b_3 ;
    wire \ALU.madd_167_0 ;
    wire \ALU.b_6_ns_1_5_cascade_ ;
    wire \ALU.b_3_ns_1_5_cascade_ ;
    wire \ALU.r6_RNIBP2O1Z0Z_5 ;
    wire \ALU.r4_RNI0QNE1Z0Z_5_cascade_ ;
    wire \ALU.b_5_cascade_ ;
    wire TXbuffer_18_3_ns_1_1_cascade_;
    wire TXbuffer_RNO_5Z0Z_1_cascade_;
    wire r6_9;
    wire TXbuffer_18_6_ns_1_1_cascade_;
    wire TXbuffer_RNO_6Z0Z_1;
    wire r0_5;
    wire \ALU.a_3_ns_1_5_cascade_ ;
    wire r2_10;
    wire \ALU.a_6_ns_1_10_cascade_ ;
    wire \ALU.a_6_ns_1_11_cascade_ ;
    wire \ALU.r6_RNIT7372Z0Z_11_cascade_ ;
    wire \ALU.a_6_ns_1_7_cascade_ ;
    wire \ALU.b_6_ns_1_7_cascade_ ;
    wire \ALU.r6_RNIJ13O1Z0Z_7 ;
    wire r2_15;
    wire r2_7;
    wire TXbuffer_18_6_ns_1_7_cascade_;
    wire r3_10;
    wire r3_11;
    wire r3_15;
    wire r3_7;
    wire TXbuffer_18_13_ns_1_6_cascade_;
    wire TXbuffer_18_3_ns_1_2_cascade_;
    wire TXbuffer_RNO_5Z0Z_2;
    wire TXbuffer_18_3_ns_1_4;
    wire r6_10;
    wire r6_15;
    wire r7_10;
    wire r7_11;
    wire r7_15;
    wire TXbuffer_18_10_ns_1_6_cascade_;
    wire TXbuffer_RNO_1Z0Z_6;
    wire TXbuffer_RNO_0Z0Z_6_cascade_;
    wire TXbuffer_18_6_ns_1_6;
    wire TXbuffer_RNO_6Z0Z_6_cascade_;
    wire TXbuffer_18_15_ns_1_6;
    wire TXbuffer_18_3_ns_1_6_cascade_;
    wire TXbuffer_RNO_5Z0Z_6;
    wire \ALU.r0_12_prm_4_11_s1_c_RNOZ0 ;
    wire \ALU.r5_RNIAFVE5Z0Z_11 ;
    wire \ALU.r0_12_prm_5_11_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_11_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_11_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_11_s1_c_RNOZ0 ;
    wire TXbuffer_18_3_ns_1_5;
    wire \ALU.a4_b_4_cascade_ ;
    wire \ALU.madd_104 ;
    wire \ALU.madd_68_cascade_ ;
    wire \ALU.madd_82_0_cascade_ ;
    wire \ALU.madd_119 ;
    wire \ALU.a_6_cascade_ ;
    wire \ALU.g3 ;
    wire \ALU.madd_72_0_tz ;
    wire \ALU.madd_40_cascade_ ;
    wire \ALU.madd_72 ;
    wire \ALU.madd_95 ;
    wire \ALU.madd_72_cascade_ ;
    wire \ALU.madd_77 ;
    wire \ALU.b_8_cascade_ ;
    wire \ALU.madd_82 ;
    wire \ALU.madd_127_cascade_ ;
    wire \ALU.madd_223 ;
    wire \ALU.madd_223_0_tz ;
    wire \ALU.madd_105_0 ;
    wire \ALU.r4_RNIU5NK1Z0Z_8 ;
    wire \ALU.un9_addsub_axb_1_cascade_ ;
    wire \ALU.a7_b_3 ;
    wire \ALU.a_1_cascade_ ;
    wire \ALU.madd_228_0_tz ;
    wire \ALU.a_9_cascade_ ;
    wire \ALU.N_675_1 ;
    wire \ALU.bZ0Z_0_cascade_ ;
    wire \ALU.madd_130_0_0 ;
    wire \ALU.r6_RNIGC3D2Z0Z_7 ;
    wire \ALU.a_7_cascade_ ;
    wire \ALU.madd_76 ;
    wire \ALU.madd_213_0_tz ;
    wire \ALU.madd_209_0 ;
    wire \ALU.a8_b_4 ;
    wire \ALU.g0_7_x1_cascade_ ;
    wire \ALU.madd_76_1 ;
    wire \ALU.r6_RNIPK3D2Z0Z_9 ;
    wire \ALU.a9_b_4 ;
    wire \ALU.a_8_cascade_ ;
    wire \ALU.madd_224_0 ;
    wire \ALU.madd_224 ;
    wire \ALU.madd_121 ;
    wire \ALU.b_3_ns_1_8 ;
    wire r2_2;
    wire r3_2;
    wire \ALU.b_6_ns_1_2_cascade_ ;
    wire \ALU.b_6_ns_1_3_cascade_ ;
    wire r7_0;
    wire \ALU.b_6_ns_1_0_cascade_ ;
    wire r6_0;
    wire \ALU.a_3_ns_1_6_cascade_ ;
    wire r0_6;
    wire \ALU.a_6_ns_1_5_cascade_ ;
    wire r3_6;
    wire \ALU.a_6_ns_1_6_cascade_ ;
    wire \ALU.a_6_ns_1_9 ;
    wire \ALU.a_6_ns_1_8_cascade_ ;
    wire \ALU.r6_RNIKG3D2Z0Z_8 ;
    wire r2_8;
    wire r3_8;
    wire \ALU.b_6_ns_1_8_cascade_ ;
    wire \ALU.r6_RNIN53O1Z0Z_8 ;
    wire \ALU.a_6_ns_1_1_cascade_ ;
    wire \ALU.a_3_ns_1_10_cascade_ ;
    wire \ALU.r5_RNIVQN52Z0Z_10_cascade_ ;
    wire \ALU.a_3_ns_1_11_cascade_ ;
    wire \ALU.r5_RNI3VN52Z0Z_11 ;
    wire r3_3;
    wire \ALU.a_6_ns_1_3_cascade_ ;
    wire \ALU.a_3_ns_1_12_cascade_ ;
    wire r7_12;
    wire \ALU.a_6_ns_1_12_cascade_ ;
    wire \ALU.r6_RNI5S672Z0Z_12_cascade_ ;
    wire \ALU.r5_RNIS3672Z0Z_12 ;
    wire r2_5;
    wire r2_6;
    wire r2_9;
    wire bfn_5_13_0_;
    wire \ALU.r0_12_prm_8_15_s1_cy ;
    wire \ALU.r0_12_prm_7_15_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_15_s1 ;
    wire \ALU.r0_12_prm_6_15_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_15_s1 ;
    wire \ALU.r0_12_prm_6_15_s1 ;
    wire \ALU.r0_12_prm_4_15_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_15_s1 ;
    wire \ALU.r0_12_prm_4_15_s1 ;
    wire \ALU.r0_12_prm_3_15_s1 ;
    wire \ALU.r0_12_prm_2_15_s1 ;
    wire bfn_5_14_0_;
    wire \ALU.madd_axb_14 ;
    wire \ALU.r0_12_s1_15 ;
    wire \ALU.a_3_ns_1_13_cascade_ ;
    wire r2_13;
    wire \ALU.a_6_ns_1_13_cascade_ ;
    wire \ALU.r6_RNI90772Z0Z_13_cascade_ ;
    wire \ALU.r5_RNI10M52Z0Z_13 ;
    wire \ALU.r5_RNIPV8A9Z0Z_13_cascade_ ;
    wire r3_12;
    wire r3_5;
    wire r3_13;
    wire r6_13;
    wire TXbuffer_18_6_ns_1_5;
    wire r6_5;
    wire TXbuffer_RNO_5Z0Z_5;
    wire TXbuffer_RNO_6Z0Z_5_cascade_;
    wire r7_13;
    wire r7_5;
    wire TXbuffer_18_13_ns_1_5;
    wire TXbuffer_18_10_ns_1_5;
    wire \ALU.madd_68_0 ;
    wire \ALU.madd_46_0 ;
    wire \ALU.madd_100 ;
    wire \ALU.madd_105 ;
    wire \ALU.madd_46_0_cascade_ ;
    wire \ALU.madd_82_0 ;
    wire \ALU.a5_b_3 ;
    wire \ALU.g2_0_0_0 ;
    wire \ALU.a0_b_7 ;
    wire \ALU.a5_b_0 ;
    wire \ALU.madd_38_cascade_ ;
    wire \ALU.madd_87_cascade_ ;
    wire \ALU.madd_92_cascade_ ;
    wire \ALU.madd_78_0 ;
    wire \ALU.madd_68 ;
    wire \ALU.madd_78_0_cascade_ ;
    wire \ALU.madd_60 ;
    wire \ALU.madd_332_cascade_ ;
    wire \ALU.r6_RNIA0841Z0Z_0 ;
    wire \ALU.madd_92 ;
    wire \ALU.madd_120 ;
    wire \ALU.r6_RNII9FT1Z0Z_3 ;
    wire \ALU.b_3_cascade_ ;
    wire \ALU.un2_addsub_axb_3 ;
    wire \ALU.b_1_cascade_ ;
    wire \ALU.a4_b_1 ;
    wire \ALU.a_3_cascade_ ;
    wire \ALU.g1_1 ;
    wire \ALU.b_4_cascade_ ;
    wire \ALU.madd_214_0 ;
    wire \ALU.b_2_cascade_ ;
    wire \ALU.madd_134_0_tz_0 ;
    wire \ALU.madd_172_0 ;
    wire \ALU.madd_368 ;
    wire \ALU.a12_b_2 ;
    wire \ALU.a12_b_2_cascade_ ;
    wire \ALU.madd_372 ;
    wire \ALU.g1_2 ;
    wire \ALU.madd_311_0 ;
    wire b_1_repZ0Z1;
    wire b_1_repZ0Z2;
    wire r0_11;
    wire TXbuffer_18_3_ns_1_3_cascade_;
    wire TXbuffer_RNO_5Z0Z_3_cascade_;
    wire TXbuffer_18_15_ns_1_3;
    wire r2_11;
    wire r2_3;
    wire r6_11;
    wire TXbuffer_18_6_ns_1_3_cascade_;
    wire TXbuffer_RNO_6Z0Z_3;
    wire r4_11;
    wire bZ0Z_0;
    wire a_0_repZ0Z1;
    wire \ALU.a_6_ns_1_4_cascade_ ;
    wire r3_4;
    wire b_0_repZ0Z1;
    wire \ALU.b_6_ns_1_4_cascade_ ;
    wire \ALU.r6_RNI7L2O1Z0Z_4 ;
    wire \ALU.r6_RNI7L2O1Z0Z_4_cascade_ ;
    wire r2_12;
    wire r2_4;
    wire TXbuffer_18_6_ns_1_4_cascade_;
    wire r6_12;
    wire TXbuffer_RNO_6Z0Z_4;
    wire r1_11;
    wire r1_12;
    wire r1_13;
    wire r4_10;
    wire r4_12;
    wire r4_13;
    wire r4_5;
    wire r4_6;
    wire \ALU.a_3_ns_1_14_cascade_ ;
    wire r4_14;
    wire r2_14;
    wire r3_14;
    wire r7_14;
    wire \ALU.a_6_ns_1_14_cascade_ ;
    wire r6_14;
    wire \ALU.r6_RNID4772Z0Z_14_cascade_ ;
    wire \ALU.r5_RNI54M52Z0Z_14 ;
    wire r0_14;
    wire aZ0Z_0;
    wire aZ0Z_2;
    wire \ALU.a_3_ns_1_15_cascade_ ;
    wire \ALU.r5_RNI98M52Z0Z_15 ;
    wire \ALU.r0_12_11 ;
    wire r5_11;
    wire r5_12;
    wire r5_13;
    wire r5_14;
    wire \ALU.r0_12_15 ;
    wire r5_5;
    wire bfn_6_15_0_;
    wire \ALU.r0_12_prm_8_13_s0_cy ;
    wire \ALU.r0_12_prm_8_13_s0 ;
    wire \ALU.r0_12_prm_7_13_s0 ;
    wire \ALU.r0_12_prm_6_13_s0 ;
    wire \ALU.r0_12_prm_5_13_s0 ;
    wire \ALU.r0_12_prm_3_13_s0_sf ;
    wire \ALU.r0_12_prm_4_13_s0 ;
    wire \ALU.r0_12_prm_3_13_s0 ;
    wire \ALU.r0_12_prm_2_13_s0 ;
    wire bfn_6_16_0_;
    wire \ALU.r0_12_s0_13 ;
    wire \ALU.r0_12_13 ;
    wire r0_13;
    wire \ALU.r5_RNIK81F5Z0Z_13 ;
    wire \ALU.r0_12_prm_5_13_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_13_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_13_s0_c_RNOZ0 ;
    wire \ALU.madd_334 ;
    wire \ALU.madd_333 ;
    wire \ALU.madd_87 ;
    wire \ALU.madd_110 ;
    wire \ALU.madd_115 ;
    wire \ALU.madd_124 ;
    wire \ALU.madd_124_cascade_ ;
    wire \ALU.madd_160 ;
    wire \ALU.r6_RNIE0JB2Z0Z_6 ;
    wire \ALU.r4_RNI68Q22Z0Z_6 ;
    wire \ALU.a3_b_1 ;
    wire \ALU.a3_b_1_cascade_ ;
    wire \ALU.madd_18_cascade_ ;
    wire \ALU.madd_43_cascade_ ;
    wire \ALU.a2_b_3 ;
    wire \ALU.madd_332 ;
    wire \ALU.madd_94 ;
    wire \ALU.madd_33 ;
    wire \ALU.madd_38 ;
    wire \ALU.a0_b_6 ;
    wire \ALU.madd_51 ;
    wire \ALU.madd_51_cascade_ ;
    wire \ALU.madd_43 ;
    wire \ALU.madd_331 ;
    wire \ALU.a1_b_4 ;
    wire \ALU.madd_73_0_cascade_ ;
    wire \ALU.a1_b_5 ;
    wire \ALU.a2_b_4 ;
    wire \ALU.a1_b_5_cascade_ ;
    wire b_fastZ0Z_1;
    wire b_2_repZ0Z2;
    wire \ALU.r4_RNIMTDQZ0Z_1_cascade_ ;
    wire \ALU.b_7_ns_1_1 ;
    wire \ALU.madd_46 ;
    wire \ALU.a5_b_1 ;
    wire \ALU.a5_b_1_cascade_ ;
    wire \ALU.madd_50 ;
    wire \ALU.madd_55 ;
    wire \ALU.madd_50_cascade_ ;
    wire \ALU.madd_73 ;
    wire \ALU.madd_83 ;
    wire TXbuffer_RNO_1Z0Z_2;
    wire TXbuffer_18_15_ns_1_2;
    wire clkdivZ0Z_1;
    wire clkdivZ0Z_2;
    wire clkdivZ0Z_3;
    wire clkdivZ0Z_0;
    wire params5;
    wire \ALU.madd_axb_3_cascade_ ;
    wire \ALU.madd_14 ;
    wire \ALU.madd_cry_0_ma ;
    wire \ALU.madd_axb_0_l_ofx ;
    wire bfn_7_6_0_;
    wire \ALU.madd_cry_0 ;
    wire \ALU.madd_cry_1 ;
    wire \ALU.madd_cry_2 ;
    wire \ALU.madd_cry_3 ;
    wire \ALU.madd_axb_5_l_fx ;
    wire \ALU.madd_cry_4 ;
    wire \ALU.madd_axb_6_l_ofx ;
    wire \ALU.madd_cry_5 ;
    wire \ALU.madd_cry_6 ;
    wire \ALU.madd_cry_7 ;
    wire \ALU.madd_165 ;
    wire \ALU.madd_axb_8_l_fx ;
    wire bfn_7_7_0_;
    wire \ALU.madd_axb_9_l_ofx ;
    wire \ALU.madd_cry_9_ma ;
    wire \ALU.madd_cry_8 ;
    wire \ALU.madd_axb_10 ;
    wire \ALU.madd_cry_9_THRU_CO ;
    wire \ALU.madd_cry_9 ;
    wire \ALU.g0_13 ;
    wire \ALU.madd_axb_11_l_fx ;
    wire \ALU.madd_cry_10 ;
    wire \ALU.madd_cry_12_ma ;
    wire \ALU.madd_axb_12_l_ofx ;
    wire \ALU.mult_13 ;
    wire \ALU.madd_cry_11 ;
    wire \ALU.madd_axb_13_l_ofx ;
    wire \ALU.madd_cry_13_ma ;
    wire \ALU.madd_cry_12 ;
    wire \ALU.madd_cry_13 ;
    wire \ALU.madd_cry_13_THRU_CO ;
    wire \ALU.a13_b_1 ;
    wire \ALU.madd_373_0 ;
    wire \ALU.madd_368_0 ;
    wire \ALU.a9_b_5 ;
    wire \ALU.madd_398_0 ;
    wire \ALU.r4_RNIJJH11Z0Z_0 ;
    wire \ALU.r0_RNIBROOZ0Z_0_cascade_ ;
    wire a_fastZ0Z_1;
    wire \ALU.a_7_ns_1_0 ;
    wire r4_0;
    wire TXbuffer_18_3_ns_1_0_cascade_;
    wire TXbuffer_RNO_5Z0Z_0;
    wire TXbuffer_18_10_ns_1_0_cascade_;
    wire r5_0;
    wire TXbuffer_RNO_0Z0Z_0;
    wire r3_9;
    wire TXbuffer_18_13_ns_1_1;
    wire TXbuffer_18_10_ns_1_1_cascade_;
    wire TXbuffer_18_15_ns_1_1;
    wire TXbuffer_RNO_0Z0Z_1_cascade_;
    wire TXbuffer_RNO_1Z0Z_1;
    wire r1_10;
    wire r5_10;
    wire TXbuffer_18_10_ns_1_2_cascade_;
    wire TXbuffer_RNO_0Z0Z_2;
    wire r7_6;
    wire r7_7;
    wire r7_8;
    wire r7_9;
    wire r7_2;
    wire r7_3;
    wire r7_4;
    wire bfn_7_11_0_;
    wire \ALU.r0_12_prm_8_10_s0_cy ;
    wire \ALU.r0_12_prm_8_10_s0 ;
    wire \ALU.r0_12_prm_7_10_s0 ;
    wire \ALU.r0_12_prm_6_10_s0 ;
    wire \ALU.r0_12_prm_5_10_s0 ;
    wire \ALU.r0_12_prm_3_10_s0_sf ;
    wire \ALU.r0_12_prm_4_10_s0 ;
    wire \ALU.r0_12_prm_3_10_s0 ;
    wire \ALU.r0_12_prm_2_10_s0 ;
    wire bfn_7_12_0_;
    wire \ALU.mult_10 ;
    wire \ALU.r0_12_s0_10 ;
    wire \ALU.r0_12_10 ;
    wire r0_10;
    wire bfn_7_13_0_;
    wire \ALU.r0_12_prm_8_14_s0_cy ;
    wire \ALU.r0_12_prm_8_14_s0 ;
    wire \ALU.r0_12_prm_7_14_s0 ;
    wire \ALU.r0_12_prm_6_14_s0 ;
    wire \ALU.r0_12_prm_5_14_s0 ;
    wire \ALU.r0_12_prm_3_14_s0_sf ;
    wire \ALU.r0_12_prm_4_14_s0 ;
    wire \ALU.r0_12_prm_3_14_s0 ;
    wire \ALU.r0_12_prm_2_14_s0 ;
    wire bfn_7_14_0_;
    wire \ALU.mult_14 ;
    wire \ALU.r0_12_s0_14 ;
    wire \ALU.r0_12_14 ;
    wire r1_14;
    wire bfn_7_15_0_;
    wire \ALU.r0_12_prm_8_12_s0_cy ;
    wire \ALU.r0_12_prm_8_12_s0 ;
    wire \ALU.r0_12_prm_7_12_s0 ;
    wire \ALU.r0_12_prm_6_12_s0 ;
    wire \ALU.r0_12_prm_5_12_s0 ;
    wire \ALU.r0_12_prm_3_12_s0_sf ;
    wire \ALU.r0_12_prm_4_12_s0 ;
    wire \ALU.r0_12_prm_3_12_s0 ;
    wire \ALU.r0_12_prm_2_12_s0 ;
    wire bfn_7_16_0_;
    wire \ALU.mult_12 ;
    wire \ALU.r0_12_s0_12 ;
    wire \ALU.r0_12_12 ;
    wire r0_12;
    wire TXbuffer_RNO_1Z0Z_5;
    wire TXbuffer_RNO_0Z0Z_5;
    wire TXbuffer_18_15_ns_1_5;
    wire \ALU.a2_b_1_cascade_ ;
    wire \ALU.a1_b_2 ;
    wire \ALU.a2_b_1 ;
    wire \ALU.a1_b_2_cascade_ ;
    wire \ALU.madd_29_0 ;
    wire \ALU.madd_18 ;
    wire \ALU.madd_34 ;
    wire \ALU.madd_39_cascade_ ;
    wire \ALU.madd_39 ;
    wire \ALU.madd_23_cascade_ ;
    wire \ALU.madd_28 ;
    wire \ALU.madd_axb_4_l_fx ;
    wire \ALU.madd_8 ;
    wire \ALU.madd_19 ;
    wire \ALU.madd_66 ;
    wire a_1_repZ0Z1;
    wire \ALU.r6_RNIASIB2Z0Z_5 ;
    wire \ALU.r4_RNI24Q22Z0Z_5 ;
    wire \ALU.a0_b_4 ;
    wire \ALU.un2_addsub_axb_2 ;
    wire \ALU.madd_56 ;
    wire \ALU.madd_45 ;
    wire \ALU.madd_cry_6_ma ;
    wire r3_0;
    wire a_0_repZ0Z2;
    wire \ALU.r2_RNI18BOZ0Z_0 ;
    wire r2_0;
    wire r3_1;
    wire r2_1;
    wire \ALU.r2_RNI4H0SZ0Z_1 ;
    wire b_0_repZ0Z2;
    wire r7_1;
    wire r6_1;
    wire \ALU.r6_RNIC9P41Z0Z_1 ;
    wire \ALU.r6_RNIE5FT1Z0Z_2 ;
    wire \ALU.madd_13 ;
    wire \ALU.a2_b_0 ;
    wire \ALU.madd_3 ;
    wire \ALU.madd_4 ;
    wire \ALU.madd_3_cascade_ ;
    wire \ALU.a0_b_3 ;
    wire \ALU.a3_b_2 ;
    wire \ALU.rshift_3_ns_1_7_cascade_ ;
    wire \ALU.b_3_ns_1_7_cascade_ ;
    wire \ALU.r4_RNI82OE1Z0Z_7 ;
    wire r1_15;
    wire r5_15;
    wire TXbuffer_18_10_ns_1_7_cascade_;
    wire clkdivZ0Z_7;
    wire r0_15;
    wire clkdivZ0Z_6;
    wire TXbuffer_18_3_ns_1_7_cascade_;
    wire r4_15;
    wire clkdivZ0Z_5;
    wire TXbuffer_RNO_5Z0Z_7_cascade_;
    wire TXbuffer_RNO_6Z0Z_7;
    wire \ALU.a_3_ns_1_1_cascade_ ;
    wire r0_7;
    wire \ALU.a_3_ns_1_7_cascade_ ;
    wire \ALU.r4_RNI6BA92Z0Z_7 ;
    wire r1_8;
    wire \ALU.a_3_ns_1_8_cascade_ ;
    wire \ALU.r4_RNIAFA92Z0Z_8 ;
    wire \ALU.a_3_ns_1_3 ;
    wire \ALU.a_3_ns_1_2_cascade_ ;
    wire a_2_repZ0Z1;
    wire \ALU.a_3_ns_1_4_cascade_ ;
    wire a_fastZ0Z_2;
    wire r1_9;
    wire a_fastZ0Z_0;
    wire a_2_repZ0Z2;
    wire \ALU.a_3_ns_1_9_cascade_ ;
    wire \ALU.r4_RNIEJA92Z0Z_9 ;
    wire bfn_9_10_0_;
    wire \ALU.r0_12_prm_8_9_s0_cy ;
    wire \ALU.r0_12_prm_8_9_s0 ;
    wire \ALU.r0_12_prm_6_9_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_9_s0 ;
    wire \ALU.r0_12_prm_6_9_s0 ;
    wire \ALU.r0_12_prm_5_9_s0 ;
    wire \ALU.r0_12_prm_3_9_s0_sf ;
    wire \ALU.r0_12_prm_4_9_s0 ;
    wire \ALU.r0_12_prm_2_9_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_9_s0 ;
    wire \ALU.r0_12_prm_2_9_s0 ;
    wire bfn_9_11_0_;
    wire \ALU.mult_9 ;
    wire \ALU.r0_12_s0_9 ;
    wire r0_9;
    wire \ALU.r0_12_prm_8_11_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_12_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_2_15_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_2_13_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_1_14_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_15_s1_c_RNOZ0 ;
    wire \ALU.rshift_10_ns_1_3 ;
    wire \ALU.r5_RNI465TIZ0Z_13_cascade_ ;
    wire \ALU.r5_RNIOL1S71Z0Z_10 ;
    wire \ALU.r0_12_prm_5_12_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_11_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_12_s0_c_RNOZ0 ;
    wire bfn_9_15_0_;
    wire \ALU.r0_12_prm_8_13_s1_cy ;
    wire \ALU.r0_12_prm_7_13_s1_c_RNOZ0 ;
    wire \ALU.r5_RNID2JJ9_0Z0Z_13 ;
    wire \ALU.r0_12_prm_8_13_s1 ;
    wire \ALU.r0_12_prm_6_13_s1_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_13 ;
    wire \ALU.r0_12_prm_7_13_s1 ;
    wire \ALU.r0_12_prm_5_13_s1_c_RNOZ0 ;
    wire \ALU.r5_RNID2JJ9_1Z0Z_13 ;
    wire \ALU.r0_12_prm_6_13_s1 ;
    wire \ALU.r0_12_prm_4_13_s1_c_RNOZ0 ;
    wire \ALU.a_i_13 ;
    wire \ALU.r0_12_prm_5_13_s1 ;
    wire \ALU.r0_12_prm_4_13_s1 ;
    wire \ALU.r0_12_prm_3_13_s1 ;
    wire \ALU.r0_12_prm_2_13_s1 ;
    wire bfn_9_16_0_;
    wire \ALU.r0_12_s1_13 ;
    wire \ALU.r0_12_s1_13_THRU_CO ;
    wire \ALU.r0_12_prm_1_13_s1_c_RNOZ0 ;
    wire \ALU.rshift_3_ns_1_2_cascade_ ;
    wire \ALU.r6_RNIFJ8D2Z0Z_3 ;
    wire \ALU.r4_RNIMQ992Z0Z_3 ;
    wire \ALU.r4_RNIDI992Z0Z_1 ;
    wire \ALU.r6_RNI7B8D2Z0Z_1 ;
    wire \ALU.a1_b_3 ;
    wire \ALU.madd_135_0 ;
    wire \ALU.lshift_3_ns_1_6 ;
    wire \ALU.lshift_3_ns_1_7 ;
    wire \ALU.un9_addsub_axb_3 ;
    wire \ALU.madd_490_5 ;
    wire \ALU.rshift_3_ns_1_3_cascade_ ;
    wire \ALU.r0_12_prm_8_3_c_RNOZ0Z_3_cascade_ ;
    wire \ALU.r5_RNI67NNKZ0Z_10 ;
    wire bZ0Z_1;
    wire \ALU.r6_RNI6TET1Z0Z_0 ;
    wire \ALU.r4_RNIC5NE1Z0Z_0 ;
    wire \ALU.r6_RNIBF8D2Z0Z_2 ;
    wire \ALU.r4_RNIHM992Z0Z_2 ;
    wire \ALU.r6_RNI403D2Z0Z_4 ;
    wire \ALU.r4_RNIQU992Z0Z_4 ;
    wire aZ0Z_1;
    wire \ALU.un2_addsub_axb_4_cascade_ ;
    wire \ALU.rshift_10 ;
    wire \ALU.madd_76_0 ;
    wire \ALU.lshift_3_ns_1_11_cascade_ ;
    wire \ALU.un9_addsub_axb_4 ;
    wire \ALU.lshift_3_ns_1_9 ;
    wire r1_1;
    wire \ALU.r0_RNIE5LHZ0Z_1 ;
    wire \ALU.b_3_ns_1_0 ;
    wire r0_4;
    wire r1_4;
    wire \ALU.b_3_ns_1_4_cascade_ ;
    wire \ALU.r4_RNISLNE1Z0Z_4 ;
    wire r0_2;
    wire r1_2;
    wire \ALU.b_3_ns_1_2_cascade_ ;
    wire \ALU.r4_RNIKDNE1Z0Z_2 ;
    wire b_fastZ0Z_2;
    wire r1_3;
    wire b_fastZ0Z_0;
    wire b_2_repZ0Z1;
    wire r4_3;
    wire \ALU.b_3_ns_1_3_cascade_ ;
    wire \ALU.r4_RNIOHNE1Z0Z_3 ;
    wire r5_6;
    wire r5_7;
    wire r5_8;
    wire r5_9;
    wire r5_1;
    wire r5_2;
    wire r5_3;
    wire r5_4;
    wire bfn_10_9_0_;
    wire \ALU.r4_RNIUES39Z0Z_1 ;
    wire \ALU.un2_addsub_cry_0 ;
    wire \ALU.r4_RNIUM9JCZ0Z_2 ;
    wire \ALU.b_i_2 ;
    wire \ALU.un2_addsub_cry_1 ;
    wire \ALU.r4_RNINFAJCZ0Z_3 ;
    wire \ALU.b_i_3 ;
    wire \ALU.un2_addsub_cry_2 ;
    wire \ALU.r4_RNI20C8CZ0Z_4 ;
    wire \ALU.b_i_4 ;
    wire \ALU.un2_addsub_cry_3 ;
    wire \ALU.r4_RNI8B628_1Z0Z_5 ;
    wire \ALU.un2_addsub_cry_4 ;
    wire \ALU.r4_RNI2BKQ8_1Z0Z_6 ;
    wire \ALU.un2_addsub_cry_5 ;
    wire \ALU.un2_addsub_cry_6 ;
    wire \ALU.un2_addsub_cry_7 ;
    wire \ALU.r4_RNIKUMQ8_1Z0Z_8 ;
    wire bfn_10_10_0_;
    wire \ALU.un2_addsub_cry_8 ;
    wire \ALU.r5_RNIUF9K8_2Z0Z_10 ;
    wire \ALU.un2_addsub_cry_9 ;
    wire \ALU.r5_RNIE0AK8_2Z0Z_11 ;
    wire \ALU.un2_addsub_cry_10 ;
    wire \ALU.r5_RNISP2L9_2Z0Z_12 ;
    wire \ALU.un2_addsub_cry_11 ;
    wire \ALU.r5_RNID2JJ9_2Z0Z_13 ;
    wire \ALU.un2_addsub_cry_12 ;
    wire \ALU.r2_RNINPPC9_2Z0Z_14 ;
    wire \ALU.un2_addsub_cry_13 ;
    wire \ALU.un2_addsub_cry_14 ;
    wire r4_7;
    wire r4_8;
    wire \ALU.r0_12_9 ;
    wire r4_9;
    wire r4_1;
    wire r4_2;
    wire r4_4;
    wire \ALU.r5_RNIVF7TIZ0Z_13 ;
    wire \ALU.lshift_15_ns_1_15_cascade_ ;
    wire \ALU.r0_12_prm_8_11_s1_c_RNOZ0Z_1 ;
    wire \ALU.r0_12_prm_2_11_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_1_10_s0_c_RNOZ0 ;
    wire \ALU.N_884_i ;
    wire \ALU.r0_12_prm_8_12_s0_c_RNOZ0 ;
    wire \ALU.lshift_3_ns_1_3_cascade_ ;
    wire \ALU.r4_RNI1RK3KZ0Z_9 ;
    wire \ALU.r4_RNIOK1781Z0Z_9_cascade_ ;
    wire \ALU.lshift_11 ;
    wire \ALU.r5_RNI27VE5Z0Z_10 ;
    wire \ALU.un2_addsub_cry_12_c_RNI74A7EZ0 ;
    wire \ALU.r0_12_prm_2_13_s1_c_RNOZ0 ;
    wire \ALU.rshift_11 ;
    wire \ALU.r0_12_prm_8_10_s1_c_RNOZ0Z_1 ;
    wire bfn_10_15_0_;
    wire \ALU.r0_12_prm_8_10_s1_cy ;
    wire \ALU.r0_12_prm_7_10_s1_c_RNOZ0 ;
    wire \ALU.r5_RNIUF9K8_0Z0Z_10 ;
    wire \ALU.r0_12_prm_8_10_s1 ;
    wire \ALU.r0_12_prm_6_10_s1_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_10 ;
    wire \ALU.r0_12_prm_7_10_s1 ;
    wire \ALU.r0_12_prm_5_10_s1_c_RNOZ0 ;
    wire \ALU.r5_RNIUF9K8_1Z0Z_10 ;
    wire \ALU.r0_12_prm_6_10_s1 ;
    wire \ALU.r0_12_prm_4_10_s1_c_RNOZ0 ;
    wire \ALU.a_i_10 ;
    wire \ALU.r0_12_prm_5_10_s1 ;
    wire \ALU.r0_12_prm_4_10_s1 ;
    wire \ALU.r0_12_prm_2_10_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_10_s1 ;
    wire \ALU.r0_12_prm_2_10_s1 ;
    wire bfn_10_16_0_;
    wire \ALU.r0_12_s1_10 ;
    wire \ALU.r0_12_s1_10_THRU_CO ;
    wire \ALU.r0_12_prm_1_13_s0_c_RNOZ0 ;
    wire bfn_11_1_0_;
    wire \ALU.r0_12_prm_8_6_s1_c_THRU_CO ;
    wire \ALU.r0_12_prm_7_6_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_6_s1 ;
    wire \ALU.r0_12_prm_6_6_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_6_s1 ;
    wire \ALU.r0_12_prm_5_6_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_6_s1 ;
    wire \ALU.r0_12_prm_4_6_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_6_s1 ;
    wire \ALU.r0_12_prm_4_6_s1 ;
    wire \ALU.r0_12_prm_2_6_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_6_s1 ;
    wire \ALU.r0_12_prm_2_6_s1 ;
    wire bfn_11_2_0_;
    wire \ALU.r0_12_s1_6 ;
    wire \ALU.lshift_6_cascade_ ;
    wire \ALU.r0_12_prm_8_6_s1_c_RNOZ0 ;
    wire bfn_11_3_0_;
    wire \ALU.r0_12_prm_7_0_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_0_s0 ;
    wire \ALU.r0_12_prm_6_0_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_0_s0 ;
    wire \ALU.r0_12_prm_5_0_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_0_s0 ;
    wire \ALU.r2_RNIKG5N5Z0Z_0 ;
    wire \ALU.r0_12_prm_5_0_s0 ;
    wire \ALU.r0_12_prm_3_0_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_4_0_s0 ;
    wire \ALU.r0_12_prm_3_0_s0 ;
    wire \ALU.r0_12_prm_1_0_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_2_0_s0 ;
    wire \ALU.r0_12_s0_0 ;
    wire \ALU.rshift_0 ;
    wire bfn_11_4_0_;
    wire r1_0;
    wire \ALU.lshift_3_ns_1_8_cascade_ ;
    wire \ALU.r4_RNILIPV9Z0Z_6_cascade_ ;
    wire \ALU.r4_RNI1G9PKZ0Z_6_cascade_ ;
    wire r0_1;
    wire r0_3;
    wire \ALU.r0_12_0 ;
    wire r0_0;
    wire \ALU.r5_RNI9S2TIZ0Z_11_cascade_ ;
    wire \ALU.lshift_15_ns_1_13_cascade_ ;
    wire \ALU.un9_addsub_axb_2 ;
    wire \ALU.un14_log_0_i_11 ;
    wire \ALU.a6_b_0 ;
    wire bfn_11_8_0_;
    wire \ALU.r4_RNI90J9EZ0Z_1 ;
    wire \ALU.un9_addsub_cry_0 ;
    wire \ALU.r4_RNI468UDZ0Z_2 ;
    wire \ALU.un9_addsub_cry_1 ;
    wire \ALU.r4_RNIUU8UDZ0Z_3 ;
    wire \ALU.un9_addsub_cry_2 ;
    wire \ALU.r4_RNIQK1EDZ0Z_4 ;
    wire \ALU.un9_addsub_cry_3 ;
    wire \ALU.un9_addsub_cry_4 ;
    wire \ALU.un9_addsub_cry_5 ;
    wire \ALU.un9_addsub_cry_6 ;
    wire \ALU.un9_addsub_cry_7 ;
    wire bfn_11_9_0_;
    wire \ALU.un9_addsub_cry_8 ;
    wire \ALU.un9_addsub_cry_9 ;
    wire \ALU.b_11 ;
    wire \ALU.un9_addsub_cry_10 ;
    wire \ALU.un9_addsub_cry_11 ;
    wire \ALU.b_13 ;
    wire \ALU.un9_addsub_cry_12_c_RNISR30AZ0 ;
    wire \ALU.un9_addsub_cry_12 ;
    wire \ALU.un9_addsub_cry_13 ;
    wire \ALU.un9_addsub_cry_14 ;
    wire \ALU.r0_12_prm_6_10_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_13_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_2_12_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_1_9_s0_c_RNOZ0 ;
    wire \ALU.lshift_3_ns_1_13 ;
    wire \ALU.rshift_12 ;
    wire \ALU.un2_addsub_cry_9_c_RNIS67KDZ0 ;
    wire \ALU.r0_12_prm_2_10_s0_c_RNOZ0 ;
    wire \ALU.un2_addsub_cry_10_c_RNIS4T7DZ0 ;
    wire \ALU.r0_12_prm_2_11_s1_c_RNOZ0 ;
    wire \ALU.r5_RNIAP7U9Z0Z_10 ;
    wire \ALU.r5_RNIKU3HJZ0Z_10_cascade_ ;
    wire \ALU.r4_RNIQK1V71Z0Z_5_cascade_ ;
    wire \ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09 ;
    wire \ALU.r0_12_prm_1_11_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_2_14_s0_c_RNOZ0 ;
    wire \ALU.rshift_15 ;
    wire bfn_11_14_0_;
    wire \ALU.lshift_15 ;
    wire \ALU.r0_12_prm_8_15_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_15_s0_cy ;
    wire \ALU.r2_RNI7AQC9_0Z0Z_15 ;
    wire \ALU.r0_12_prm_8_15_s0 ;
    wire \ALU.r0_12_prm_6_15_s0_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_15 ;
    wire \ALU.r0_12_prm_7_15_s0 ;
    wire \ALU.r0_12_prm_5_15_s0_c_RNOZ0 ;
    wire \ALU.r2_RNI7AQC9_1Z0Z_15 ;
    wire \ALU.r0_12_prm_6_15_s0 ;
    wire \ALU.r5_RNI5P1F5Z0Z_15 ;
    wire \ALU.a_i_15 ;
    wire \ALU.r0_12_prm_5_15_s0 ;
    wire \ALU.r0_12_prm_3_15_s0_sf ;
    wire \ALU.r0_12_prm_4_15_s0 ;
    wire \ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9 ;
    wire \ALU.r0_12_prm_2_15_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_15_s0 ;
    wire \ALU.r0_12_prm_2_15_s0 ;
    wire \ALU.r0_12_prm_1_15_s0_c_RNOZ0 ;
    wire bfn_11_15_0_;
    wire \ALU.r0_12_s0_15 ;
    wire \ALU.r0_12_s0_15_THRU_CO ;
    wire \ALU.r5_RNIB8HG5Z0Z_12 ;
    wire \ALU.lshift_13 ;
    wire \ALU.r0_12_prm_8_13_s1_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8 ;
    wire \ALU.r0_12_prm_1_10_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_1_12_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_1_6_s1_c_RNOZ0 ;
    wire \ALU.rshift_3_ns_1_4_cascade_ ;
    wire bfn_12_2_0_;
    wire \ALU.r0_12_prm_7_0_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_0_s1 ;
    wire \ALU.r0_12_prm_6_0_s1_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_0 ;
    wire \ALU.r0_12_prm_7_0_s1 ;
    wire \ALU.r0_12_prm_5_0_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_0_s1 ;
    wire \ALU.r0_12_prm_4_0_s1_c_RNOZ0 ;
    wire \ALU.N_883_i ;
    wire \ALU.r0_12_prm_5_0_s1 ;
    wire \ALU.r0_12_prm_3_0_s1_c_RNOZ0 ;
    wire \ALU.mult_0 ;
    wire \ALU.r0_12_prm_4_0_s1 ;
    wire \ALU.r0_12_prm_3_0_s1 ;
    wire \ALU.r0_12_prm_1_0_s1_c_RNOZ0 ;
    wire \ALU.un9_addsub_axb_0 ;
    wire \ALU.r0_12_prm_2_0_s1 ;
    wire \ALU.r0_12_s1_0 ;
    wire bfn_12_3_0_;
    wire \ALU.r0_12_s1_0_THRU_CO ;
    wire \ALU.rshift_15_ns_1_0 ;
    wire \ALU.r0_12_prm_2_0_s0_c_RNOZ0 ;
    wire \ALU.rshift_15_ns_1_6 ;
    wire \ALU.rshift_3_ns_1_5 ;
    wire \ALU.r4_RNI9OH6AZ0Z_1_cascade_ ;
    wire \ALU.r5_RNIVQN52Z0Z_10 ;
    wire \ALU.r6_RNIP3372Z0Z_10 ;
    wire a_1_repZ0Z2;
    wire \ALU.a10_b_4 ;
    wire \ALU.lshift_3_ns_1_5 ;
    wire \ALU.lshift_15_ns_1_9 ;
    wire \ALU.r4_RNIF01FKZ0Z_2_cascade_ ;
    wire \ALU.r4_RNI2H9PKZ0Z_6 ;
    wire \ALU.lshift_9_cascade_ ;
    wire \ALU.r0_12_prm_8_9_s0_c_RNOZ0 ;
    wire bfn_12_6_0_;
    wire \ALU.r0_12_prm_8_7_s0_c_THRU_CO ;
    wire \ALU.r0_12_prm_8_7_s0 ;
    wire \ALU.r0_12_prm_6_7_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_7_s0 ;
    wire \ALU.r0_12_prm_6_7_s0 ;
    wire \ALU.r4_RNIFR136Z0Z_7 ;
    wire \ALU.r0_12_prm_5_7_s0 ;
    wire \ALU.r0_12_prm_3_7_s0_sf ;
    wire \ALU.r0_12_prm_4_7_s0 ;
    wire \ALU.r0_12_prm_3_7_s0 ;
    wire \ALU.r0_12_prm_2_7_s0 ;
    wire \ALU.r0_12_prm_1_7_s0_c_RNOZ0 ;
    wire bfn_12_7_0_;
    wire \ALU.mult_7 ;
    wire \ALU.r0_12_s0_7 ;
    wire r1_7;
    wire bfn_12_8_0_;
    wire \ALU.r0_12_prm_8_5_s0_cy ;
    wire \ALU.r0_12_prm_7_5_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_5_s0 ;
    wire \ALU.r0_12_prm_6_5_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_5_s0 ;
    wire \ALU.r0_12_prm_5_5_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_5_s0 ;
    wire \ALU.r4_RNIM8HG5Z0Z_5 ;
    wire \ALU.r0_12_prm_5_5_s0 ;
    wire \ALU.r0_12_prm_3_5_s0_sf ;
    wire \ALU.r0_12_prm_4_5_s0 ;
    wire \ALU.r0_12_prm_2_5_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_5_s0 ;
    wire \ALU.r0_12_prm_2_5_s0 ;
    wire bfn_12_9_0_;
    wire \ALU.mult_5 ;
    wire \ALU.r0_12_s0_5 ;
    wire \ALU.r0_12_5 ;
    wire r1_5;
    wire bfn_12_10_0_;
    wire \ALU.r0_12_prm_8_8_s0_cy ;
    wire \ALU.r0_12_prm_8_8_s0 ;
    wire \ALU.r0_12_prm_6_8_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_8_s0 ;
    wire \ALU.r0_12_prm_6_8_s0 ;
    wire \ALU.r0_12_prm_5_8_s0 ;
    wire \ALU.r0_12_prm_3_8_s0_sf ;
    wire \ALU.r0_12_prm_4_8_s0 ;
    wire \ALU.r0_12_prm_3_8_s0 ;
    wire \ALU.r0_12_prm_2_8_s0 ;
    wire bfn_12_11_0_;
    wire \ALU.r0_12_s0_8 ;
    wire \ALU.r0_12_prm_1_8_s0_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9 ;
    wire \ALU.r0_12_prm_1_15_s1_c_RNOZ0 ;
    wire \ALU.r4_RNIQK1V71Z0Z_5 ;
    wire bfn_12_13_0_;
    wire \ALU.r0_12_prm_8_12_s1_c_RNOZ0 ;
    wire \ALU.lshift_12 ;
    wire \ALU.r0_12_prm_8_12_s1_cy ;
    wire \ALU.r0_12_prm_7_12_s1_c_RNOZ0 ;
    wire \ALU.r5_RNISP2L9_0Z0Z_12 ;
    wire \ALU.r0_12_prm_8_12_s1 ;
    wire \ALU.un14_log_0_i_12 ;
    wire \ALU.r0_12_prm_7_12_s1 ;
    wire \ALU.r0_12_prm_5_12_s1_c_RNOZ0 ;
    wire \ALU.r5_RNISP2L9_1Z0Z_12 ;
    wire \ALU.r0_12_prm_6_12_s1 ;
    wire \ALU.r0_12_prm_4_12_s1_c_RNOZ0 ;
    wire \ALU.a_i_12 ;
    wire \ALU.r0_12_prm_5_12_s1 ;
    wire \ALU.r0_12_prm_4_12_s1 ;
    wire \ALU.un2_addsub_cry_11_c_RNICP8AEZ0 ;
    wire \ALU.r0_12_prm_2_12_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_12_s1 ;
    wire \ALU.r0_12_prm_2_12_s1 ;
    wire \ALU.r0_12_prm_1_12_s1_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_11_c_RNIAHI1AZ0 ;
    wire bfn_12_14_0_;
    wire \ALU.r0_12_s1_12 ;
    wire \ALU.r0_12_s1_12_THRU_CO ;
    wire \ALU.r0_12_prm_5_15_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_15_s1_c_RNOZ0Z_1 ;
    wire \ALU.r0_12_prm_8_0_s1_c_RNOZ0 ;
    wire \ALU.r5_RNIAV175Z0Z_15 ;
    wire \ALU.r0_12_prm_2_0_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_2_c_RNOZ0Z_3 ;
    wire \ALU.r4_RNI1G9PKZ0Z_6 ;
    wire \ALU.N_845_1 ;
    wire \ALU.rshift_15_ns_1_2_cascade_ ;
    wire \ALU.r5_RNI8R2TIZ0Z_11 ;
    wire \ALU.bZ0Z_0 ;
    wire \ALU.r4_RNID26E8_0Z0Z_0 ;
    wire \ALU.rshift_6 ;
    wire bfn_13_3_0_;
    wire \ALU.lshift_6 ;
    wire \ALU.r0_12_prm_8_6_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_6_s0_c_THRU_CO ;
    wire \ALU.r0_12_prm_8_6_s0 ;
    wire \ALU.un14_log_0_i_6 ;
    wire \ALU.r0_12_prm_7_6_s0 ;
    wire \ALU.r4_RNI2BKQ8_0Z0Z_6 ;
    wire \ALU.r0_12_prm_6_6_s0 ;
    wire \ALU.r4_RNIUGHG5Z0Z_6 ;
    wire \ALU.a_i_6 ;
    wire \ALU.r0_12_prm_5_6_s0 ;
    wire \ALU.r0_12_prm_3_6_s0_sf ;
    wire \ALU.r0_12_prm_4_6_s0 ;
    wire \ALU.un2_addsub_cry_5_c_RNIO30SDZ0 ;
    wire \ALU.r0_12_prm_2_6_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_6_s0 ;
    wire \ALU.r0_12_prm_2_6_s0 ;
    wire \ALU.un9_addsub_cry_5_c_RNI3CZ0Z019 ;
    wire \ALU.r0_12_prm_1_6_s0_c_RNOZ0 ;
    wire bfn_13_4_0_;
    wire \ALU.r0_12_s1_6_THRU_CO ;
    wire \ALU.mult_6 ;
    wire \ALU.r0_12_s0_6 ;
    wire r1_6;
    wire bfn_13_5_0_;
    wire \ALU.r0_12_prm_8_4_c_THRU_CO ;
    wire \ALU.a4_b_4 ;
    wire \ALU.r0_12_prm_7_4_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_4 ;
    wire \ALU.r0_12_prm_6_4_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_4 ;
    wire \ALU.r0_12_prm_7_4 ;
    wire \ALU.r0_12_prm_5_4_c_RNOZ0Z_0 ;
    wire \ALU.r0_12_prm_6_4 ;
    wire \ALU.a_i_4 ;
    wire \ALU.r0_12_prm_5_4 ;
    wire \ALU.mult_4 ;
    wire \ALU.r0_12_prm_4_4 ;
    wire \ALU.r0_12_prm_3_4 ;
    wire \ALU.r0_12_prm_2_4 ;
    wire bfn_13_6_0_;
    wire \ALU.r0_12_4 ;
    wire \ALU.r5_RNIKS4A9Z0Z_11 ;
    wire \ALU.r4_RNIVLAIAZ0Z_9 ;
    wire \ALU.r5_RNI0QK3KZ0Z_11_cascade_ ;
    wire \ALU.rshift_8 ;
    wire \ALU.un2_addsub_cry_3_c_RNI8MVBGZ0 ;
    wire \ALU.r0_12_prm_2_4_c_RNOZ0 ;
    wire \ALU.madd_axb_3 ;
    wire \ALU.madd_cry_2_THRU_CO ;
    wire \ALU.r0_12_prm_3_4_c_RNOZ0 ;
    wire \ALU.r0_12_prm_2_7_s0_c_RNOZ0 ;
    wire \ALU.r4_RNIODO6KZ0Z_5 ;
    wire \ALU.lshift_8_cascade_ ;
    wire \ALU.r0_12_prm_8_8_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_12_s1_c_RNOZ0Z_1 ;
    wire \ALU.r0_12_prm_7_8_s0_c_RNOZ0 ;
    wire \ALU.rshift_5 ;
    wire \ALU.r0_12_6 ;
    wire r6_6;
    wire \ALU.r0_12_7 ;
    wire r6_7;
    wire r6_8;
    wire r6_2;
    wire r6_3;
    wire \ALU.r0_12_4_THRU_CO ;
    wire r6_4;
    wire \ALU.r4_RNIN3236Z0Z_8 ;
    wire \ALU.rshift_3_ns_1_1 ;
    wire \ALU.r0_12_prm_8_1_c_RNOZ0Z_3_cascade_ ;
    wire \ALU.rshift_15_ns_1_1_cascade_ ;
    wire \ALU.r0_12_prm_8_8_s1_c_RNOZ0Z_1 ;
    wire bfn_13_10_0_;
    wire \ALU.lshift_8 ;
    wire \ALU.r0_12_prm_8_8_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_8_s1_cy ;
    wire \ALU.a8_b_8 ;
    wire \ALU.r0_12_prm_8_8_s1 ;
    wire \ALU.un14_log_0_i_8 ;
    wire \ALU.r0_12_prm_7_8_s1 ;
    wire \ALU.r0_12_prm_6_8_s1 ;
    wire \ALU.r0_12_prm_4_8_s1_c_RNOZ0 ;
    wire \ALU.a_i_8 ;
    wire \ALU.r0_12_prm_5_8_s1 ;
    wire \ALU.r0_12_prm_4_8_s1 ;
    wire \ALU.r0_12_prm_2_8_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_8_s1 ;
    wire \ALU.r0_12_prm_2_8_s1 ;
    wire \ALU.un9_addsub_cry_7_c_RNINZ0Z3519 ;
    wire \ALU.r0_12_prm_1_8_s1_c_RNOZ0 ;
    wire bfn_13_11_0_;
    wire \ALU.madd_cry_6_THRU_CO ;
    wire \ALU.madd_axb_7 ;
    wire \ALU.r0_12_s0_8_THRU_CO ;
    wire \ALU.r0_12_s1_8 ;
    wire \ALU.r0_12_8 ;
    wire r0_8;
    wire \ALU.un2_addsub_cry_7_c_RNI5ELEEZ0 ;
    wire \ALU.r0_12_prm_2_8_s0_c_RNOZ0 ;
    wire \ALU.r5_RNITTMB9Z0Z_12 ;
    wire \ALU.r5_RNITTMB9Z0Z_12_cascade_ ;
    wire \ALU.r5_RNITG1F5Z0Z_14 ;
    wire \ALU.r0_12_prm_5_14_s0_c_RNOZ0 ;
    wire \ALU.rshift_13 ;
    wire \ALU.r0_12_prm_6_14_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_14_s0_c_RNOZ0 ;
    wire \ALU.a_15 ;
    wire \ALU.b_15 ;
    wire \ALU.r0_12_prm_7_15_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_13_s1_c_RNOZ0Z_1 ;
    wire \ALU.b_12 ;
    wire \ALU.r0_12_prm_6_12_s1_c_RNOZ0 ;
    wire \ALU.r5_RNIPV8A9_0Z0Z_13 ;
    wire \ALU.rshift_2 ;
    wire bfn_14_1_0_;
    wire \ALU.r0_12_prm_8_2_c_THRU_CO ;
    wire \ALU.r0_12_prm_8_2 ;
    wire \ALU.r0_12_prm_7_2 ;
    wire \ALU.r0_12_prm_5_2_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_2 ;
    wire \ALU.r4_RNIL9636Z0Z_2 ;
    wire \ALU.a_i_2 ;
    wire \ALU.r0_12_prm_5_2 ;
    wire \ALU.r0_12_prm_4_2 ;
    wire \ALU.r0_12_prm_3_2 ;
    wire \ALU.r0_12_prm_2_2 ;
    wire bfn_14_2_0_;
    wire \ALU.r0_12_2 ;
    wire \ALU.r0_12_2_THRU_CO ;
    wire \ALU.lshift_2 ;
    wire \ALU.r0_12_prm_8_2_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_0_s0_c_RNOZ0 ;
    wire \ALU.a2_b_2 ;
    wire \ALU.r0_12_prm_7_2_c_RNOZ0 ;
    wire \ALU.lshift_0 ;
    wire \ALU.r4_RNIHENK8_1Z0Z_7 ;
    wire \ALU.b_i_0 ;
    wire \ALU.un2_addsub_axb_0_i ;
    wire \ALU.un2_addsub_cry_1_c_RNI1H7SGZ0 ;
    wire \ALU.r0_12_prm_2_2_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_2_c_RNOZ0 ;
    wire \ALU.b_4 ;
    wire \ALU.r0_12_prm_5_4_c_RNOZ0 ;
    wire \ALU.rshift_3_ns_1_9_cascade_ ;
    wire \ALU.a_11 ;
    wire \ALU.r0_12_prm_5_8_s0_c_RNOZ0 ;
    wire \ALU.N_610_1_cascade_ ;
    wire \ALU.r4_RNIVFRGQ_0Z0Z_2_cascade_ ;
    wire \ALU.lshift_4 ;
    wire \ALU.r0_12_prm_6_6_s0_c_RNOZ0 ;
    wire \ALU.a_13 ;
    wire \ALU.a_12 ;
    wire \ALU.r4_RNI9H7SJZ0Z_6 ;
    wire \ALU.r5_RNI0QK3KZ0Z_11 ;
    wire \ALU.r0_12_prm_8_4_c_RNOZ0Z_2_cascade_ ;
    wire \ALU.rshift_4 ;
    wire \ALU.lshift_15_ns_1_8 ;
    wire \ALU.lshift_3_ns_1_4 ;
    wire \ALU.r4_RNI6PL1LZ0Z_2 ;
    wire \ALU.r4_RNI6PL1LZ0Z_2_cascade_ ;
    wire \ALU.r4_RNIVFRGQZ0Z_2 ;
    wire \ALU.r4_RNIVFRGQ_0Z0Z_2 ;
    wire \ALU.r0_12_prm_8_4_c_RNOZ0 ;
    wire \ALU.r4_RNIODO6KZ0Z_7 ;
    wire \ALU.r0_12_prm_8_4_c_RNOZ0Z_3 ;
    wire \ALU.un9_addsub_cry_3_c_RNIV8DFIZ0 ;
    wire \ALU.r0_12_prm_1_4_c_RNOZ0 ;
    wire \ALU.r5_RNI7NOB9Z0Z_13 ;
    wire \ALU.r5_RNIUE7TIZ0Z_13 ;
    wire \ALU.r4_RNIRL1V71Z0Z_7 ;
    wire \ALU.a6_b_6 ;
    wire \ALU.r0_12_prm_7_6_s0_c_RNOZ0 ;
    wire \ALU.rshift_1 ;
    wire bfn_14_8_0_;
    wire \ALU.lshift_1 ;
    wire \ALU.r0_12_prm_8_1_c_THRU_CO ;
    wire \ALU.a1_b_1 ;
    wire \ALU.r0_12_prm_7_1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_1 ;
    wire \ALU.r0_12_prm_6_1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_1 ;
    wire \ALU.r0_12_prm_5_1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_1 ;
    wire \ALU.r4_RNID1636Z0Z_1 ;
    wire \ALU.a_i_1 ;
    wire \ALU.r0_12_prm_5_1 ;
    wire \ALU.r0_12_prm_3_1_c_RNOZ0 ;
    wire \ALU.mult_1 ;
    wire \ALU.r0_12_prm_4_1 ;
    wire \ALU.r0_12_prm_3_1 ;
    wire \ALU.r0_12_prm_2_1 ;
    wire bfn_14_9_0_;
    wire \ALU.r0_12_1 ;
    wire \ALU.r0_12_1_THRU_CO ;
    wire \ALU.un9_addsub_cry_0_c_RNIG8GLJZ0 ;
    wire \ALU.r0_12_prm_1_1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_9_s0_c_RNOZ0 ;
    wire \ALU.r4_RNIKUMQ8_0Z0Z_8 ;
    wire \ALU.r0_12_prm_6_8_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_10_s0_c_RNOZ0 ;
    wire \ALU.lshift_3_ns_1_10 ;
    wire \ALU.r4_RNI67NNKZ0Z_7_cascade_ ;
    wire \ALU.lshift_10 ;
    wire \ALU.N_610_1 ;
    wire \ALU.r4_RNIAHIIAZ0Z_2 ;
    wire \ALU.r4_RNI38O1GZ0Z_2 ;
    wire \ALU.r4_RNI38O1GZ0Z_2_cascade_ ;
    wire \ALU.r4_RNICN8R81Z0Z_7 ;
    wire \ALU.r0_12_prm_8_10_s1_c_RNOZ0 ;
    wire \ALU.r4_RNI67NNKZ0Z_7 ;
    wire \ALU.r5_RNI355TIZ0Z_13 ;
    wire \ALU.r4_RNIO7CSJZ0Z_4 ;
    wire \ALU.lshift_15_ns_1_14_cascade_ ;
    wire \ALU.r4_RNILVIQFZ0Z_2 ;
    wire \ALU.r0_12_prm_8_9_s1_c_RNOZ0Z_1 ;
    wire bfn_14_12_0_;
    wire \ALU.r0_12_prm_8_9_s1_c_RNOZ0 ;
    wire \ALU.lshift_9 ;
    wire \ALU.r0_12_prm_8_9_s1_cy ;
    wire \ALU.r0_12_prm_7_9_s1_c_RNOZ0 ;
    wire \ALU.r4_RNISU5D9_0Z0Z_9 ;
    wire \ALU.r0_12_prm_8_9_s1 ;
    wire \ALU.r0_12_prm_6_9_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_9_s1 ;
    wire \ALU.r4_RNISU5D9_1Z0Z_9 ;
    wire \ALU.r0_12_prm_5_9_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_9_s1 ;
    wire \ALU.a_i_9 ;
    wire \ALU.r0_12_prm_5_9_s1 ;
    wire \ALU.r0_12_prm_4_9_s1 ;
    wire \ALU.r0_12_prm_2_9_s1_c_RNOZ0 ;
    wire \ALU.un2_addsub_cry_8_c_RNINO51FZ0 ;
    wire \ALU.r0_12_prm_3_9_s1 ;
    wire \ALU.r0_12_prm_2_9_s1 ;
    wire \ALU.r0_12_prm_1_9_s1_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9 ;
    wire bfn_14_13_0_;
    wire \ALU.r0_12_s1_9 ;
    wire \ALU.r0_12_s1_9_THRU_CO ;
    wire \ALU.r0_12_prm_7_14_s0_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_2 ;
    wire \ALU.mult_2 ;
    wire \ALU.madd_cry_0_THRU_CO ;
    wire \ALU.madd_axb_1 ;
    wire \ALU.r0_12_prm_3_2_c_RNOZ0 ;
    wire \ALU.a_4 ;
    wire \ALU.r4_RNI87HO5Z0Z_4 ;
    wire \ALU.b_2 ;
    wire \ALU.r0_12_prm_5_2_c_RNOZ0Z_0 ;
    wire \ALU.un9_addsub_cry_1_c_RNIKO6AJZ0 ;
    wire \ALU.r0_12_prm_1_2_c_RNOZ0 ;
    wire \ALU.b_6 ;
    wire \ALU.a_6 ;
    wire \ALU.r0_12_prm_5_6_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_7_s0_c_RNOZ0 ;
    wire \ALU.r5_RNILM5AEZ0Z_15 ;
    wire \ALU.r5_RNILV3HJZ0Z_12 ;
    wire \ALU.rshift_9 ;
    wire \ALU.r4_RNI9H7SJZ0Z_5 ;
    wire \ALU.lshift_7_cascade_ ;
    wire \ALU.r0_12_prm_8_7_s0_c_RNOZ0 ;
    wire \ALU.rshift_7 ;
    wire bfn_15_4_0_;
    wire \ALU.r0_12_prm_8_7_s1_c_RNOZ0 ;
    wire \ALU.lshift_7 ;
    wire \ALU.r0_12_prm_8_7_s1_c_THRU_CO ;
    wire \ALU.r0_12_prm_8_7_s1 ;
    wire \ALU.un14_log_0_i_7 ;
    wire \ALU.r0_12_prm_7_7_s1 ;
    wire \ALU.r0_12_prm_5_7_s1_c_RNOZ0 ;
    wire \ALU.r4_RNIHENK8_0Z0Z_7 ;
    wire \ALU.r0_12_prm_6_7_s1 ;
    wire \ALU.r0_12_prm_4_7_s1_c_RNOZ0 ;
    wire \ALU.a_i_7 ;
    wire \ALU.r0_12_prm_5_7_s1 ;
    wire \ALU.r0_12_prm_4_7_s1 ;
    wire \ALU.un2_addsub_cry_6_c_RNIPJK8EZ0 ;
    wire \ALU.r0_12_prm_2_7_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_7_s1 ;
    wire \ALU.r0_12_prm_2_7_s1 ;
    wire bfn_15_5_0_;
    wire \ALU.r0_12_s1_7 ;
    wire \ALU.r0_12_s1_7_THRU_CO ;
    wire \ALU.r5_RNISMSV4Z0Z_15 ;
    wire \ALU.rshift_15_ns_1_3 ;
    wire \ALU.r5_RNI465TIZ0Z_13 ;
    wire \ALU.r4_RNIF01FKZ0Z_2 ;
    wire \ALU.b_7 ;
    wire \ALU.a_7 ;
    wire \ALU.r0_12_prm_6_7_s1_c_RNOZ0 ;
    wire \ALU.b_3 ;
    wire \ALU.r0_12_prm_1_5_s0_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_9 ;
    wire \ALU.a_5 ;
    wire \ALU.b_5 ;
    wire \ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8 ;
    wire \ALU.r0_12_prm_1_7_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_5_s1_c_RNOZ0Z_1 ;
    wire bfn_15_7_0_;
    wire \ALU.r0_12_prm_8_5_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_5_s1_cy ;
    wire \ALU.r0_12_prm_8_5_s1 ;
    wire \ALU.r0_12_prm_6_5_s1_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_5 ;
    wire \ALU.r0_12_prm_7_5_s1 ;
    wire \ALU.r4_RNI8B628_0Z0Z_5 ;
    wire \ALU.r0_12_prm_5_5_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_6_5_s1 ;
    wire \ALU.r0_12_prm_4_5_s1_c_RNOZ0 ;
    wire \ALU.a_i_5 ;
    wire \ALU.r0_12_prm_5_5_s1 ;
    wire \ALU.r0_12_prm_4_5_s1 ;
    wire \ALU.r0_12_prm_2_5_s1_c_RNOZ0 ;
    wire \ALU.un2_addsub_cry_4_c_RNILPG3DZ0 ;
    wire \ALU.r0_12_prm_3_5_s1 ;
    wire \ALU.r0_12_prm_2_5_s1 ;
    wire \ALU.r0_12_prm_1_5_s1_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88 ;
    wire bfn_15_8_0_;
    wire \ALU.r0_12_s1_5 ;
    wire \ALU.r0_12_s1_5_THRU_CO ;
    wire \ALU.r0_12_prm_5_8_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_10_s0_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_1_c_RNOZ0Z_0 ;
    wire \ALU.rshift_14 ;
    wire \ALU.N_622_1 ;
    wire \ALU.r0_12_prm_8_1_c_RNOZ0 ;
    wire \ALU.b_8 ;
    wire \ALU.a_8 ;
    wire \ALU.r0_12_prm_7_8_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_9_s0_c_RNOZ0 ;
    wire \ALU.un1_yindexZ0Z_1 ;
    wire \ALU.un1_yindexZ0Z_2 ;
    wire \ALU.un1_yindexZ0Z_3 ;
    wire \ALU.un1_yindexZ0Z_4 ;
    wire \ALU.un1_yindexZ0Z_5 ;
    wire \ALU.un1_yindexZ0Z_6 ;
    wire \ALU.un1_yindexZ0Z_7 ;
    wire \ALU.b_9 ;
    wire \ALU.r4_RNISU5D9_2Z0Z_9 ;
    wire \ALU.a5_b_5 ;
    wire \ALU.r0_12_prm_7_5_s1_c_RNOZ0 ;
    wire \ALU.b_14 ;
    wire \ALU.a_14 ;
    wire \ALU.r0_12_prm_7_7_s1_c_RNOZ0 ;
    wire \ALU.b_1 ;
    wire \ALU.un14_log_0_i_1 ;
    wire \ALU.a7_b_7 ;
    wire \ALU.r0_12_prm_7_7_s0_c_RNOZ0 ;
    wire bfn_15_13_0_;
    wire \ALU.r0_12_prm_8_14_s1_c_RNOZ0 ;
    wire \ALU.lshift_14 ;
    wire \ALU.r0_12_prm_8_14_s1_cy ;
    wire \ALU.r0_12_prm_7_14_s1_c_RNOZ0 ;
    wire \ALU.r2_RNINPPC9_0Z0Z_14 ;
    wire \ALU.r0_12_prm_8_14_s1 ;
    wire \ALU.r0_12_prm_6_14_s1_c_RNOZ0 ;
    wire \ALU.un14_log_0_i_14 ;
    wire \ALU.r0_12_prm_7_14_s1 ;
    wire \ALU.r0_12_prm_5_14_s1_c_RNOZ0 ;
    wire \ALU.r2_RNINPPC9_1Z0Z_14 ;
    wire \ALU.r0_12_prm_6_14_s1 ;
    wire \ALU.r0_12_prm_4_14_s1_c_RNOZ0 ;
    wire \ALU.a_i_14 ;
    wire \ALU.r0_12_prm_5_14_s1 ;
    wire \ALU.r0_12_prm_4_14_s1 ;
    wire \ALU.un2_addsub_cry_13_c_RNIR5I0EZ0 ;
    wire \ALU.r0_12_prm_2_14_s1_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_14_s1 ;
    wire \ALU.r0_12_prm_2_14_s1 ;
    wire \ALU.r0_12_prm_1_14_s1_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9 ;
    wire bfn_15_14_0_;
    wire \ALU.r0_12_s1_14 ;
    wire \ALU.r0_12_s1_14_THRU_CO ;
    wire \ALU.aZ0Z_0 ;
    wire \ALU.a_1 ;
    wire \ALU.a_2 ;
    wire \ALU.rshift_3_ns_1_0_cascade_ ;
    wire \ALU.r4_RNII2A0LZ0Z_2 ;
    wire \ALU.lshift_5 ;
    wire \ALU.r0_12_prm_8_5_s0_c_RNOZ0 ;
    wire \ALU.r4_RNI0C236Z0Z_9 ;
    wire \ALU.rshift_3 ;
    wire bfn_16_5_0_;
    wire \ALU.r0_12_prm_8_3_c_RNOZ0 ;
    wire \ALU.r0_12_prm_8_3_c_THRU_CO ;
    wire \ALU.r0_12_prm_7_3_c_RNOZ0 ;
    wire \ALU.a3_b_3 ;
    wire \ALU.r0_12_prm_8_3 ;
    wire \ALU.un14_log_0_i_3 ;
    wire \ALU.r0_12_prm_6_3_c_RNOZ0 ;
    wire \ALU.r0_12_prm_7_3 ;
    wire \ALU.r0_12_prm_5_3_c_RNOZ0 ;
    wire \ALU.r0_12_prm_5_3_c_RNOZ0Z_0 ;
    wire \ALU.r0_12_prm_6_3 ;
    wire \ALU.r4_RNIUH636Z0Z_3 ;
    wire \ALU.a_3 ;
    wire \ALU.a_i_3 ;
    wire \ALU.r0_12_prm_5_3 ;
    wire \ALU.r0_12_prm_4_3 ;
    wire \ALU.r0_12_prm_3_3 ;
    wire \ALU.r0_12_prm_2_3 ;
    wire \ALU.r0_12_prm_1_3_c_RNOZ0 ;
    wire \ALU.un9_addsub_cry_2_c_RNIOR8AJZ0 ;
    wire bfn_16_6_0_;
    wire \ALU.r0_12_3 ;
    wire \ALU.r0_12_3_THRU_CO ;
    wire \ALU.un2_addsub_cry_2_c_RNI3K9SGZ0 ;
    wire \ALU.r0_12_prm_2_3_c_RNOZ0 ;
    wire \ALU.r0_12_prm_3_3_c_RNOZ0 ;
    wire \ALU.madd_axb_2 ;
    wire \ALU.madd_cry_1_THRU_CO ;
    wire \ALU.mult_3 ;
    wire TXbuffer_RNO_1Z0Z_7;
    wire TXbuffer_RNO_0Z0Z_7;
    wire clkdivZ0Z_4;
    wire TXbuffer_18_15_ns_1_7;
    wire yZ0Z_2;
    wire \ALU.un1_yindexZ0Z_8 ;
    wire yZ0Z_0;
    wire yZ0Z_1;
    wire TXbufferZ0Z_7;
    wire \INVFTDI.TXshift_7C_net ;
    wire TXbufferZ0Z_1;
    wire TXbufferZ0Z_2;
    wire \FTDI.TXshiftZ0Z_2 ;
    wire \INVFTDI.TXshift_1C_net ;
    wire TXbufferZ0Z_4;
    wire \FTDI.TXshiftZ0Z_4 ;
    wire TXbufferZ0Z_3;
    wire \FTDI.TXshiftZ0Z_3 ;
    wire \FTDI.TXshiftZ0Z_7 ;
    wire TXbufferZ0Z_6;
    wire \FTDI.TXshiftZ0Z_6 ;
    wire TXbufferZ0Z_5;
    wire \FTDI.TXshiftZ0Z_5 ;
    wire \INVFTDI.TXshift_4C_net ;
    wire \ALU.b_10 ;
    wire \ALU.a_10 ;
    wire \ALU.r0_12_prm_7_10_s0_c_RNOZ0 ;
    wire paramsZ0Z_3;
    wire paramsZ0Z_2;
    wire \ALU.r4_RNII2A0LZ0Z_1 ;
    wire \ALU.lshift_3 ;
    wire \ALU.lshift63Z0Z_2 ;
    wire \ALU.r5_RNIAG9A9Z0Z_15 ;
    wire \ALU.r0_12_prm_8_14_s1_c_RNOZ0Z_1 ;
    wire op_i_0;
    wire \ALU.un2_addsub_cry_0_c_RNIJPSHDZ0 ;
    wire \ALU.r0_12_prm_2_1_c_RNOZ0 ;
    wire bfn_17_7_0_;
    wire op_1_cry_1;
    wire op_1_cry_2;
    wire op_1_cry_3;
    wire CLK_c_g;
    wire params5_g;
    wire \FTDI.N_208_0_cascade_ ;
    wire \FTDI.N_185_0_cascade_ ;
    wire \FTDI.N_207_0 ;
    wire \INVFTDI.TXstate_1C_net ;
    wire opZ0Z_0;
    wire opZ0Z_3;
    wire opZ0Z_1;
    wire \ALU.un1_op_1Z0Z_1_cascade_ ;
    wire opZ0Z_4;
    wire \ALU.un1_op_1_0 ;
    wire paramsZ0Z_1;
    wire paramsZ0Z_0;
    wire opZ0Z_2;
    wire \ALU.a_9 ;
    wire \ALU.r0_12_prm_4_9_s1_c_RNOZ0 ;
    wire \FTDI.TXstate_cnst_0_0_2_cascade_ ;
    wire \INVFTDI.TXstate_2C_net ;
    wire TXstartZ0;
    wire \FTDI.TXshiftZ0Z_1 ;
    wire TXbufferZ0Z_0;
    wire \INVFTDI.TXshift_0C_net ;
    wire \FTDI.un1_TXstate_0_sqmuxa_0_i ;
    wire bfn_18_6_0_;
    wire \FTDI.un3_TX_axb_3 ;
    wire \FTDI.un3_TX_cry_2 ;
    wire \FTDI.TXshiftZ0Z_0 ;
    wire \FTDI.un3_TX_cry_3 ;
    wire FTDI_TX_0_i;
    wire CONSTANT_ONE_NET;
    wire \FTDI.un3_TX_0_i ;
    wire \FTDI.N_185_0 ;
    wire \INVFTDI.TXstate_0C_net ;
    wire \FTDI.TXstateZ1Z_1 ;
    wire \FTDI.N_186_0 ;
    wire \FTDI.TXstate_e_1_3 ;
    wire \FTDI.N_186_0_cascade_ ;
    wire \FTDI.un3_TX_0 ;
    wire \INVFTDI.TXstate_3C_net ;
    wire \FTDI.TXstateZ1Z_0 ;
    wire \FTDI.TXstateZ0Z_3 ;
    wire \FTDI.baudAccZ0Z_2 ;
    wire \FTDI.TXstate_e_1_0 ;
    wire \FTDI.TXready ;
    wire \FTDI.baudAccZ0Z_0 ;
    wire \FTDI.baudAccZ0Z_1 ;
    wire \INVFTDI.baudAcc_0C_net ;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__57005),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__57007),
            .DIN(N__57006),
            .DOUT(N__57005),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__57007),
            .PADOUT(N__57006),
            .PADIN(N__57005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TX_obuf_iopad (
            .OE(N__56996),
            .DIN(N__56995),
            .DOUT(N__56994),
            .PACKAGEPIN(TX));
    defparam TX_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TX_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TX_obuf_preio (
            .PADOEN(N__56996),
            .PADOUT(N__56995),
            .PADIN(N__56994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__56524),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO3_obuf_iopad (
            .OE(N__56987),
            .DIN(N__56986),
            .DOUT(N__56985),
            .PACKAGEPIN(GPIO3));
    defparam GPIO3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO3_obuf_preio (
            .PADOEN(N__56987),
            .PADOUT(N__56986),
            .PADIN(N__56985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO11_obuf_iopad (
            .OE(N__56978),
            .DIN(N__56977),
            .DOUT(N__56976),
            .PACKAGEPIN(GPIO11));
    defparam GPIO11_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO11_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO11_obuf_preio (
            .PADOEN(N__56978),
            .PADOUT(N__56977),
            .PADIN(N__56976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO9_obuf_iopad (
            .OE(N__56969),
            .DIN(N__56968),
            .DOUT(N__56967),
            .PACKAGEPIN(GPIO9));
    defparam GPIO9_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO9_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO9_obuf_preio (
            .PADOEN(N__56969),
            .PADOUT(N__56968),
            .PADIN(N__56967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__56397),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__14264 (
            .O(N__56950),
            .I(N__56942));
    InMux I__14263 (
            .O(N__56949),
            .I(N__56937));
    InMux I__14262 (
            .O(N__56948),
            .I(N__56937));
    InMux I__14261 (
            .O(N__56947),
            .I(N__56932));
    InMux I__14260 (
            .O(N__56946),
            .I(N__56932));
    InMux I__14259 (
            .O(N__56945),
            .I(N__56929));
    LocalMux I__14258 (
            .O(N__56942),
            .I(\FTDI.TXstateZ1Z_1 ));
    LocalMux I__14257 (
            .O(N__56937),
            .I(\FTDI.TXstateZ1Z_1 ));
    LocalMux I__14256 (
            .O(N__56932),
            .I(\FTDI.TXstateZ1Z_1 ));
    LocalMux I__14255 (
            .O(N__56929),
            .I(\FTDI.TXstateZ1Z_1 ));
    InMux I__14254 (
            .O(N__56920),
            .I(N__56917));
    LocalMux I__14253 (
            .O(N__56917),
            .I(\FTDI.N_186_0 ));
    InMux I__14252 (
            .O(N__56914),
            .I(N__56911));
    LocalMux I__14251 (
            .O(N__56911),
            .I(\FTDI.TXstate_e_1_3 ));
    CascadeMux I__14250 (
            .O(N__56908),
            .I(\FTDI.N_186_0_cascade_ ));
    InMux I__14249 (
            .O(N__56905),
            .I(N__56901));
    CascadeMux I__14248 (
            .O(N__56904),
            .I(N__56897));
    LocalMux I__14247 (
            .O(N__56901),
            .I(N__56891));
    InMux I__14246 (
            .O(N__56900),
            .I(N__56888));
    InMux I__14245 (
            .O(N__56897),
            .I(N__56885));
    InMux I__14244 (
            .O(N__56896),
            .I(N__56882));
    InMux I__14243 (
            .O(N__56895),
            .I(N__56877));
    InMux I__14242 (
            .O(N__56894),
            .I(N__56877));
    Odrv4 I__14241 (
            .O(N__56891),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__14240 (
            .O(N__56888),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__14239 (
            .O(N__56885),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__14238 (
            .O(N__56882),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__14237 (
            .O(N__56877),
            .I(\FTDI.un3_TX_0 ));
    InMux I__14236 (
            .O(N__56866),
            .I(N__56858));
    InMux I__14235 (
            .O(N__56865),
            .I(N__56851));
    InMux I__14234 (
            .O(N__56864),
            .I(N__56851));
    InMux I__14233 (
            .O(N__56863),
            .I(N__56851));
    InMux I__14232 (
            .O(N__56862),
            .I(N__56846));
    InMux I__14231 (
            .O(N__56861),
            .I(N__56846));
    LocalMux I__14230 (
            .O(N__56858),
            .I(\FTDI.TXstateZ1Z_0 ));
    LocalMux I__14229 (
            .O(N__56851),
            .I(\FTDI.TXstateZ1Z_0 ));
    LocalMux I__14228 (
            .O(N__56846),
            .I(\FTDI.TXstateZ1Z_0 ));
    InMux I__14227 (
            .O(N__56839),
            .I(N__56826));
    InMux I__14226 (
            .O(N__56838),
            .I(N__56826));
    InMux I__14225 (
            .O(N__56837),
            .I(N__56817));
    InMux I__14224 (
            .O(N__56836),
            .I(N__56817));
    InMux I__14223 (
            .O(N__56835),
            .I(N__56817));
    InMux I__14222 (
            .O(N__56834),
            .I(N__56817));
    InMux I__14221 (
            .O(N__56833),
            .I(N__56811));
    InMux I__14220 (
            .O(N__56832),
            .I(N__56811));
    InMux I__14219 (
            .O(N__56831),
            .I(N__56807));
    LocalMux I__14218 (
            .O(N__56826),
            .I(N__56804));
    LocalMux I__14217 (
            .O(N__56817),
            .I(N__56801));
    CascadeMux I__14216 (
            .O(N__56816),
            .I(N__56792));
    LocalMux I__14215 (
            .O(N__56811),
            .I(N__56789));
    InMux I__14214 (
            .O(N__56810),
            .I(N__56786));
    LocalMux I__14213 (
            .O(N__56807),
            .I(N__56781));
    Span4Mux_v I__14212 (
            .O(N__56804),
            .I(N__56781));
    Span4Mux_h I__14211 (
            .O(N__56801),
            .I(N__56778));
    InMux I__14210 (
            .O(N__56800),
            .I(N__56773));
    InMux I__14209 (
            .O(N__56799),
            .I(N__56773));
    InMux I__14208 (
            .O(N__56798),
            .I(N__56768));
    InMux I__14207 (
            .O(N__56797),
            .I(N__56768));
    InMux I__14206 (
            .O(N__56796),
            .I(N__56763));
    InMux I__14205 (
            .O(N__56795),
            .I(N__56763));
    InMux I__14204 (
            .O(N__56792),
            .I(N__56760));
    Odrv4 I__14203 (
            .O(N__56789),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__14202 (
            .O(N__56786),
            .I(\FTDI.TXstateZ0Z_3 ));
    Odrv4 I__14201 (
            .O(N__56781),
            .I(\FTDI.TXstateZ0Z_3 ));
    Odrv4 I__14200 (
            .O(N__56778),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__14199 (
            .O(N__56773),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__14198 (
            .O(N__56768),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__14197 (
            .O(N__56763),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__14196 (
            .O(N__56760),
            .I(\FTDI.TXstateZ0Z_3 ));
    InMux I__14195 (
            .O(N__56743),
            .I(N__56732));
    InMux I__14194 (
            .O(N__56742),
            .I(N__56732));
    InMux I__14193 (
            .O(N__56741),
            .I(N__56727));
    InMux I__14192 (
            .O(N__56740),
            .I(N__56727));
    InMux I__14191 (
            .O(N__56739),
            .I(N__56720));
    InMux I__14190 (
            .O(N__56738),
            .I(N__56720));
    InMux I__14189 (
            .O(N__56737),
            .I(N__56720));
    LocalMux I__14188 (
            .O(N__56732),
            .I(\FTDI.baudAccZ0Z_2 ));
    LocalMux I__14187 (
            .O(N__56727),
            .I(\FTDI.baudAccZ0Z_2 ));
    LocalMux I__14186 (
            .O(N__56720),
            .I(\FTDI.baudAccZ0Z_2 ));
    CascadeMux I__14185 (
            .O(N__56713),
            .I(N__56710));
    InMux I__14184 (
            .O(N__56710),
            .I(N__56707));
    LocalMux I__14183 (
            .O(N__56707),
            .I(\FTDI.TXstate_e_1_0 ));
    InMux I__14182 (
            .O(N__56704),
            .I(N__56696));
    InMux I__14181 (
            .O(N__56703),
            .I(N__56696));
    CascadeMux I__14180 (
            .O(N__56702),
            .I(N__56692));
    InMux I__14179 (
            .O(N__56701),
            .I(N__56689));
    LocalMux I__14178 (
            .O(N__56696),
            .I(N__56686));
    InMux I__14177 (
            .O(N__56695),
            .I(N__56681));
    InMux I__14176 (
            .O(N__56692),
            .I(N__56681));
    LocalMux I__14175 (
            .O(N__56689),
            .I(\FTDI.TXready ));
    Odrv4 I__14174 (
            .O(N__56686),
            .I(\FTDI.TXready ));
    LocalMux I__14173 (
            .O(N__56681),
            .I(\FTDI.TXready ));
    CascadeMux I__14172 (
            .O(N__56674),
            .I(N__56670));
    InMux I__14171 (
            .O(N__56673),
            .I(N__56666));
    InMux I__14170 (
            .O(N__56670),
            .I(N__56661));
    InMux I__14169 (
            .O(N__56669),
            .I(N__56661));
    LocalMux I__14168 (
            .O(N__56666),
            .I(\FTDI.baudAccZ0Z_0 ));
    LocalMux I__14167 (
            .O(N__56661),
            .I(\FTDI.baudAccZ0Z_0 ));
    InMux I__14166 (
            .O(N__56656),
            .I(N__56652));
    InMux I__14165 (
            .O(N__56655),
            .I(N__56649));
    LocalMux I__14164 (
            .O(N__56652),
            .I(\FTDI.baudAccZ0Z_1 ));
    LocalMux I__14163 (
            .O(N__56649),
            .I(\FTDI.baudAccZ0Z_1 ));
    CascadeMux I__14162 (
            .O(N__56644),
            .I(\FTDI.TXstate_cnst_0_0_2_cascade_ ));
    InMux I__14161 (
            .O(N__56641),
            .I(N__56635));
    InMux I__14160 (
            .O(N__56640),
            .I(N__56635));
    LocalMux I__14159 (
            .O(N__56635),
            .I(N__56632));
    Span4Mux_v I__14158 (
            .O(N__56632),
            .I(N__56629));
    Span4Mux_v I__14157 (
            .O(N__56629),
            .I(N__56626));
    Sp12to4 I__14156 (
            .O(N__56626),
            .I(N__56623));
    Span12Mux_h I__14155 (
            .O(N__56623),
            .I(N__56620));
    Odrv12 I__14154 (
            .O(N__56620),
            .I(TXstartZ0));
    InMux I__14153 (
            .O(N__56617),
            .I(N__56614));
    LocalMux I__14152 (
            .O(N__56614),
            .I(\FTDI.TXshiftZ0Z_1 ));
    InMux I__14151 (
            .O(N__56611),
            .I(N__56608));
    LocalMux I__14150 (
            .O(N__56608),
            .I(N__56605));
    Span4Mux_v I__14149 (
            .O(N__56605),
            .I(N__56602));
    Sp12to4 I__14148 (
            .O(N__56602),
            .I(N__56599));
    Span12Mux_h I__14147 (
            .O(N__56599),
            .I(N__56596));
    Odrv12 I__14146 (
            .O(N__56596),
            .I(TXbufferZ0Z_0));
    CEMux I__14145 (
            .O(N__56593),
            .I(N__56590));
    LocalMux I__14144 (
            .O(N__56590),
            .I(N__56587));
    Span4Mux_v I__14143 (
            .O(N__56587),
            .I(N__56583));
    CEMux I__14142 (
            .O(N__56586),
            .I(N__56580));
    Span4Mux_v I__14141 (
            .O(N__56583),
            .I(N__56573));
    LocalMux I__14140 (
            .O(N__56580),
            .I(N__56573));
    CEMux I__14139 (
            .O(N__56579),
            .I(N__56570));
    CEMux I__14138 (
            .O(N__56578),
            .I(N__56567));
    Span4Mux_v I__14137 (
            .O(N__56573),
            .I(N__56564));
    LocalMux I__14136 (
            .O(N__56570),
            .I(N__56561));
    LocalMux I__14135 (
            .O(N__56567),
            .I(N__56558));
    Span4Mux_v I__14134 (
            .O(N__56564),
            .I(N__56555));
    Span4Mux_v I__14133 (
            .O(N__56561),
            .I(N__56550));
    Span4Mux_h I__14132 (
            .O(N__56558),
            .I(N__56550));
    Odrv4 I__14131 (
            .O(N__56555),
            .I(\FTDI.un1_TXstate_0_sqmuxa_0_i ));
    Odrv4 I__14130 (
            .O(N__56550),
            .I(\FTDI.un1_TXstate_0_sqmuxa_0_i ));
    InMux I__14129 (
            .O(N__56545),
            .I(N__56542));
    LocalMux I__14128 (
            .O(N__56542),
            .I(\FTDI.un3_TX_axb_3 ));
    InMux I__14127 (
            .O(N__56539),
            .I(N__56536));
    LocalMux I__14126 (
            .O(N__56536),
            .I(N__56533));
    Span4Mux_v I__14125 (
            .O(N__56533),
            .I(N__56530));
    Odrv4 I__14124 (
            .O(N__56530),
            .I(\FTDI.TXshiftZ0Z_0 ));
    InMux I__14123 (
            .O(N__56527),
            .I(\FTDI.un3_TX_cry_3 ));
    IoInMux I__14122 (
            .O(N__56524),
            .I(N__56521));
    LocalMux I__14121 (
            .O(N__56521),
            .I(N__56518));
    Span12Mux_s5_v I__14120 (
            .O(N__56518),
            .I(N__56515));
    Odrv12 I__14119 (
            .O(N__56515),
            .I(FTDI_TX_0_i));
    CascadeMux I__14118 (
            .O(N__56512),
            .I(N__56509));
    InMux I__14117 (
            .O(N__56509),
            .I(N__56501));
    CascadeMux I__14116 (
            .O(N__56508),
            .I(N__56498));
    CascadeMux I__14115 (
            .O(N__56507),
            .I(N__56495));
    CascadeMux I__14114 (
            .O(N__56506),
            .I(N__56492));
    InMux I__14113 (
            .O(N__56505),
            .I(N__56489));
    CascadeMux I__14112 (
            .O(N__56504),
            .I(N__56485));
    LocalMux I__14111 (
            .O(N__56501),
            .I(N__56482));
    InMux I__14110 (
            .O(N__56498),
            .I(N__56478));
    InMux I__14109 (
            .O(N__56495),
            .I(N__56472));
    InMux I__14108 (
            .O(N__56492),
            .I(N__56469));
    LocalMux I__14107 (
            .O(N__56489),
            .I(N__56466));
    InMux I__14106 (
            .O(N__56488),
            .I(N__56463));
    InMux I__14105 (
            .O(N__56485),
            .I(N__56460));
    Span4Mux_s1_v I__14104 (
            .O(N__56482),
            .I(N__56457));
    CascadeMux I__14103 (
            .O(N__56481),
            .I(N__56454));
    LocalMux I__14102 (
            .O(N__56478),
            .I(N__56451));
    CascadeMux I__14101 (
            .O(N__56477),
            .I(N__56448));
    CascadeMux I__14100 (
            .O(N__56476),
            .I(N__56445));
    CascadeMux I__14099 (
            .O(N__56475),
            .I(N__56442));
    LocalMux I__14098 (
            .O(N__56472),
            .I(N__56437));
    LocalMux I__14097 (
            .O(N__56469),
            .I(N__56437));
    Span4Mux_v I__14096 (
            .O(N__56466),
            .I(N__56434));
    LocalMux I__14095 (
            .O(N__56463),
            .I(N__56431));
    LocalMux I__14094 (
            .O(N__56460),
            .I(N__56426));
    Span4Mux_h I__14093 (
            .O(N__56457),
            .I(N__56426));
    InMux I__14092 (
            .O(N__56454),
            .I(N__56423));
    Span4Mux_v I__14091 (
            .O(N__56451),
            .I(N__56420));
    InMux I__14090 (
            .O(N__56448),
            .I(N__56417));
    InMux I__14089 (
            .O(N__56445),
            .I(N__56414));
    InMux I__14088 (
            .O(N__56442),
            .I(N__56410));
    Span4Mux_v I__14087 (
            .O(N__56437),
            .I(N__56399));
    Span4Mux_h I__14086 (
            .O(N__56434),
            .I(N__56399));
    Span4Mux_v I__14085 (
            .O(N__56431),
            .I(N__56399));
    Span4Mux_v I__14084 (
            .O(N__56426),
            .I(N__56399));
    LocalMux I__14083 (
            .O(N__56423),
            .I(N__56399));
    Span4Mux_v I__14082 (
            .O(N__56420),
            .I(N__56394));
    LocalMux I__14081 (
            .O(N__56417),
            .I(N__56389));
    LocalMux I__14080 (
            .O(N__56414),
            .I(N__56389));
    CascadeMux I__14079 (
            .O(N__56413),
            .I(N__56386));
    LocalMux I__14078 (
            .O(N__56410),
            .I(N__56381));
    Span4Mux_v I__14077 (
            .O(N__56399),
            .I(N__56381));
    InMux I__14076 (
            .O(N__56398),
            .I(N__56378));
    IoInMux I__14075 (
            .O(N__56397),
            .I(N__56375));
    Span4Mux_v I__14074 (
            .O(N__56394),
            .I(N__56372));
    Span4Mux_v I__14073 (
            .O(N__56389),
            .I(N__56369));
    InMux I__14072 (
            .O(N__56386),
            .I(N__56366));
    Span4Mux_h I__14071 (
            .O(N__56381),
            .I(N__56363));
    LocalMux I__14070 (
            .O(N__56378),
            .I(N__56360));
    LocalMux I__14069 (
            .O(N__56375),
            .I(N__56357));
    Sp12to4 I__14068 (
            .O(N__56372),
            .I(N__56354));
    Span4Mux_h I__14067 (
            .O(N__56369),
            .I(N__56351));
    LocalMux I__14066 (
            .O(N__56366),
            .I(N__56348));
    Span4Mux_h I__14065 (
            .O(N__56363),
            .I(N__56343));
    Span4Mux_v I__14064 (
            .O(N__56360),
            .I(N__56343));
    Span12Mux_s10_v I__14063 (
            .O(N__56357),
            .I(N__56334));
    Span12Mux_h I__14062 (
            .O(N__56354),
            .I(N__56334));
    Sp12to4 I__14061 (
            .O(N__56351),
            .I(N__56334));
    Sp12to4 I__14060 (
            .O(N__56348),
            .I(N__56334));
    Sp12to4 I__14059 (
            .O(N__56343),
            .I(N__56331));
    Span12Mux_v I__14058 (
            .O(N__56334),
            .I(N__56326));
    Span12Mux_s5_h I__14057 (
            .O(N__56331),
            .I(N__56326));
    Odrv12 I__14056 (
            .O(N__56326),
            .I(CONSTANT_ONE_NET));
    InMux I__14055 (
            .O(N__56323),
            .I(N__56319));
    InMux I__14054 (
            .O(N__56322),
            .I(N__56316));
    LocalMux I__14053 (
            .O(N__56319),
            .I(\FTDI.un3_TX_0_i ));
    LocalMux I__14052 (
            .O(N__56316),
            .I(\FTDI.un3_TX_0_i ));
    InMux I__14051 (
            .O(N__56311),
            .I(N__56308));
    LocalMux I__14050 (
            .O(N__56308),
            .I(\FTDI.N_185_0 ));
    ClkMux I__14049 (
            .O(N__56305),
            .I(N__56065));
    ClkMux I__14048 (
            .O(N__56304),
            .I(N__56065));
    ClkMux I__14047 (
            .O(N__56303),
            .I(N__56065));
    ClkMux I__14046 (
            .O(N__56302),
            .I(N__56065));
    ClkMux I__14045 (
            .O(N__56301),
            .I(N__56065));
    ClkMux I__14044 (
            .O(N__56300),
            .I(N__56065));
    ClkMux I__14043 (
            .O(N__56299),
            .I(N__56065));
    ClkMux I__14042 (
            .O(N__56298),
            .I(N__56065));
    ClkMux I__14041 (
            .O(N__56297),
            .I(N__56065));
    ClkMux I__14040 (
            .O(N__56296),
            .I(N__56065));
    ClkMux I__14039 (
            .O(N__56295),
            .I(N__56065));
    ClkMux I__14038 (
            .O(N__56294),
            .I(N__56065));
    ClkMux I__14037 (
            .O(N__56293),
            .I(N__56065));
    ClkMux I__14036 (
            .O(N__56292),
            .I(N__56065));
    ClkMux I__14035 (
            .O(N__56291),
            .I(N__56065));
    ClkMux I__14034 (
            .O(N__56290),
            .I(N__56065));
    ClkMux I__14033 (
            .O(N__56289),
            .I(N__56065));
    ClkMux I__14032 (
            .O(N__56288),
            .I(N__56065));
    ClkMux I__14031 (
            .O(N__56287),
            .I(N__56065));
    ClkMux I__14030 (
            .O(N__56286),
            .I(N__56065));
    ClkMux I__14029 (
            .O(N__56285),
            .I(N__56065));
    ClkMux I__14028 (
            .O(N__56284),
            .I(N__56065));
    ClkMux I__14027 (
            .O(N__56283),
            .I(N__56065));
    ClkMux I__14026 (
            .O(N__56282),
            .I(N__56065));
    ClkMux I__14025 (
            .O(N__56281),
            .I(N__56065));
    ClkMux I__14024 (
            .O(N__56280),
            .I(N__56065));
    ClkMux I__14023 (
            .O(N__56279),
            .I(N__56065));
    ClkMux I__14022 (
            .O(N__56278),
            .I(N__56065));
    ClkMux I__14021 (
            .O(N__56277),
            .I(N__56065));
    ClkMux I__14020 (
            .O(N__56276),
            .I(N__56065));
    ClkMux I__14019 (
            .O(N__56275),
            .I(N__56065));
    ClkMux I__14018 (
            .O(N__56274),
            .I(N__56065));
    ClkMux I__14017 (
            .O(N__56273),
            .I(N__56065));
    ClkMux I__14016 (
            .O(N__56272),
            .I(N__56065));
    ClkMux I__14015 (
            .O(N__56271),
            .I(N__56065));
    ClkMux I__14014 (
            .O(N__56270),
            .I(N__56065));
    ClkMux I__14013 (
            .O(N__56269),
            .I(N__56065));
    ClkMux I__14012 (
            .O(N__56268),
            .I(N__56065));
    ClkMux I__14011 (
            .O(N__56267),
            .I(N__56065));
    ClkMux I__14010 (
            .O(N__56266),
            .I(N__56065));
    ClkMux I__14009 (
            .O(N__56265),
            .I(N__56065));
    ClkMux I__14008 (
            .O(N__56264),
            .I(N__56065));
    ClkMux I__14007 (
            .O(N__56263),
            .I(N__56065));
    ClkMux I__14006 (
            .O(N__56262),
            .I(N__56065));
    ClkMux I__14005 (
            .O(N__56261),
            .I(N__56065));
    ClkMux I__14004 (
            .O(N__56260),
            .I(N__56065));
    ClkMux I__14003 (
            .O(N__56259),
            .I(N__56065));
    ClkMux I__14002 (
            .O(N__56258),
            .I(N__56065));
    ClkMux I__14001 (
            .O(N__56257),
            .I(N__56065));
    ClkMux I__14000 (
            .O(N__56256),
            .I(N__56065));
    ClkMux I__13999 (
            .O(N__56255),
            .I(N__56065));
    ClkMux I__13998 (
            .O(N__56254),
            .I(N__56065));
    ClkMux I__13997 (
            .O(N__56253),
            .I(N__56065));
    ClkMux I__13996 (
            .O(N__56252),
            .I(N__56065));
    ClkMux I__13995 (
            .O(N__56251),
            .I(N__56065));
    ClkMux I__13994 (
            .O(N__56250),
            .I(N__56065));
    ClkMux I__13993 (
            .O(N__56249),
            .I(N__56065));
    ClkMux I__13992 (
            .O(N__56248),
            .I(N__56065));
    ClkMux I__13991 (
            .O(N__56247),
            .I(N__56065));
    ClkMux I__13990 (
            .O(N__56246),
            .I(N__56065));
    ClkMux I__13989 (
            .O(N__56245),
            .I(N__56065));
    ClkMux I__13988 (
            .O(N__56244),
            .I(N__56065));
    ClkMux I__13987 (
            .O(N__56243),
            .I(N__56065));
    ClkMux I__13986 (
            .O(N__56242),
            .I(N__56065));
    ClkMux I__13985 (
            .O(N__56241),
            .I(N__56065));
    ClkMux I__13984 (
            .O(N__56240),
            .I(N__56065));
    ClkMux I__13983 (
            .O(N__56239),
            .I(N__56065));
    ClkMux I__13982 (
            .O(N__56238),
            .I(N__56065));
    ClkMux I__13981 (
            .O(N__56237),
            .I(N__56065));
    ClkMux I__13980 (
            .O(N__56236),
            .I(N__56065));
    ClkMux I__13979 (
            .O(N__56235),
            .I(N__56065));
    ClkMux I__13978 (
            .O(N__56234),
            .I(N__56065));
    ClkMux I__13977 (
            .O(N__56233),
            .I(N__56065));
    ClkMux I__13976 (
            .O(N__56232),
            .I(N__56065));
    ClkMux I__13975 (
            .O(N__56231),
            .I(N__56065));
    ClkMux I__13974 (
            .O(N__56230),
            .I(N__56065));
    ClkMux I__13973 (
            .O(N__56229),
            .I(N__56065));
    ClkMux I__13972 (
            .O(N__56228),
            .I(N__56065));
    ClkMux I__13971 (
            .O(N__56227),
            .I(N__56065));
    ClkMux I__13970 (
            .O(N__56226),
            .I(N__56065));
    GlobalMux I__13969 (
            .O(N__56065),
            .I(N__56062));
    gio2CtrlBuf I__13968 (
            .O(N__56062),
            .I(CLK_c_g));
    CEMux I__13967 (
            .O(N__56059),
            .I(N__55987));
    CEMux I__13966 (
            .O(N__56058),
            .I(N__55987));
    CEMux I__13965 (
            .O(N__56057),
            .I(N__55987));
    CEMux I__13964 (
            .O(N__56056),
            .I(N__55987));
    CEMux I__13963 (
            .O(N__56055),
            .I(N__55987));
    CEMux I__13962 (
            .O(N__56054),
            .I(N__55987));
    CEMux I__13961 (
            .O(N__56053),
            .I(N__55987));
    CEMux I__13960 (
            .O(N__56052),
            .I(N__55987));
    CEMux I__13959 (
            .O(N__56051),
            .I(N__55987));
    CEMux I__13958 (
            .O(N__56050),
            .I(N__55987));
    CEMux I__13957 (
            .O(N__56049),
            .I(N__55987));
    CEMux I__13956 (
            .O(N__56048),
            .I(N__55987));
    CEMux I__13955 (
            .O(N__56047),
            .I(N__55987));
    CEMux I__13954 (
            .O(N__56046),
            .I(N__55987));
    CEMux I__13953 (
            .O(N__56045),
            .I(N__55987));
    CEMux I__13952 (
            .O(N__56044),
            .I(N__55987));
    CEMux I__13951 (
            .O(N__56043),
            .I(N__55987));
    CEMux I__13950 (
            .O(N__56042),
            .I(N__55987));
    CEMux I__13949 (
            .O(N__56041),
            .I(N__55987));
    CEMux I__13948 (
            .O(N__56040),
            .I(N__55987));
    CEMux I__13947 (
            .O(N__56039),
            .I(N__55987));
    CEMux I__13946 (
            .O(N__56038),
            .I(N__55987));
    CEMux I__13945 (
            .O(N__56037),
            .I(N__55987));
    CEMux I__13944 (
            .O(N__56036),
            .I(N__55987));
    GlobalMux I__13943 (
            .O(N__55987),
            .I(N__55984));
    gio2CtrlBuf I__13942 (
            .O(N__55984),
            .I(params5_g));
    CascadeMux I__13941 (
            .O(N__55981),
            .I(\FTDI.N_208_0_cascade_ ));
    CascadeMux I__13940 (
            .O(N__55978),
            .I(\FTDI.N_185_0_cascade_ ));
    InMux I__13939 (
            .O(N__55975),
            .I(N__55972));
    LocalMux I__13938 (
            .O(N__55972),
            .I(\FTDI.N_207_0 ));
    InMux I__13937 (
            .O(N__55969),
            .I(N__55965));
    InMux I__13936 (
            .O(N__55968),
            .I(N__55962));
    LocalMux I__13935 (
            .O(N__55965),
            .I(N__55952));
    LocalMux I__13934 (
            .O(N__55962),
            .I(N__55947));
    CascadeMux I__13933 (
            .O(N__55961),
            .I(N__55943));
    InMux I__13932 (
            .O(N__55960),
            .I(N__55934));
    InMux I__13931 (
            .O(N__55959),
            .I(N__55934));
    InMux I__13930 (
            .O(N__55958),
            .I(N__55924));
    InMux I__13929 (
            .O(N__55957),
            .I(N__55921));
    CascadeMux I__13928 (
            .O(N__55956),
            .I(N__55916));
    CascadeMux I__13927 (
            .O(N__55955),
            .I(N__55913));
    Span4Mux_h I__13926 (
            .O(N__55952),
            .I(N__55910));
    InMux I__13925 (
            .O(N__55951),
            .I(N__55905));
    InMux I__13924 (
            .O(N__55950),
            .I(N__55905));
    Span4Mux_h I__13923 (
            .O(N__55947),
            .I(N__55896));
    InMux I__13922 (
            .O(N__55946),
            .I(N__55893));
    InMux I__13921 (
            .O(N__55943),
            .I(N__55888));
    InMux I__13920 (
            .O(N__55942),
            .I(N__55888));
    InMux I__13919 (
            .O(N__55941),
            .I(N__55885));
    InMux I__13918 (
            .O(N__55940),
            .I(N__55882));
    InMux I__13917 (
            .O(N__55939),
            .I(N__55879));
    LocalMux I__13916 (
            .O(N__55934),
            .I(N__55876));
    InMux I__13915 (
            .O(N__55933),
            .I(N__55871));
    InMux I__13914 (
            .O(N__55932),
            .I(N__55871));
    InMux I__13913 (
            .O(N__55931),
            .I(N__55862));
    InMux I__13912 (
            .O(N__55930),
            .I(N__55862));
    InMux I__13911 (
            .O(N__55929),
            .I(N__55862));
    InMux I__13910 (
            .O(N__55928),
            .I(N__55862));
    InMux I__13909 (
            .O(N__55927),
            .I(N__55858));
    LocalMux I__13908 (
            .O(N__55924),
            .I(N__55853));
    LocalMux I__13907 (
            .O(N__55921),
            .I(N__55853));
    InMux I__13906 (
            .O(N__55920),
            .I(N__55848));
    InMux I__13905 (
            .O(N__55919),
            .I(N__55848));
    InMux I__13904 (
            .O(N__55916),
            .I(N__55842));
    InMux I__13903 (
            .O(N__55913),
            .I(N__55842));
    Span4Mux_h I__13902 (
            .O(N__55910),
            .I(N__55834));
    LocalMux I__13901 (
            .O(N__55905),
            .I(N__55834));
    InMux I__13900 (
            .O(N__55904),
            .I(N__55831));
    InMux I__13899 (
            .O(N__55903),
            .I(N__55826));
    InMux I__13898 (
            .O(N__55902),
            .I(N__55826));
    InMux I__13897 (
            .O(N__55901),
            .I(N__55819));
    InMux I__13896 (
            .O(N__55900),
            .I(N__55819));
    InMux I__13895 (
            .O(N__55899),
            .I(N__55819));
    Span4Mux_h I__13894 (
            .O(N__55896),
            .I(N__55814));
    LocalMux I__13893 (
            .O(N__55893),
            .I(N__55809));
    LocalMux I__13892 (
            .O(N__55888),
            .I(N__55809));
    LocalMux I__13891 (
            .O(N__55885),
            .I(N__55802));
    LocalMux I__13890 (
            .O(N__55882),
            .I(N__55787));
    LocalMux I__13889 (
            .O(N__55879),
            .I(N__55787));
    Span4Mux_v I__13888 (
            .O(N__55876),
            .I(N__55787));
    LocalMux I__13887 (
            .O(N__55871),
            .I(N__55787));
    LocalMux I__13886 (
            .O(N__55862),
            .I(N__55787));
    InMux I__13885 (
            .O(N__55861),
            .I(N__55784));
    LocalMux I__13884 (
            .O(N__55858),
            .I(N__55777));
    Span4Mux_v I__13883 (
            .O(N__55853),
            .I(N__55777));
    LocalMux I__13882 (
            .O(N__55848),
            .I(N__55777));
    CascadeMux I__13881 (
            .O(N__55847),
            .I(N__55773));
    LocalMux I__13880 (
            .O(N__55842),
            .I(N__55769));
    InMux I__13879 (
            .O(N__55841),
            .I(N__55766));
    InMux I__13878 (
            .O(N__55840),
            .I(N__55763));
    CascadeMux I__13877 (
            .O(N__55839),
            .I(N__55760));
    Span4Mux_h I__13876 (
            .O(N__55834),
            .I(N__55754));
    LocalMux I__13875 (
            .O(N__55831),
            .I(N__55754));
    LocalMux I__13874 (
            .O(N__55826),
            .I(N__55749));
    LocalMux I__13873 (
            .O(N__55819),
            .I(N__55749));
    InMux I__13872 (
            .O(N__55818),
            .I(N__55744));
    InMux I__13871 (
            .O(N__55817),
            .I(N__55744));
    Span4Mux_v I__13870 (
            .O(N__55814),
            .I(N__55741));
    Span4Mux_h I__13869 (
            .O(N__55809),
            .I(N__55738));
    InMux I__13868 (
            .O(N__55808),
            .I(N__55731));
    InMux I__13867 (
            .O(N__55807),
            .I(N__55731));
    InMux I__13866 (
            .O(N__55806),
            .I(N__55724));
    InMux I__13865 (
            .O(N__55805),
            .I(N__55724));
    Span4Mux_h I__13864 (
            .O(N__55802),
            .I(N__55719));
    InMux I__13863 (
            .O(N__55801),
            .I(N__55716));
    InMux I__13862 (
            .O(N__55800),
            .I(N__55709));
    InMux I__13861 (
            .O(N__55799),
            .I(N__55709));
    InMux I__13860 (
            .O(N__55798),
            .I(N__55709));
    Span4Mux_v I__13859 (
            .O(N__55787),
            .I(N__55706));
    LocalMux I__13858 (
            .O(N__55784),
            .I(N__55701));
    Span4Mux_v I__13857 (
            .O(N__55777),
            .I(N__55701));
    InMux I__13856 (
            .O(N__55776),
            .I(N__55694));
    InMux I__13855 (
            .O(N__55773),
            .I(N__55694));
    InMux I__13854 (
            .O(N__55772),
            .I(N__55694));
    Span4Mux_h I__13853 (
            .O(N__55769),
            .I(N__55690));
    LocalMux I__13852 (
            .O(N__55766),
            .I(N__55685));
    LocalMux I__13851 (
            .O(N__55763),
            .I(N__55685));
    InMux I__13850 (
            .O(N__55760),
            .I(N__55682));
    InMux I__13849 (
            .O(N__55759),
            .I(N__55679));
    Span4Mux_h I__13848 (
            .O(N__55754),
            .I(N__55676));
    Span4Mux_v I__13847 (
            .O(N__55749),
            .I(N__55671));
    LocalMux I__13846 (
            .O(N__55744),
            .I(N__55671));
    Span4Mux_h I__13845 (
            .O(N__55741),
            .I(N__55666));
    Span4Mux_v I__13844 (
            .O(N__55738),
            .I(N__55666));
    InMux I__13843 (
            .O(N__55737),
            .I(N__55663));
    InMux I__13842 (
            .O(N__55736),
            .I(N__55660));
    LocalMux I__13841 (
            .O(N__55731),
            .I(N__55656));
    InMux I__13840 (
            .O(N__55730),
            .I(N__55653));
    InMux I__13839 (
            .O(N__55729),
            .I(N__55650));
    LocalMux I__13838 (
            .O(N__55724),
            .I(N__55647));
    InMux I__13837 (
            .O(N__55723),
            .I(N__55642));
    InMux I__13836 (
            .O(N__55722),
            .I(N__55642));
    Span4Mux_h I__13835 (
            .O(N__55719),
            .I(N__55631));
    LocalMux I__13834 (
            .O(N__55716),
            .I(N__55631));
    LocalMux I__13833 (
            .O(N__55709),
            .I(N__55631));
    Span4Mux_h I__13832 (
            .O(N__55706),
            .I(N__55631));
    Sp12to4 I__13831 (
            .O(N__55701),
            .I(N__55626));
    LocalMux I__13830 (
            .O(N__55694),
            .I(N__55626));
    InMux I__13829 (
            .O(N__55693),
            .I(N__55623));
    Span4Mux_h I__13828 (
            .O(N__55690),
            .I(N__55618));
    Span4Mux_h I__13827 (
            .O(N__55685),
            .I(N__55618));
    LocalMux I__13826 (
            .O(N__55682),
            .I(N__55609));
    LocalMux I__13825 (
            .O(N__55679),
            .I(N__55609));
    Span4Mux_v I__13824 (
            .O(N__55676),
            .I(N__55609));
    Span4Mux_h I__13823 (
            .O(N__55671),
            .I(N__55609));
    Span4Mux_v I__13822 (
            .O(N__55666),
            .I(N__55604));
    LocalMux I__13821 (
            .O(N__55663),
            .I(N__55604));
    LocalMux I__13820 (
            .O(N__55660),
            .I(N__55601));
    InMux I__13819 (
            .O(N__55659),
            .I(N__55598));
    Span4Mux_h I__13818 (
            .O(N__55656),
            .I(N__55589));
    LocalMux I__13817 (
            .O(N__55653),
            .I(N__55589));
    LocalMux I__13816 (
            .O(N__55650),
            .I(N__55589));
    Span4Mux_h I__13815 (
            .O(N__55647),
            .I(N__55589));
    LocalMux I__13814 (
            .O(N__55642),
            .I(N__55586));
    InMux I__13813 (
            .O(N__55641),
            .I(N__55582));
    InMux I__13812 (
            .O(N__55640),
            .I(N__55579));
    Sp12to4 I__13811 (
            .O(N__55631),
            .I(N__55574));
    Span12Mux_h I__13810 (
            .O(N__55626),
            .I(N__55574));
    LocalMux I__13809 (
            .O(N__55623),
            .I(N__55567));
    Span4Mux_h I__13808 (
            .O(N__55618),
            .I(N__55567));
    Span4Mux_v I__13807 (
            .O(N__55609),
            .I(N__55567));
    Span4Mux_h I__13806 (
            .O(N__55604),
            .I(N__55564));
    Span4Mux_h I__13805 (
            .O(N__55601),
            .I(N__55555));
    LocalMux I__13804 (
            .O(N__55598),
            .I(N__55555));
    Span4Mux_v I__13803 (
            .O(N__55589),
            .I(N__55555));
    Span4Mux_s2_v I__13802 (
            .O(N__55586),
            .I(N__55555));
    InMux I__13801 (
            .O(N__55585),
            .I(N__55552));
    LocalMux I__13800 (
            .O(N__55582),
            .I(opZ0Z_0));
    LocalMux I__13799 (
            .O(N__55579),
            .I(opZ0Z_0));
    Odrv12 I__13798 (
            .O(N__55574),
            .I(opZ0Z_0));
    Odrv4 I__13797 (
            .O(N__55567),
            .I(opZ0Z_0));
    Odrv4 I__13796 (
            .O(N__55564),
            .I(opZ0Z_0));
    Odrv4 I__13795 (
            .O(N__55555),
            .I(opZ0Z_0));
    LocalMux I__13794 (
            .O(N__55552),
            .I(opZ0Z_0));
    CascadeMux I__13793 (
            .O(N__55537),
            .I(N__55530));
    CascadeMux I__13792 (
            .O(N__55536),
            .I(N__55524));
    InMux I__13791 (
            .O(N__55535),
            .I(N__55518));
    CascadeMux I__13790 (
            .O(N__55534),
            .I(N__55514));
    InMux I__13789 (
            .O(N__55533),
            .I(N__55510));
    InMux I__13788 (
            .O(N__55530),
            .I(N__55507));
    InMux I__13787 (
            .O(N__55529),
            .I(N__55503));
    InMux I__13786 (
            .O(N__55528),
            .I(N__55500));
    InMux I__13785 (
            .O(N__55527),
            .I(N__55497));
    InMux I__13784 (
            .O(N__55524),
            .I(N__55492));
    InMux I__13783 (
            .O(N__55523),
            .I(N__55492));
    CascadeMux I__13782 (
            .O(N__55522),
            .I(N__55485));
    InMux I__13781 (
            .O(N__55521),
            .I(N__55482));
    LocalMux I__13780 (
            .O(N__55518),
            .I(N__55477));
    InMux I__13779 (
            .O(N__55517),
            .I(N__55473));
    InMux I__13778 (
            .O(N__55514),
            .I(N__55468));
    InMux I__13777 (
            .O(N__55513),
            .I(N__55468));
    LocalMux I__13776 (
            .O(N__55510),
            .I(N__55465));
    LocalMux I__13775 (
            .O(N__55507),
            .I(N__55462));
    InMux I__13774 (
            .O(N__55506),
            .I(N__55459));
    LocalMux I__13773 (
            .O(N__55503),
            .I(N__55449));
    LocalMux I__13772 (
            .O(N__55500),
            .I(N__55449));
    LocalMux I__13771 (
            .O(N__55497),
            .I(N__55449));
    LocalMux I__13770 (
            .O(N__55492),
            .I(N__55449));
    InMux I__13769 (
            .O(N__55491),
            .I(N__55441));
    InMux I__13768 (
            .O(N__55490),
            .I(N__55441));
    InMux I__13767 (
            .O(N__55489),
            .I(N__55438));
    InMux I__13766 (
            .O(N__55488),
            .I(N__55435));
    InMux I__13765 (
            .O(N__55485),
            .I(N__55431));
    LocalMux I__13764 (
            .O(N__55482),
            .I(N__55428));
    InMux I__13763 (
            .O(N__55481),
            .I(N__55423));
    InMux I__13762 (
            .O(N__55480),
            .I(N__55423));
    Span4Mux_h I__13761 (
            .O(N__55477),
            .I(N__55420));
    InMux I__13760 (
            .O(N__55476),
            .I(N__55417));
    LocalMux I__13759 (
            .O(N__55473),
            .I(N__55414));
    LocalMux I__13758 (
            .O(N__55468),
            .I(N__55411));
    Span4Mux_v I__13757 (
            .O(N__55465),
            .I(N__55404));
    Span4Mux_h I__13756 (
            .O(N__55462),
            .I(N__55404));
    LocalMux I__13755 (
            .O(N__55459),
            .I(N__55404));
    InMux I__13754 (
            .O(N__55458),
            .I(N__55401));
    Span4Mux_v I__13753 (
            .O(N__55449),
            .I(N__55396));
    InMux I__13752 (
            .O(N__55448),
            .I(N__55393));
    InMux I__13751 (
            .O(N__55447),
            .I(N__55388));
    InMux I__13750 (
            .O(N__55446),
            .I(N__55388));
    LocalMux I__13749 (
            .O(N__55441),
            .I(N__55383));
    LocalMux I__13748 (
            .O(N__55438),
            .I(N__55383));
    LocalMux I__13747 (
            .O(N__55435),
            .I(N__55378));
    InMux I__13746 (
            .O(N__55434),
            .I(N__55375));
    LocalMux I__13745 (
            .O(N__55431),
            .I(N__55366));
    Span4Mux_h I__13744 (
            .O(N__55428),
            .I(N__55366));
    LocalMux I__13743 (
            .O(N__55423),
            .I(N__55366));
    Span4Mux_v I__13742 (
            .O(N__55420),
            .I(N__55366));
    LocalMux I__13741 (
            .O(N__55417),
            .I(N__55359));
    Span4Mux_v I__13740 (
            .O(N__55414),
            .I(N__55359));
    Span4Mux_v I__13739 (
            .O(N__55411),
            .I(N__55359));
    Span4Mux_h I__13738 (
            .O(N__55404),
            .I(N__55356));
    LocalMux I__13737 (
            .O(N__55401),
            .I(N__55353));
    InMux I__13736 (
            .O(N__55400),
            .I(N__55348));
    InMux I__13735 (
            .O(N__55399),
            .I(N__55348));
    Span4Mux_h I__13734 (
            .O(N__55396),
            .I(N__55345));
    LocalMux I__13733 (
            .O(N__55393),
            .I(N__55342));
    LocalMux I__13732 (
            .O(N__55388),
            .I(N__55337));
    Span4Mux_s2_v I__13731 (
            .O(N__55383),
            .I(N__55337));
    InMux I__13730 (
            .O(N__55382),
            .I(N__55334));
    InMux I__13729 (
            .O(N__55381),
            .I(N__55331));
    Span12Mux_h I__13728 (
            .O(N__55378),
            .I(N__55328));
    LocalMux I__13727 (
            .O(N__55375),
            .I(N__55325));
    Span4Mux_v I__13726 (
            .O(N__55366),
            .I(N__55322));
    Span4Mux_h I__13725 (
            .O(N__55359),
            .I(N__55319));
    Span4Mux_v I__13724 (
            .O(N__55356),
            .I(N__55316));
    Span12Mux_s6_v I__13723 (
            .O(N__55353),
            .I(N__55311));
    LocalMux I__13722 (
            .O(N__55348),
            .I(N__55311));
    Span4Mux_h I__13721 (
            .O(N__55345),
            .I(N__55306));
    Span4Mux_h I__13720 (
            .O(N__55342),
            .I(N__55306));
    Span4Mux_h I__13719 (
            .O(N__55337),
            .I(N__55303));
    LocalMux I__13718 (
            .O(N__55334),
            .I(opZ0Z_3));
    LocalMux I__13717 (
            .O(N__55331),
            .I(opZ0Z_3));
    Odrv12 I__13716 (
            .O(N__55328),
            .I(opZ0Z_3));
    Odrv4 I__13715 (
            .O(N__55325),
            .I(opZ0Z_3));
    Odrv4 I__13714 (
            .O(N__55322),
            .I(opZ0Z_3));
    Odrv4 I__13713 (
            .O(N__55319),
            .I(opZ0Z_3));
    Odrv4 I__13712 (
            .O(N__55316),
            .I(opZ0Z_3));
    Odrv12 I__13711 (
            .O(N__55311),
            .I(opZ0Z_3));
    Odrv4 I__13710 (
            .O(N__55306),
            .I(opZ0Z_3));
    Odrv4 I__13709 (
            .O(N__55303),
            .I(opZ0Z_3));
    InMux I__13708 (
            .O(N__55282),
            .I(N__55276));
    InMux I__13707 (
            .O(N__55281),
            .I(N__55273));
    InMux I__13706 (
            .O(N__55280),
            .I(N__55269));
    InMux I__13705 (
            .O(N__55279),
            .I(N__55265));
    LocalMux I__13704 (
            .O(N__55276),
            .I(N__55256));
    LocalMux I__13703 (
            .O(N__55273),
            .I(N__55253));
    InMux I__13702 (
            .O(N__55272),
            .I(N__55250));
    LocalMux I__13701 (
            .O(N__55269),
            .I(N__55247));
    InMux I__13700 (
            .O(N__55268),
            .I(N__55244));
    LocalMux I__13699 (
            .O(N__55265),
            .I(N__55241));
    InMux I__13698 (
            .O(N__55264),
            .I(N__55238));
    InMux I__13697 (
            .O(N__55263),
            .I(N__55235));
    InMux I__13696 (
            .O(N__55262),
            .I(N__55231));
    InMux I__13695 (
            .O(N__55261),
            .I(N__55227));
    InMux I__13694 (
            .O(N__55260),
            .I(N__55224));
    CascadeMux I__13693 (
            .O(N__55259),
            .I(N__55217));
    Span4Mux_v I__13692 (
            .O(N__55256),
            .I(N__55205));
    Span4Mux_h I__13691 (
            .O(N__55253),
            .I(N__55205));
    LocalMux I__13690 (
            .O(N__55250),
            .I(N__55205));
    Span4Mux_v I__13689 (
            .O(N__55247),
            .I(N__55205));
    LocalMux I__13688 (
            .O(N__55244),
            .I(N__55205));
    Span4Mux_v I__13687 (
            .O(N__55241),
            .I(N__55202));
    LocalMux I__13686 (
            .O(N__55238),
            .I(N__55199));
    LocalMux I__13685 (
            .O(N__55235),
            .I(N__55196));
    InMux I__13684 (
            .O(N__55234),
            .I(N__55193));
    LocalMux I__13683 (
            .O(N__55231),
            .I(N__55189));
    InMux I__13682 (
            .O(N__55230),
            .I(N__55186));
    LocalMux I__13681 (
            .O(N__55227),
            .I(N__55182));
    LocalMux I__13680 (
            .O(N__55224),
            .I(N__55179));
    InMux I__13679 (
            .O(N__55223),
            .I(N__55176));
    InMux I__13678 (
            .O(N__55222),
            .I(N__55173));
    InMux I__13677 (
            .O(N__55221),
            .I(N__55169));
    InMux I__13676 (
            .O(N__55220),
            .I(N__55163));
    InMux I__13675 (
            .O(N__55217),
            .I(N__55159));
    InMux I__13674 (
            .O(N__55216),
            .I(N__55156));
    Span4Mux_v I__13673 (
            .O(N__55205),
            .I(N__55153));
    Span4Mux_h I__13672 (
            .O(N__55202),
            .I(N__55150));
    Span4Mux_h I__13671 (
            .O(N__55199),
            .I(N__55143));
    Span4Mux_h I__13670 (
            .O(N__55196),
            .I(N__55143));
    LocalMux I__13669 (
            .O(N__55193),
            .I(N__55143));
    InMux I__13668 (
            .O(N__55192),
            .I(N__55139));
    Span4Mux_v I__13667 (
            .O(N__55189),
            .I(N__55133));
    LocalMux I__13666 (
            .O(N__55186),
            .I(N__55133));
    InMux I__13665 (
            .O(N__55185),
            .I(N__55130));
    Span4Mux_v I__13664 (
            .O(N__55182),
            .I(N__55123));
    Span4Mux_h I__13663 (
            .O(N__55179),
            .I(N__55123));
    LocalMux I__13662 (
            .O(N__55176),
            .I(N__55123));
    LocalMux I__13661 (
            .O(N__55173),
            .I(N__55120));
    InMux I__13660 (
            .O(N__55172),
            .I(N__55117));
    LocalMux I__13659 (
            .O(N__55169),
            .I(N__55114));
    InMux I__13658 (
            .O(N__55168),
            .I(N__55111));
    InMux I__13657 (
            .O(N__55167),
            .I(N__55108));
    InMux I__13656 (
            .O(N__55166),
            .I(N__55105));
    LocalMux I__13655 (
            .O(N__55163),
            .I(N__55102));
    InMux I__13654 (
            .O(N__55162),
            .I(N__55099));
    LocalMux I__13653 (
            .O(N__55159),
            .I(N__55095));
    LocalMux I__13652 (
            .O(N__55156),
            .I(N__55092));
    Span4Mux_h I__13651 (
            .O(N__55153),
            .I(N__55085));
    Span4Mux_h I__13650 (
            .O(N__55150),
            .I(N__55085));
    Span4Mux_v I__13649 (
            .O(N__55143),
            .I(N__55085));
    InMux I__13648 (
            .O(N__55142),
            .I(N__55082));
    LocalMux I__13647 (
            .O(N__55139),
            .I(N__55079));
    InMux I__13646 (
            .O(N__55138),
            .I(N__55076));
    Span4Mux_v I__13645 (
            .O(N__55133),
            .I(N__55073));
    LocalMux I__13644 (
            .O(N__55130),
            .I(N__55068));
    Span4Mux_v I__13643 (
            .O(N__55123),
            .I(N__55065));
    Span4Mux_h I__13642 (
            .O(N__55120),
            .I(N__55062));
    LocalMux I__13641 (
            .O(N__55117),
            .I(N__55057));
    Span4Mux_h I__13640 (
            .O(N__55114),
            .I(N__55057));
    LocalMux I__13639 (
            .O(N__55111),
            .I(N__55048));
    LocalMux I__13638 (
            .O(N__55108),
            .I(N__55048));
    LocalMux I__13637 (
            .O(N__55105),
            .I(N__55048));
    Sp12to4 I__13636 (
            .O(N__55102),
            .I(N__55048));
    LocalMux I__13635 (
            .O(N__55099),
            .I(N__55045));
    InMux I__13634 (
            .O(N__55098),
            .I(N__55042));
    Span12Mux_s4_h I__13633 (
            .O(N__55095),
            .I(N__55035));
    Span12Mux_v I__13632 (
            .O(N__55092),
            .I(N__55035));
    Sp12to4 I__13631 (
            .O(N__55085),
            .I(N__55035));
    LocalMux I__13630 (
            .O(N__55082),
            .I(N__55030));
    Span4Mux_h I__13629 (
            .O(N__55079),
            .I(N__55030));
    LocalMux I__13628 (
            .O(N__55076),
            .I(N__55027));
    Span4Mux_h I__13627 (
            .O(N__55073),
            .I(N__55024));
    InMux I__13626 (
            .O(N__55072),
            .I(N__55021));
    InMux I__13625 (
            .O(N__55071),
            .I(N__55018));
    Span4Mux_h I__13624 (
            .O(N__55068),
            .I(N__55015));
    Span4Mux_v I__13623 (
            .O(N__55065),
            .I(N__55008));
    Span4Mux_v I__13622 (
            .O(N__55062),
            .I(N__55008));
    Span4Mux_v I__13621 (
            .O(N__55057),
            .I(N__55008));
    Span12Mux_v I__13620 (
            .O(N__55048),
            .I(N__55003));
    Span12Mux_s6_h I__13619 (
            .O(N__55045),
            .I(N__55003));
    LocalMux I__13618 (
            .O(N__55042),
            .I(N__54998));
    Span12Mux_h I__13617 (
            .O(N__55035),
            .I(N__54998));
    Span4Mux_v I__13616 (
            .O(N__55030),
            .I(N__54991));
    Span4Mux_h I__13615 (
            .O(N__55027),
            .I(N__54991));
    Span4Mux_h I__13614 (
            .O(N__55024),
            .I(N__54991));
    LocalMux I__13613 (
            .O(N__55021),
            .I(opZ0Z_1));
    LocalMux I__13612 (
            .O(N__55018),
            .I(opZ0Z_1));
    Odrv4 I__13611 (
            .O(N__55015),
            .I(opZ0Z_1));
    Odrv4 I__13610 (
            .O(N__55008),
            .I(opZ0Z_1));
    Odrv12 I__13609 (
            .O(N__55003),
            .I(opZ0Z_1));
    Odrv12 I__13608 (
            .O(N__54998),
            .I(opZ0Z_1));
    Odrv4 I__13607 (
            .O(N__54991),
            .I(opZ0Z_1));
    CascadeMux I__13606 (
            .O(N__54976),
            .I(\ALU.un1_op_1Z0Z_1_cascade_ ));
    InMux I__13605 (
            .O(N__54973),
            .I(N__54969));
    InMux I__13604 (
            .O(N__54972),
            .I(N__54966));
    LocalMux I__13603 (
            .O(N__54969),
            .I(opZ0Z_4));
    LocalMux I__13602 (
            .O(N__54966),
            .I(opZ0Z_4));
    InMux I__13601 (
            .O(N__54961),
            .I(N__54940));
    InMux I__13600 (
            .O(N__54960),
            .I(N__54940));
    InMux I__13599 (
            .O(N__54959),
            .I(N__54940));
    InMux I__13598 (
            .O(N__54958),
            .I(N__54940));
    InMux I__13597 (
            .O(N__54957),
            .I(N__54940));
    InMux I__13596 (
            .O(N__54956),
            .I(N__54940));
    InMux I__13595 (
            .O(N__54955),
            .I(N__54940));
    LocalMux I__13594 (
            .O(N__54940),
            .I(N__54937));
    Span4Mux_h I__13593 (
            .O(N__54937),
            .I(N__54933));
    InMux I__13592 (
            .O(N__54936),
            .I(N__54930));
    Odrv4 I__13591 (
            .O(N__54933),
            .I(\ALU.un1_op_1_0 ));
    LocalMux I__13590 (
            .O(N__54930),
            .I(\ALU.un1_op_1_0 ));
    InMux I__13589 (
            .O(N__54925),
            .I(N__54916));
    CascadeMux I__13588 (
            .O(N__54924),
            .I(N__54911));
    CascadeMux I__13587 (
            .O(N__54923),
            .I(N__54908));
    InMux I__13586 (
            .O(N__54922),
            .I(N__54902));
    CascadeMux I__13585 (
            .O(N__54921),
            .I(N__54895));
    CascadeMux I__13584 (
            .O(N__54920),
            .I(N__54891));
    InMux I__13583 (
            .O(N__54919),
            .I(N__54881));
    LocalMux I__13582 (
            .O(N__54916),
            .I(N__54878));
    InMux I__13581 (
            .O(N__54915),
            .I(N__54871));
    InMux I__13580 (
            .O(N__54914),
            .I(N__54871));
    InMux I__13579 (
            .O(N__54911),
            .I(N__54871));
    InMux I__13578 (
            .O(N__54908),
            .I(N__54864));
    InMux I__13577 (
            .O(N__54907),
            .I(N__54864));
    InMux I__13576 (
            .O(N__54906),
            .I(N__54864));
    InMux I__13575 (
            .O(N__54905),
            .I(N__54861));
    LocalMux I__13574 (
            .O(N__54902),
            .I(N__54855));
    InMux I__13573 (
            .O(N__54901),
            .I(N__54850));
    InMux I__13572 (
            .O(N__54900),
            .I(N__54850));
    InMux I__13571 (
            .O(N__54899),
            .I(N__54843));
    InMux I__13570 (
            .O(N__54898),
            .I(N__54843));
    InMux I__13569 (
            .O(N__54895),
            .I(N__54843));
    InMux I__13568 (
            .O(N__54894),
            .I(N__54838));
    InMux I__13567 (
            .O(N__54891),
            .I(N__54838));
    InMux I__13566 (
            .O(N__54890),
            .I(N__54830));
    CascadeMux I__13565 (
            .O(N__54889),
            .I(N__54824));
    CascadeMux I__13564 (
            .O(N__54888),
            .I(N__54818));
    CascadeMux I__13563 (
            .O(N__54887),
            .I(N__54814));
    CascadeMux I__13562 (
            .O(N__54886),
            .I(N__54807));
    CascadeMux I__13561 (
            .O(N__54885),
            .I(N__54797));
    CascadeMux I__13560 (
            .O(N__54884),
            .I(N__54792));
    LocalMux I__13559 (
            .O(N__54881),
            .I(N__54770));
    Span4Mux_h I__13558 (
            .O(N__54878),
            .I(N__54770));
    LocalMux I__13557 (
            .O(N__54871),
            .I(N__54770));
    LocalMux I__13556 (
            .O(N__54864),
            .I(N__54765));
    LocalMux I__13555 (
            .O(N__54861),
            .I(N__54765));
    InMux I__13554 (
            .O(N__54860),
            .I(N__54760));
    InMux I__13553 (
            .O(N__54859),
            .I(N__54760));
    InMux I__13552 (
            .O(N__54858),
            .I(N__54757));
    Span4Mux_v I__13551 (
            .O(N__54855),
            .I(N__54754));
    LocalMux I__13550 (
            .O(N__54850),
            .I(N__54749));
    LocalMux I__13549 (
            .O(N__54843),
            .I(N__54749));
    LocalMux I__13548 (
            .O(N__54838),
            .I(N__54746));
    InMux I__13547 (
            .O(N__54837),
            .I(N__54739));
    InMux I__13546 (
            .O(N__54836),
            .I(N__54739));
    InMux I__13545 (
            .O(N__54835),
            .I(N__54739));
    InMux I__13544 (
            .O(N__54834),
            .I(N__54734));
    InMux I__13543 (
            .O(N__54833),
            .I(N__54734));
    LocalMux I__13542 (
            .O(N__54830),
            .I(N__54731));
    InMux I__13541 (
            .O(N__54829),
            .I(N__54728));
    InMux I__13540 (
            .O(N__54828),
            .I(N__54725));
    InMux I__13539 (
            .O(N__54827),
            .I(N__54720));
    InMux I__13538 (
            .O(N__54824),
            .I(N__54720));
    CascadeMux I__13537 (
            .O(N__54823),
            .I(N__54715));
    InMux I__13536 (
            .O(N__54822),
            .I(N__54708));
    InMux I__13535 (
            .O(N__54821),
            .I(N__54708));
    InMux I__13534 (
            .O(N__54818),
            .I(N__54708));
    InMux I__13533 (
            .O(N__54817),
            .I(N__54703));
    InMux I__13532 (
            .O(N__54814),
            .I(N__54703));
    CascadeMux I__13531 (
            .O(N__54813),
            .I(N__54698));
    InMux I__13530 (
            .O(N__54812),
            .I(N__54694));
    InMux I__13529 (
            .O(N__54811),
            .I(N__54691));
    InMux I__13528 (
            .O(N__54810),
            .I(N__54686));
    InMux I__13527 (
            .O(N__54807),
            .I(N__54686));
    InMux I__13526 (
            .O(N__54806),
            .I(N__54681));
    InMux I__13525 (
            .O(N__54805),
            .I(N__54681));
    InMux I__13524 (
            .O(N__54804),
            .I(N__54672));
    InMux I__13523 (
            .O(N__54803),
            .I(N__54672));
    InMux I__13522 (
            .O(N__54802),
            .I(N__54672));
    InMux I__13521 (
            .O(N__54801),
            .I(N__54672));
    CascadeMux I__13520 (
            .O(N__54800),
            .I(N__54669));
    InMux I__13519 (
            .O(N__54797),
            .I(N__54664));
    InMux I__13518 (
            .O(N__54796),
            .I(N__54664));
    InMux I__13517 (
            .O(N__54795),
            .I(N__54659));
    InMux I__13516 (
            .O(N__54792),
            .I(N__54659));
    CascadeMux I__13515 (
            .O(N__54791),
            .I(N__54655));
    CascadeMux I__13514 (
            .O(N__54790),
            .I(N__54652));
    CascadeMux I__13513 (
            .O(N__54789),
            .I(N__54648));
    CascadeMux I__13512 (
            .O(N__54788),
            .I(N__54645));
    CascadeMux I__13511 (
            .O(N__54787),
            .I(N__54642));
    InMux I__13510 (
            .O(N__54786),
            .I(N__54633));
    InMux I__13509 (
            .O(N__54785),
            .I(N__54633));
    CascadeMux I__13508 (
            .O(N__54784),
            .I(N__54622));
    InMux I__13507 (
            .O(N__54783),
            .I(N__54619));
    InMux I__13506 (
            .O(N__54782),
            .I(N__54612));
    CascadeMux I__13505 (
            .O(N__54781),
            .I(N__54608));
    CascadeMux I__13504 (
            .O(N__54780),
            .I(N__54600));
    CascadeMux I__13503 (
            .O(N__54779),
            .I(N__54597));
    CascadeMux I__13502 (
            .O(N__54778),
            .I(N__54587));
    CascadeMux I__13501 (
            .O(N__54777),
            .I(N__54577));
    Span4Mux_v I__13500 (
            .O(N__54770),
            .I(N__54568));
    Span4Mux_v I__13499 (
            .O(N__54765),
            .I(N__54568));
    LocalMux I__13498 (
            .O(N__54760),
            .I(N__54568));
    LocalMux I__13497 (
            .O(N__54757),
            .I(N__54568));
    Span4Mux_h I__13496 (
            .O(N__54754),
            .I(N__54563));
    Span4Mux_v I__13495 (
            .O(N__54749),
            .I(N__54563));
    Span4Mux_s3_v I__13494 (
            .O(N__54746),
            .I(N__54558));
    LocalMux I__13493 (
            .O(N__54739),
            .I(N__54558));
    LocalMux I__13492 (
            .O(N__54734),
            .I(N__54547));
    Span4Mux_v I__13491 (
            .O(N__54731),
            .I(N__54547));
    LocalMux I__13490 (
            .O(N__54728),
            .I(N__54540));
    LocalMux I__13489 (
            .O(N__54725),
            .I(N__54540));
    LocalMux I__13488 (
            .O(N__54720),
            .I(N__54540));
    InMux I__13487 (
            .O(N__54719),
            .I(N__54533));
    InMux I__13486 (
            .O(N__54718),
            .I(N__54533));
    InMux I__13485 (
            .O(N__54715),
            .I(N__54533));
    LocalMux I__13484 (
            .O(N__54708),
            .I(N__54528));
    LocalMux I__13483 (
            .O(N__54703),
            .I(N__54528));
    InMux I__13482 (
            .O(N__54702),
            .I(N__54521));
    InMux I__13481 (
            .O(N__54701),
            .I(N__54521));
    InMux I__13480 (
            .O(N__54698),
            .I(N__54521));
    CascadeMux I__13479 (
            .O(N__54697),
            .I(N__54517));
    LocalMux I__13478 (
            .O(N__54694),
            .I(N__54512));
    LocalMux I__13477 (
            .O(N__54691),
            .I(N__54512));
    LocalMux I__13476 (
            .O(N__54686),
            .I(N__54509));
    LocalMux I__13475 (
            .O(N__54681),
            .I(N__54504));
    LocalMux I__13474 (
            .O(N__54672),
            .I(N__54504));
    InMux I__13473 (
            .O(N__54669),
            .I(N__54501));
    LocalMux I__13472 (
            .O(N__54664),
            .I(N__54496));
    LocalMux I__13471 (
            .O(N__54659),
            .I(N__54496));
    InMux I__13470 (
            .O(N__54658),
            .I(N__54489));
    InMux I__13469 (
            .O(N__54655),
            .I(N__54489));
    InMux I__13468 (
            .O(N__54652),
            .I(N__54489));
    InMux I__13467 (
            .O(N__54651),
            .I(N__54484));
    InMux I__13466 (
            .O(N__54648),
            .I(N__54484));
    InMux I__13465 (
            .O(N__54645),
            .I(N__54479));
    InMux I__13464 (
            .O(N__54642),
            .I(N__54479));
    InMux I__13463 (
            .O(N__54641),
            .I(N__54475));
    InMux I__13462 (
            .O(N__54640),
            .I(N__54470));
    InMux I__13461 (
            .O(N__54639),
            .I(N__54470));
    CascadeMux I__13460 (
            .O(N__54638),
            .I(N__54467));
    LocalMux I__13459 (
            .O(N__54633),
            .I(N__54464));
    InMux I__13458 (
            .O(N__54632),
            .I(N__54461));
    InMux I__13457 (
            .O(N__54631),
            .I(N__54448));
    InMux I__13456 (
            .O(N__54630),
            .I(N__54448));
    InMux I__13455 (
            .O(N__54629),
            .I(N__54448));
    InMux I__13454 (
            .O(N__54628),
            .I(N__54448));
    InMux I__13453 (
            .O(N__54627),
            .I(N__54448));
    InMux I__13452 (
            .O(N__54626),
            .I(N__54448));
    InMux I__13451 (
            .O(N__54625),
            .I(N__54442));
    InMux I__13450 (
            .O(N__54622),
            .I(N__54442));
    LocalMux I__13449 (
            .O(N__54619),
            .I(N__54439));
    InMux I__13448 (
            .O(N__54618),
            .I(N__54432));
    InMux I__13447 (
            .O(N__54617),
            .I(N__54432));
    InMux I__13446 (
            .O(N__54616),
            .I(N__54432));
    InMux I__13445 (
            .O(N__54615),
            .I(N__54429));
    LocalMux I__13444 (
            .O(N__54612),
            .I(N__54426));
    InMux I__13443 (
            .O(N__54611),
            .I(N__54423));
    InMux I__13442 (
            .O(N__54608),
            .I(N__54420));
    CascadeMux I__13441 (
            .O(N__54607),
            .I(N__54417));
    InMux I__13440 (
            .O(N__54606),
            .I(N__54414));
    InMux I__13439 (
            .O(N__54605),
            .I(N__54409));
    InMux I__13438 (
            .O(N__54604),
            .I(N__54409));
    InMux I__13437 (
            .O(N__54603),
            .I(N__54406));
    InMux I__13436 (
            .O(N__54600),
            .I(N__54403));
    InMux I__13435 (
            .O(N__54597),
            .I(N__54396));
    InMux I__13434 (
            .O(N__54596),
            .I(N__54396));
    InMux I__13433 (
            .O(N__54595),
            .I(N__54396));
    InMux I__13432 (
            .O(N__54594),
            .I(N__54393));
    InMux I__13431 (
            .O(N__54593),
            .I(N__54384));
    InMux I__13430 (
            .O(N__54592),
            .I(N__54384));
    InMux I__13429 (
            .O(N__54591),
            .I(N__54384));
    InMux I__13428 (
            .O(N__54590),
            .I(N__54384));
    InMux I__13427 (
            .O(N__54587),
            .I(N__54376));
    InMux I__13426 (
            .O(N__54586),
            .I(N__54376));
    InMux I__13425 (
            .O(N__54585),
            .I(N__54376));
    InMux I__13424 (
            .O(N__54584),
            .I(N__54373));
    InMux I__13423 (
            .O(N__54583),
            .I(N__54370));
    InMux I__13422 (
            .O(N__54582),
            .I(N__54365));
    InMux I__13421 (
            .O(N__54581),
            .I(N__54365));
    InMux I__13420 (
            .O(N__54580),
            .I(N__54362));
    InMux I__13419 (
            .O(N__54577),
            .I(N__54359));
    Span4Mux_h I__13418 (
            .O(N__54568),
            .I(N__54352));
    Span4Mux_h I__13417 (
            .O(N__54563),
            .I(N__54352));
    Span4Mux_v I__13416 (
            .O(N__54558),
            .I(N__54352));
    CascadeMux I__13415 (
            .O(N__54557),
            .I(N__54349));
    InMux I__13414 (
            .O(N__54556),
            .I(N__54346));
    InMux I__13413 (
            .O(N__54555),
            .I(N__54343));
    InMux I__13412 (
            .O(N__54554),
            .I(N__54338));
    InMux I__13411 (
            .O(N__54553),
            .I(N__54338));
    InMux I__13410 (
            .O(N__54552),
            .I(N__54335));
    Span4Mux_v I__13409 (
            .O(N__54547),
            .I(N__54328));
    Span4Mux_v I__13408 (
            .O(N__54540),
            .I(N__54328));
    LocalMux I__13407 (
            .O(N__54533),
            .I(N__54328));
    Span4Mux_h I__13406 (
            .O(N__54528),
            .I(N__54325));
    LocalMux I__13405 (
            .O(N__54521),
            .I(N__54322));
    InMux I__13404 (
            .O(N__54520),
            .I(N__54319));
    InMux I__13403 (
            .O(N__54517),
            .I(N__54316));
    Span4Mux_h I__13402 (
            .O(N__54512),
            .I(N__54301));
    Span4Mux_s2_v I__13401 (
            .O(N__54509),
            .I(N__54301));
    Span4Mux_s2_v I__13400 (
            .O(N__54504),
            .I(N__54301));
    LocalMux I__13399 (
            .O(N__54501),
            .I(N__54301));
    Span4Mux_v I__13398 (
            .O(N__54496),
            .I(N__54301));
    LocalMux I__13397 (
            .O(N__54489),
            .I(N__54301));
    LocalMux I__13396 (
            .O(N__54484),
            .I(N__54301));
    LocalMux I__13395 (
            .O(N__54479),
            .I(N__54298));
    CascadeMux I__13394 (
            .O(N__54478),
            .I(N__54295));
    LocalMux I__13393 (
            .O(N__54475),
            .I(N__54290));
    LocalMux I__13392 (
            .O(N__54470),
            .I(N__54290));
    InMux I__13391 (
            .O(N__54467),
            .I(N__54287));
    Span4Mux_s2_v I__13390 (
            .O(N__54464),
            .I(N__54280));
    LocalMux I__13389 (
            .O(N__54461),
            .I(N__54280));
    LocalMux I__13388 (
            .O(N__54448),
            .I(N__54280));
    InMux I__13387 (
            .O(N__54447),
            .I(N__54277));
    LocalMux I__13386 (
            .O(N__54442),
            .I(N__54274));
    Span4Mux_s2_v I__13385 (
            .O(N__54439),
            .I(N__54269));
    LocalMux I__13384 (
            .O(N__54432),
            .I(N__54269));
    LocalMux I__13383 (
            .O(N__54429),
            .I(N__54260));
    Span4Mux_h I__13382 (
            .O(N__54426),
            .I(N__54260));
    LocalMux I__13381 (
            .O(N__54423),
            .I(N__54260));
    LocalMux I__13380 (
            .O(N__54420),
            .I(N__54260));
    InMux I__13379 (
            .O(N__54417),
            .I(N__54257));
    LocalMux I__13378 (
            .O(N__54414),
            .I(N__54250));
    LocalMux I__13377 (
            .O(N__54409),
            .I(N__54250));
    LocalMux I__13376 (
            .O(N__54406),
            .I(N__54250));
    LocalMux I__13375 (
            .O(N__54403),
            .I(N__54247));
    LocalMux I__13374 (
            .O(N__54396),
            .I(N__54244));
    LocalMux I__13373 (
            .O(N__54393),
            .I(N__54239));
    LocalMux I__13372 (
            .O(N__54384),
            .I(N__54239));
    InMux I__13371 (
            .O(N__54383),
            .I(N__54236));
    LocalMux I__13370 (
            .O(N__54376),
            .I(N__54233));
    LocalMux I__13369 (
            .O(N__54373),
            .I(N__54230));
    LocalMux I__13368 (
            .O(N__54370),
            .I(N__54219));
    LocalMux I__13367 (
            .O(N__54365),
            .I(N__54219));
    LocalMux I__13366 (
            .O(N__54362),
            .I(N__54219));
    LocalMux I__13365 (
            .O(N__54359),
            .I(N__54219));
    Span4Mux_v I__13364 (
            .O(N__54352),
            .I(N__54219));
    InMux I__13363 (
            .O(N__54349),
            .I(N__54216));
    LocalMux I__13362 (
            .O(N__54346),
            .I(N__54212));
    LocalMux I__13361 (
            .O(N__54343),
            .I(N__54209));
    LocalMux I__13360 (
            .O(N__54338),
            .I(N__54204));
    LocalMux I__13359 (
            .O(N__54335),
            .I(N__54204));
    Span4Mux_h I__13358 (
            .O(N__54328),
            .I(N__54193));
    Span4Mux_v I__13357 (
            .O(N__54325),
            .I(N__54193));
    Span4Mux_v I__13356 (
            .O(N__54322),
            .I(N__54193));
    LocalMux I__13355 (
            .O(N__54319),
            .I(N__54193));
    LocalMux I__13354 (
            .O(N__54316),
            .I(N__54193));
    Span4Mux_h I__13353 (
            .O(N__54301),
            .I(N__54188));
    Span4Mux_s2_v I__13352 (
            .O(N__54298),
            .I(N__54188));
    InMux I__13351 (
            .O(N__54295),
            .I(N__54185));
    Span4Mux_v I__13350 (
            .O(N__54290),
            .I(N__54178));
    LocalMux I__13349 (
            .O(N__54287),
            .I(N__54178));
    Span4Mux_v I__13348 (
            .O(N__54280),
            .I(N__54178));
    LocalMux I__13347 (
            .O(N__54277),
            .I(N__54167));
    Span4Mux_h I__13346 (
            .O(N__54274),
            .I(N__54167));
    Span4Mux_v I__13345 (
            .O(N__54269),
            .I(N__54167));
    Span4Mux_v I__13344 (
            .O(N__54260),
            .I(N__54167));
    LocalMux I__13343 (
            .O(N__54257),
            .I(N__54167));
    Span4Mux_v I__13342 (
            .O(N__54250),
            .I(N__54164));
    Span4Mux_h I__13341 (
            .O(N__54247),
            .I(N__54155));
    Span4Mux_h I__13340 (
            .O(N__54244),
            .I(N__54155));
    Span4Mux_v I__13339 (
            .O(N__54239),
            .I(N__54155));
    LocalMux I__13338 (
            .O(N__54236),
            .I(N__54155));
    Span4Mux_v I__13337 (
            .O(N__54233),
            .I(N__54152));
    Span4Mux_h I__13336 (
            .O(N__54230),
            .I(N__54145));
    Span4Mux_v I__13335 (
            .O(N__54219),
            .I(N__54145));
    LocalMux I__13334 (
            .O(N__54216),
            .I(N__54145));
    CascadeMux I__13333 (
            .O(N__54215),
            .I(N__54142));
    Span4Mux_s0_v I__13332 (
            .O(N__54212),
            .I(N__54133));
    Span4Mux_h I__13331 (
            .O(N__54209),
            .I(N__54133));
    Span4Mux_h I__13330 (
            .O(N__54204),
            .I(N__54133));
    Span4Mux_h I__13329 (
            .O(N__54193),
            .I(N__54133));
    Span4Mux_h I__13328 (
            .O(N__54188),
            .I(N__54130));
    LocalMux I__13327 (
            .O(N__54185),
            .I(N__54125));
    Span4Mux_h I__13326 (
            .O(N__54178),
            .I(N__54120));
    Span4Mux_v I__13325 (
            .O(N__54167),
            .I(N__54120));
    Span4Mux_h I__13324 (
            .O(N__54164),
            .I(N__54111));
    Span4Mux_v I__13323 (
            .O(N__54155),
            .I(N__54111));
    Span4Mux_h I__13322 (
            .O(N__54152),
            .I(N__54111));
    Span4Mux_h I__13321 (
            .O(N__54145),
            .I(N__54111));
    InMux I__13320 (
            .O(N__54142),
            .I(N__54108));
    Sp12to4 I__13319 (
            .O(N__54133),
            .I(N__54105));
    Span4Mux_v I__13318 (
            .O(N__54130),
            .I(N__54102));
    InMux I__13317 (
            .O(N__54129),
            .I(N__54099));
    InMux I__13316 (
            .O(N__54128),
            .I(N__54096));
    Span4Mux_v I__13315 (
            .O(N__54125),
            .I(N__54091));
    Span4Mux_h I__13314 (
            .O(N__54120),
            .I(N__54091));
    Span4Mux_v I__13313 (
            .O(N__54111),
            .I(N__54086));
    LocalMux I__13312 (
            .O(N__54108),
            .I(N__54086));
    Span12Mux_s6_v I__13311 (
            .O(N__54105),
            .I(N__54081));
    Sp12to4 I__13310 (
            .O(N__54102),
            .I(N__54081));
    LocalMux I__13309 (
            .O(N__54099),
            .I(paramsZ0Z_1));
    LocalMux I__13308 (
            .O(N__54096),
            .I(paramsZ0Z_1));
    Odrv4 I__13307 (
            .O(N__54091),
            .I(paramsZ0Z_1));
    Odrv4 I__13306 (
            .O(N__54086),
            .I(paramsZ0Z_1));
    Odrv12 I__13305 (
            .O(N__54081),
            .I(paramsZ0Z_1));
    CascadeMux I__13304 (
            .O(N__54070),
            .I(N__54066));
    CascadeMux I__13303 (
            .O(N__54069),
            .I(N__54063));
    InMux I__13302 (
            .O(N__54066),
            .I(N__54042));
    InMux I__13301 (
            .O(N__54063),
            .I(N__54042));
    InMux I__13300 (
            .O(N__54062),
            .I(N__54033));
    CascadeMux I__13299 (
            .O(N__54061),
            .I(N__54029));
    InMux I__13298 (
            .O(N__54060),
            .I(N__54017));
    InMux I__13297 (
            .O(N__54059),
            .I(N__54014));
    InMux I__13296 (
            .O(N__54058),
            .I(N__54009));
    InMux I__13295 (
            .O(N__54057),
            .I(N__54009));
    InMux I__13294 (
            .O(N__54056),
            .I(N__54006));
    InMux I__13293 (
            .O(N__54055),
            .I(N__54003));
    InMux I__13292 (
            .O(N__54054),
            .I(N__53987));
    InMux I__13291 (
            .O(N__54053),
            .I(N__53987));
    InMux I__13290 (
            .O(N__54052),
            .I(N__53987));
    InMux I__13289 (
            .O(N__54051),
            .I(N__53987));
    InMux I__13288 (
            .O(N__54050),
            .I(N__53980));
    InMux I__13287 (
            .O(N__54049),
            .I(N__53980));
    CascadeMux I__13286 (
            .O(N__54048),
            .I(N__53977));
    CascadeMux I__13285 (
            .O(N__54047),
            .I(N__53952));
    LocalMux I__13284 (
            .O(N__54042),
            .I(N__53942));
    InMux I__13283 (
            .O(N__54041),
            .I(N__53939));
    InMux I__13282 (
            .O(N__54040),
            .I(N__53930));
    InMux I__13281 (
            .O(N__54039),
            .I(N__53930));
    InMux I__13280 (
            .O(N__54038),
            .I(N__53930));
    InMux I__13279 (
            .O(N__54037),
            .I(N__53930));
    InMux I__13278 (
            .O(N__54036),
            .I(N__53920));
    LocalMux I__13277 (
            .O(N__54033),
            .I(N__53917));
    InMux I__13276 (
            .O(N__54032),
            .I(N__53914));
    InMux I__13275 (
            .O(N__54029),
            .I(N__53908));
    InMux I__13274 (
            .O(N__54028),
            .I(N__53901));
    InMux I__13273 (
            .O(N__54027),
            .I(N__53901));
    InMux I__13272 (
            .O(N__54026),
            .I(N__53901));
    InMux I__13271 (
            .O(N__54025),
            .I(N__53890));
    InMux I__13270 (
            .O(N__54024),
            .I(N__53887));
    InMux I__13269 (
            .O(N__54023),
            .I(N__53880));
    InMux I__13268 (
            .O(N__54022),
            .I(N__53880));
    InMux I__13267 (
            .O(N__54021),
            .I(N__53875));
    InMux I__13266 (
            .O(N__54020),
            .I(N__53875));
    LocalMux I__13265 (
            .O(N__54017),
            .I(N__53864));
    LocalMux I__13264 (
            .O(N__54014),
            .I(N__53864));
    LocalMux I__13263 (
            .O(N__54009),
            .I(N__53864));
    LocalMux I__13262 (
            .O(N__54006),
            .I(N__53861));
    LocalMux I__13261 (
            .O(N__54003),
            .I(N__53858));
    InMux I__13260 (
            .O(N__54002),
            .I(N__53853));
    InMux I__13259 (
            .O(N__54001),
            .I(N__53848));
    InMux I__13258 (
            .O(N__54000),
            .I(N__53848));
    InMux I__13257 (
            .O(N__53999),
            .I(N__53843));
    InMux I__13256 (
            .O(N__53998),
            .I(N__53843));
    InMux I__13255 (
            .O(N__53997),
            .I(N__53838));
    InMux I__13254 (
            .O(N__53996),
            .I(N__53838));
    LocalMux I__13253 (
            .O(N__53987),
            .I(N__53835));
    InMux I__13252 (
            .O(N__53986),
            .I(N__53832));
    InMux I__13251 (
            .O(N__53985),
            .I(N__53829));
    LocalMux I__13250 (
            .O(N__53980),
            .I(N__53826));
    InMux I__13249 (
            .O(N__53977),
            .I(N__53823));
    InMux I__13248 (
            .O(N__53976),
            .I(N__53816));
    InMux I__13247 (
            .O(N__53975),
            .I(N__53816));
    InMux I__13246 (
            .O(N__53974),
            .I(N__53816));
    InMux I__13245 (
            .O(N__53973),
            .I(N__53813));
    InMux I__13244 (
            .O(N__53972),
            .I(N__53808));
    InMux I__13243 (
            .O(N__53971),
            .I(N__53799));
    InMux I__13242 (
            .O(N__53970),
            .I(N__53799));
    InMux I__13241 (
            .O(N__53969),
            .I(N__53792));
    InMux I__13240 (
            .O(N__53968),
            .I(N__53792));
    InMux I__13239 (
            .O(N__53967),
            .I(N__53792));
    InMux I__13238 (
            .O(N__53966),
            .I(N__53783));
    InMux I__13237 (
            .O(N__53965),
            .I(N__53783));
    InMux I__13236 (
            .O(N__53964),
            .I(N__53783));
    InMux I__13235 (
            .O(N__53963),
            .I(N__53783));
    InMux I__13234 (
            .O(N__53962),
            .I(N__53771));
    InMux I__13233 (
            .O(N__53961),
            .I(N__53771));
    InMux I__13232 (
            .O(N__53960),
            .I(N__53771));
    InMux I__13231 (
            .O(N__53959),
            .I(N__53766));
    InMux I__13230 (
            .O(N__53958),
            .I(N__53766));
    InMux I__13229 (
            .O(N__53957),
            .I(N__53763));
    InMux I__13228 (
            .O(N__53956),
            .I(N__53760));
    InMux I__13227 (
            .O(N__53955),
            .I(N__53754));
    InMux I__13226 (
            .O(N__53952),
            .I(N__53748));
    InMux I__13225 (
            .O(N__53951),
            .I(N__53748));
    InMux I__13224 (
            .O(N__53950),
            .I(N__53743));
    InMux I__13223 (
            .O(N__53949),
            .I(N__53743));
    InMux I__13222 (
            .O(N__53948),
            .I(N__53735));
    InMux I__13221 (
            .O(N__53947),
            .I(N__53735));
    InMux I__13220 (
            .O(N__53946),
            .I(N__53735));
    InMux I__13219 (
            .O(N__53945),
            .I(N__53732));
    Span4Mux_s2_v I__13218 (
            .O(N__53942),
            .I(N__53725));
    LocalMux I__13217 (
            .O(N__53939),
            .I(N__53725));
    LocalMux I__13216 (
            .O(N__53930),
            .I(N__53725));
    InMux I__13215 (
            .O(N__53929),
            .I(N__53718));
    InMux I__13214 (
            .O(N__53928),
            .I(N__53718));
    InMux I__13213 (
            .O(N__53927),
            .I(N__53718));
    InMux I__13212 (
            .O(N__53926),
            .I(N__53709));
    InMux I__13211 (
            .O(N__53925),
            .I(N__53709));
    InMux I__13210 (
            .O(N__53924),
            .I(N__53709));
    InMux I__13209 (
            .O(N__53923),
            .I(N__53709));
    LocalMux I__13208 (
            .O(N__53920),
            .I(N__53702));
    Span4Mux_v I__13207 (
            .O(N__53917),
            .I(N__53702));
    LocalMux I__13206 (
            .O(N__53914),
            .I(N__53702));
    InMux I__13205 (
            .O(N__53913),
            .I(N__53695));
    InMux I__13204 (
            .O(N__53912),
            .I(N__53695));
    InMux I__13203 (
            .O(N__53911),
            .I(N__53695));
    LocalMux I__13202 (
            .O(N__53908),
            .I(N__53690));
    LocalMux I__13201 (
            .O(N__53901),
            .I(N__53690));
    InMux I__13200 (
            .O(N__53900),
            .I(N__53687));
    CascadeMux I__13199 (
            .O(N__53899),
            .I(N__53682));
    InMux I__13198 (
            .O(N__53898),
            .I(N__53677));
    InMux I__13197 (
            .O(N__53897),
            .I(N__53672));
    InMux I__13196 (
            .O(N__53896),
            .I(N__53669));
    InMux I__13195 (
            .O(N__53895),
            .I(N__53662));
    InMux I__13194 (
            .O(N__53894),
            .I(N__53662));
    InMux I__13193 (
            .O(N__53893),
            .I(N__53662));
    LocalMux I__13192 (
            .O(N__53890),
            .I(N__53657));
    LocalMux I__13191 (
            .O(N__53887),
            .I(N__53657));
    InMux I__13190 (
            .O(N__53886),
            .I(N__53652));
    InMux I__13189 (
            .O(N__53885),
            .I(N__53652));
    LocalMux I__13188 (
            .O(N__53880),
            .I(N__53647));
    LocalMux I__13187 (
            .O(N__53875),
            .I(N__53647));
    InMux I__13186 (
            .O(N__53874),
            .I(N__53641));
    InMux I__13185 (
            .O(N__53873),
            .I(N__53636));
    InMux I__13184 (
            .O(N__53872),
            .I(N__53636));
    InMux I__13183 (
            .O(N__53871),
            .I(N__53633));
    Span4Mux_v I__13182 (
            .O(N__53864),
            .I(N__53630));
    Span4Mux_s3_v I__13181 (
            .O(N__53861),
            .I(N__53625));
    Span4Mux_h I__13180 (
            .O(N__53858),
            .I(N__53625));
    InMux I__13179 (
            .O(N__53857),
            .I(N__53620));
    InMux I__13178 (
            .O(N__53856),
            .I(N__53620));
    LocalMux I__13177 (
            .O(N__53853),
            .I(N__53613));
    LocalMux I__13176 (
            .O(N__53848),
            .I(N__53613));
    LocalMux I__13175 (
            .O(N__53843),
            .I(N__53613));
    LocalMux I__13174 (
            .O(N__53838),
            .I(N__53610));
    Span4Mux_h I__13173 (
            .O(N__53835),
            .I(N__53607));
    LocalMux I__13172 (
            .O(N__53832),
            .I(N__53594));
    LocalMux I__13171 (
            .O(N__53829),
            .I(N__53594));
    Span4Mux_h I__13170 (
            .O(N__53826),
            .I(N__53594));
    LocalMux I__13169 (
            .O(N__53823),
            .I(N__53594));
    LocalMux I__13168 (
            .O(N__53816),
            .I(N__53594));
    LocalMux I__13167 (
            .O(N__53813),
            .I(N__53594));
    CascadeMux I__13166 (
            .O(N__53812),
            .I(N__53591));
    InMux I__13165 (
            .O(N__53811),
            .I(N__53587));
    LocalMux I__13164 (
            .O(N__53808),
            .I(N__53584));
    InMux I__13163 (
            .O(N__53807),
            .I(N__53579));
    InMux I__13162 (
            .O(N__53806),
            .I(N__53579));
    InMux I__13161 (
            .O(N__53805),
            .I(N__53576));
    InMux I__13160 (
            .O(N__53804),
            .I(N__53573));
    LocalMux I__13159 (
            .O(N__53799),
            .I(N__53570));
    LocalMux I__13158 (
            .O(N__53792),
            .I(N__53565));
    LocalMux I__13157 (
            .O(N__53783),
            .I(N__53565));
    InMux I__13156 (
            .O(N__53782),
            .I(N__53562));
    InMux I__13155 (
            .O(N__53781),
            .I(N__53559));
    InMux I__13154 (
            .O(N__53780),
            .I(N__53552));
    InMux I__13153 (
            .O(N__53779),
            .I(N__53552));
    InMux I__13152 (
            .O(N__53778),
            .I(N__53552));
    LocalMux I__13151 (
            .O(N__53771),
            .I(N__53543));
    LocalMux I__13150 (
            .O(N__53766),
            .I(N__53543));
    LocalMux I__13149 (
            .O(N__53763),
            .I(N__53543));
    LocalMux I__13148 (
            .O(N__53760),
            .I(N__53543));
    InMux I__13147 (
            .O(N__53759),
            .I(N__53540));
    InMux I__13146 (
            .O(N__53758),
            .I(N__53535));
    InMux I__13145 (
            .O(N__53757),
            .I(N__53535));
    LocalMux I__13144 (
            .O(N__53754),
            .I(N__53532));
    InMux I__13143 (
            .O(N__53753),
            .I(N__53529));
    LocalMux I__13142 (
            .O(N__53748),
            .I(N__53526));
    LocalMux I__13141 (
            .O(N__53743),
            .I(N__53523));
    InMux I__13140 (
            .O(N__53742),
            .I(N__53520));
    LocalMux I__13139 (
            .O(N__53735),
            .I(N__53517));
    LocalMux I__13138 (
            .O(N__53732),
            .I(N__53513));
    Span4Mux_v I__13137 (
            .O(N__53725),
            .I(N__53510));
    LocalMux I__13136 (
            .O(N__53718),
            .I(N__53505));
    LocalMux I__13135 (
            .O(N__53709),
            .I(N__53505));
    Span4Mux_s2_v I__13134 (
            .O(N__53702),
            .I(N__53500));
    LocalMux I__13133 (
            .O(N__53695),
            .I(N__53500));
    Span4Mux_v I__13132 (
            .O(N__53690),
            .I(N__53495));
    LocalMux I__13131 (
            .O(N__53687),
            .I(N__53495));
    InMux I__13130 (
            .O(N__53686),
            .I(N__53486));
    InMux I__13129 (
            .O(N__53685),
            .I(N__53486));
    InMux I__13128 (
            .O(N__53682),
            .I(N__53486));
    InMux I__13127 (
            .O(N__53681),
            .I(N__53486));
    InMux I__13126 (
            .O(N__53680),
            .I(N__53483));
    LocalMux I__13125 (
            .O(N__53677),
            .I(N__53480));
    InMux I__13124 (
            .O(N__53676),
            .I(N__53475));
    InMux I__13123 (
            .O(N__53675),
            .I(N__53475));
    LocalMux I__13122 (
            .O(N__53672),
            .I(N__53466));
    LocalMux I__13121 (
            .O(N__53669),
            .I(N__53466));
    LocalMux I__13120 (
            .O(N__53662),
            .I(N__53466));
    Span4Mux_v I__13119 (
            .O(N__53657),
            .I(N__53466));
    LocalMux I__13118 (
            .O(N__53652),
            .I(N__53461));
    Span4Mux_v I__13117 (
            .O(N__53647),
            .I(N__53461));
    InMux I__13116 (
            .O(N__53646),
            .I(N__53454));
    InMux I__13115 (
            .O(N__53645),
            .I(N__53454));
    InMux I__13114 (
            .O(N__53644),
            .I(N__53454));
    LocalMux I__13113 (
            .O(N__53641),
            .I(N__53447));
    LocalMux I__13112 (
            .O(N__53636),
            .I(N__53447));
    LocalMux I__13111 (
            .O(N__53633),
            .I(N__53447));
    Span4Mux_h I__13110 (
            .O(N__53630),
            .I(N__53442));
    Span4Mux_v I__13109 (
            .O(N__53625),
            .I(N__53442));
    LocalMux I__13108 (
            .O(N__53620),
            .I(N__53435));
    Span4Mux_h I__13107 (
            .O(N__53613),
            .I(N__53435));
    Span4Mux_h I__13106 (
            .O(N__53610),
            .I(N__53435));
    Span4Mux_v I__13105 (
            .O(N__53607),
            .I(N__53430));
    Span4Mux_v I__13104 (
            .O(N__53594),
            .I(N__53430));
    InMux I__13103 (
            .O(N__53591),
            .I(N__53425));
    InMux I__13102 (
            .O(N__53590),
            .I(N__53425));
    LocalMux I__13101 (
            .O(N__53587),
            .I(N__53422));
    Span4Mux_v I__13100 (
            .O(N__53584),
            .I(N__53418));
    LocalMux I__13099 (
            .O(N__53579),
            .I(N__53415));
    LocalMux I__13098 (
            .O(N__53576),
            .I(N__53412));
    LocalMux I__13097 (
            .O(N__53573),
            .I(N__53401));
    Span4Mux_h I__13096 (
            .O(N__53570),
            .I(N__53401));
    Span4Mux_s2_v I__13095 (
            .O(N__53565),
            .I(N__53401));
    LocalMux I__13094 (
            .O(N__53562),
            .I(N__53401));
    LocalMux I__13093 (
            .O(N__53559),
            .I(N__53401));
    LocalMux I__13092 (
            .O(N__53552),
            .I(N__53396));
    Span4Mux_v I__13091 (
            .O(N__53543),
            .I(N__53396));
    LocalMux I__13090 (
            .O(N__53540),
            .I(N__53387));
    LocalMux I__13089 (
            .O(N__53535),
            .I(N__53387));
    Span4Mux_h I__13088 (
            .O(N__53532),
            .I(N__53387));
    LocalMux I__13087 (
            .O(N__53529),
            .I(N__53387));
    Span4Mux_s2_v I__13086 (
            .O(N__53526),
            .I(N__53380));
    Span4Mux_s2_v I__13085 (
            .O(N__53523),
            .I(N__53380));
    LocalMux I__13084 (
            .O(N__53520),
            .I(N__53380));
    Span4Mux_s2_v I__13083 (
            .O(N__53517),
            .I(N__53377));
    InMux I__13082 (
            .O(N__53516),
            .I(N__53374));
    Span4Mux_v I__13081 (
            .O(N__53513),
            .I(N__53365));
    Span4Mux_h I__13080 (
            .O(N__53510),
            .I(N__53365));
    Span4Mux_v I__13079 (
            .O(N__53505),
            .I(N__53365));
    Span4Mux_v I__13078 (
            .O(N__53500),
            .I(N__53365));
    Span4Mux_h I__13077 (
            .O(N__53495),
            .I(N__53358));
    LocalMux I__13076 (
            .O(N__53486),
            .I(N__53358));
    LocalMux I__13075 (
            .O(N__53483),
            .I(N__53358));
    Span4Mux_h I__13074 (
            .O(N__53480),
            .I(N__53351));
    LocalMux I__13073 (
            .O(N__53475),
            .I(N__53351));
    Span4Mux_v I__13072 (
            .O(N__53466),
            .I(N__53342));
    Span4Mux_h I__13071 (
            .O(N__53461),
            .I(N__53342));
    LocalMux I__13070 (
            .O(N__53454),
            .I(N__53342));
    Span4Mux_v I__13069 (
            .O(N__53447),
            .I(N__53342));
    Span4Mux_h I__13068 (
            .O(N__53442),
            .I(N__53335));
    Span4Mux_h I__13067 (
            .O(N__53435),
            .I(N__53335));
    Span4Mux_h I__13066 (
            .O(N__53430),
            .I(N__53335));
    LocalMux I__13065 (
            .O(N__53425),
            .I(N__53330));
    Span4Mux_v I__13064 (
            .O(N__53422),
            .I(N__53330));
    InMux I__13063 (
            .O(N__53421),
            .I(N__53327));
    Span4Mux_h I__13062 (
            .O(N__53418),
            .I(N__53320));
    Span4Mux_v I__13061 (
            .O(N__53415),
            .I(N__53320));
    Span4Mux_v I__13060 (
            .O(N__53412),
            .I(N__53320));
    Span4Mux_h I__13059 (
            .O(N__53401),
            .I(N__53317));
    Span4Mux_h I__13058 (
            .O(N__53396),
            .I(N__53310));
    Span4Mux_v I__13057 (
            .O(N__53387),
            .I(N__53310));
    Span4Mux_v I__13056 (
            .O(N__53380),
            .I(N__53310));
    Span4Mux_h I__13055 (
            .O(N__53377),
            .I(N__53305));
    LocalMux I__13054 (
            .O(N__53374),
            .I(N__53305));
    Span4Mux_h I__13053 (
            .O(N__53365),
            .I(N__53302));
    Span4Mux_v I__13052 (
            .O(N__53358),
            .I(N__53299));
    InMux I__13051 (
            .O(N__53357),
            .I(N__53294));
    InMux I__13050 (
            .O(N__53356),
            .I(N__53294));
    Span4Mux_v I__13049 (
            .O(N__53351),
            .I(N__53289));
    Span4Mux_h I__13048 (
            .O(N__53342),
            .I(N__53289));
    Span4Mux_v I__13047 (
            .O(N__53335),
            .I(N__53282));
    Span4Mux_s3_v I__13046 (
            .O(N__53330),
            .I(N__53282));
    LocalMux I__13045 (
            .O(N__53327),
            .I(N__53282));
    Span4Mux_h I__13044 (
            .O(N__53320),
            .I(N__53275));
    Span4Mux_v I__13043 (
            .O(N__53317),
            .I(N__53275));
    Span4Mux_v I__13042 (
            .O(N__53310),
            .I(N__53275));
    Span4Mux_v I__13041 (
            .O(N__53305),
            .I(N__53268));
    Span4Mux_h I__13040 (
            .O(N__53302),
            .I(N__53268));
    Span4Mux_v I__13039 (
            .O(N__53299),
            .I(N__53268));
    LocalMux I__13038 (
            .O(N__53294),
            .I(paramsZ0Z_0));
    Odrv4 I__13037 (
            .O(N__53289),
            .I(paramsZ0Z_0));
    Odrv4 I__13036 (
            .O(N__53282),
            .I(paramsZ0Z_0));
    Odrv4 I__13035 (
            .O(N__53275),
            .I(paramsZ0Z_0));
    Odrv4 I__13034 (
            .O(N__53268),
            .I(paramsZ0Z_0));
    CascadeMux I__13033 (
            .O(N__53257),
            .I(N__53251));
    InMux I__13032 (
            .O(N__53256),
            .I(N__53247));
    InMux I__13031 (
            .O(N__53255),
            .I(N__53244));
    InMux I__13030 (
            .O(N__53254),
            .I(N__53233));
    InMux I__13029 (
            .O(N__53251),
            .I(N__53225));
    CascadeMux I__13028 (
            .O(N__53250),
            .I(N__53209));
    LocalMux I__13027 (
            .O(N__53247),
            .I(N__53200));
    LocalMux I__13026 (
            .O(N__53244),
            .I(N__53200));
    CascadeMux I__13025 (
            .O(N__53243),
            .I(N__53197));
    CascadeMux I__13024 (
            .O(N__53242),
            .I(N__53190));
    CascadeMux I__13023 (
            .O(N__53241),
            .I(N__53187));
    CascadeMux I__13022 (
            .O(N__53240),
            .I(N__53184));
    CascadeMux I__13021 (
            .O(N__53239),
            .I(N__53177));
    InMux I__13020 (
            .O(N__53238),
            .I(N__53170));
    InMux I__13019 (
            .O(N__53237),
            .I(N__53170));
    CascadeMux I__13018 (
            .O(N__53236),
            .I(N__53155));
    LocalMux I__13017 (
            .O(N__53233),
            .I(N__53149));
    CascadeMux I__13016 (
            .O(N__53232),
            .I(N__53146));
    CascadeMux I__13015 (
            .O(N__53231),
            .I(N__53140));
    CascadeMux I__13014 (
            .O(N__53230),
            .I(N__53136));
    CascadeMux I__13013 (
            .O(N__53229),
            .I(N__53131));
    CascadeMux I__13012 (
            .O(N__53228),
            .I(N__53126));
    LocalMux I__13011 (
            .O(N__53225),
            .I(N__53123));
    CascadeMux I__13010 (
            .O(N__53224),
            .I(N__53115));
    CascadeMux I__13009 (
            .O(N__53223),
            .I(N__53111));
    CascadeMux I__13008 (
            .O(N__53222),
            .I(N__53108));
    CascadeMux I__13007 (
            .O(N__53221),
            .I(N__53105));
    CascadeMux I__13006 (
            .O(N__53220),
            .I(N__53099));
    CascadeMux I__13005 (
            .O(N__53219),
            .I(N__53095));
    CascadeMux I__13004 (
            .O(N__53218),
            .I(N__53092));
    CascadeMux I__13003 (
            .O(N__53217),
            .I(N__53087));
    CascadeMux I__13002 (
            .O(N__53216),
            .I(N__53084));
    CascadeMux I__13001 (
            .O(N__53215),
            .I(N__53081));
    CascadeMux I__13000 (
            .O(N__53214),
            .I(N__53077));
    CascadeMux I__12999 (
            .O(N__53213),
            .I(N__53074));
    InMux I__12998 (
            .O(N__53212),
            .I(N__53069));
    InMux I__12997 (
            .O(N__53209),
            .I(N__53069));
    CascadeMux I__12996 (
            .O(N__53208),
            .I(N__53065));
    CascadeMux I__12995 (
            .O(N__53207),
            .I(N__53061));
    CascadeMux I__12994 (
            .O(N__53206),
            .I(N__53058));
    CascadeMux I__12993 (
            .O(N__53205),
            .I(N__53055));
    Span4Mux_h I__12992 (
            .O(N__53200),
            .I(N__53052));
    InMux I__12991 (
            .O(N__53197),
            .I(N__53045));
    InMux I__12990 (
            .O(N__53196),
            .I(N__53045));
    InMux I__12989 (
            .O(N__53195),
            .I(N__53045));
    InMux I__12988 (
            .O(N__53194),
            .I(N__53034));
    InMux I__12987 (
            .O(N__53193),
            .I(N__53034));
    InMux I__12986 (
            .O(N__53190),
            .I(N__53034));
    InMux I__12985 (
            .O(N__53187),
            .I(N__53034));
    InMux I__12984 (
            .O(N__53184),
            .I(N__53034));
    CascadeMux I__12983 (
            .O(N__53183),
            .I(N__53031));
    CascadeMux I__12982 (
            .O(N__53182),
            .I(N__53028));
    CascadeMux I__12981 (
            .O(N__53181),
            .I(N__53025));
    InMux I__12980 (
            .O(N__53180),
            .I(N__53018));
    InMux I__12979 (
            .O(N__53177),
            .I(N__53018));
    InMux I__12978 (
            .O(N__53176),
            .I(N__53018));
    InMux I__12977 (
            .O(N__53175),
            .I(N__53015));
    LocalMux I__12976 (
            .O(N__53170),
            .I(N__53011));
    CascadeMux I__12975 (
            .O(N__53169),
            .I(N__53008));
    CascadeMux I__12974 (
            .O(N__53168),
            .I(N__53005));
    CascadeMux I__12973 (
            .O(N__53167),
            .I(N__53000));
    CascadeMux I__12972 (
            .O(N__53166),
            .I(N__52997));
    CascadeMux I__12971 (
            .O(N__53165),
            .I(N__52993));
    CascadeMux I__12970 (
            .O(N__53164),
            .I(N__52989));
    CascadeMux I__12969 (
            .O(N__53163),
            .I(N__52986));
    CascadeMux I__12968 (
            .O(N__53162),
            .I(N__52979));
    CascadeMux I__12967 (
            .O(N__53161),
            .I(N__52976));
    CascadeMux I__12966 (
            .O(N__53160),
            .I(N__52973));
    InMux I__12965 (
            .O(N__53159),
            .I(N__52967));
    CascadeMux I__12964 (
            .O(N__53158),
            .I(N__52964));
    InMux I__12963 (
            .O(N__53155),
            .I(N__52960));
    CascadeMux I__12962 (
            .O(N__53154),
            .I(N__52957));
    CascadeMux I__12961 (
            .O(N__53153),
            .I(N__52954));
    CascadeMux I__12960 (
            .O(N__53152),
            .I(N__52951));
    Span4Mux_s3_h I__12959 (
            .O(N__53149),
            .I(N__52948));
    InMux I__12958 (
            .O(N__53146),
            .I(N__52945));
    InMux I__12957 (
            .O(N__53145),
            .I(N__52942));
    CascadeMux I__12956 (
            .O(N__53144),
            .I(N__52934));
    CascadeMux I__12955 (
            .O(N__53143),
            .I(N__52931));
    InMux I__12954 (
            .O(N__53140),
            .I(N__52928));
    InMux I__12953 (
            .O(N__53139),
            .I(N__52925));
    InMux I__12952 (
            .O(N__53136),
            .I(N__52922));
    InMux I__12951 (
            .O(N__53135),
            .I(N__52915));
    InMux I__12950 (
            .O(N__53134),
            .I(N__52915));
    InMux I__12949 (
            .O(N__53131),
            .I(N__52915));
    CascadeMux I__12948 (
            .O(N__53130),
            .I(N__52912));
    CascadeMux I__12947 (
            .O(N__53129),
            .I(N__52909));
    InMux I__12946 (
            .O(N__53126),
            .I(N__52906));
    Span4Mux_s2_v I__12945 (
            .O(N__53123),
            .I(N__52903));
    CascadeMux I__12944 (
            .O(N__53122),
            .I(N__52900));
    CascadeMux I__12943 (
            .O(N__53121),
            .I(N__52897));
    CascadeMux I__12942 (
            .O(N__53120),
            .I(N__52894));
    InMux I__12941 (
            .O(N__53119),
            .I(N__52890));
    InMux I__12940 (
            .O(N__53118),
            .I(N__52887));
    InMux I__12939 (
            .O(N__53115),
            .I(N__52884));
    CascadeMux I__12938 (
            .O(N__53114),
            .I(N__52881));
    InMux I__12937 (
            .O(N__53111),
            .I(N__52876));
    InMux I__12936 (
            .O(N__53108),
            .I(N__52873));
    InMux I__12935 (
            .O(N__53105),
            .I(N__52870));
    CascadeMux I__12934 (
            .O(N__53104),
            .I(N__52867));
    CascadeMux I__12933 (
            .O(N__53103),
            .I(N__52864));
    CascadeMux I__12932 (
            .O(N__53102),
            .I(N__52861));
    InMux I__12931 (
            .O(N__53099),
            .I(N__52858));
    InMux I__12930 (
            .O(N__53098),
            .I(N__52855));
    InMux I__12929 (
            .O(N__53095),
            .I(N__52848));
    InMux I__12928 (
            .O(N__53092),
            .I(N__52848));
    InMux I__12927 (
            .O(N__53091),
            .I(N__52848));
    InMux I__12926 (
            .O(N__53090),
            .I(N__52841));
    InMux I__12925 (
            .O(N__53087),
            .I(N__52841));
    InMux I__12924 (
            .O(N__53084),
            .I(N__52841));
    InMux I__12923 (
            .O(N__53081),
            .I(N__52838));
    InMux I__12922 (
            .O(N__53080),
            .I(N__52833));
    InMux I__12921 (
            .O(N__53077),
            .I(N__52833));
    InMux I__12920 (
            .O(N__53074),
            .I(N__52830));
    LocalMux I__12919 (
            .O(N__53069),
            .I(N__52827));
    CascadeMux I__12918 (
            .O(N__53068),
            .I(N__52824));
    InMux I__12917 (
            .O(N__53065),
            .I(N__52821));
    InMux I__12916 (
            .O(N__53064),
            .I(N__52816));
    InMux I__12915 (
            .O(N__53061),
            .I(N__52811));
    InMux I__12914 (
            .O(N__53058),
            .I(N__52811));
    InMux I__12913 (
            .O(N__53055),
            .I(N__52808));
    Span4Mux_h I__12912 (
            .O(N__53052),
            .I(N__52803));
    LocalMux I__12911 (
            .O(N__53045),
            .I(N__52803));
    LocalMux I__12910 (
            .O(N__53034),
            .I(N__52800));
    InMux I__12909 (
            .O(N__53031),
            .I(N__52793));
    InMux I__12908 (
            .O(N__53028),
            .I(N__52793));
    InMux I__12907 (
            .O(N__53025),
            .I(N__52793));
    LocalMux I__12906 (
            .O(N__53018),
            .I(N__52788));
    LocalMux I__12905 (
            .O(N__53015),
            .I(N__52788));
    InMux I__12904 (
            .O(N__53014),
            .I(N__52785));
    Span4Mux_s2_h I__12903 (
            .O(N__53011),
            .I(N__52782));
    InMux I__12902 (
            .O(N__53008),
            .I(N__52775));
    InMux I__12901 (
            .O(N__53005),
            .I(N__52775));
    InMux I__12900 (
            .O(N__53004),
            .I(N__52775));
    InMux I__12899 (
            .O(N__53003),
            .I(N__52766));
    InMux I__12898 (
            .O(N__53000),
            .I(N__52766));
    InMux I__12897 (
            .O(N__52997),
            .I(N__52766));
    InMux I__12896 (
            .O(N__52996),
            .I(N__52766));
    InMux I__12895 (
            .O(N__52993),
            .I(N__52759));
    InMux I__12894 (
            .O(N__52992),
            .I(N__52759));
    InMux I__12893 (
            .O(N__52989),
            .I(N__52759));
    InMux I__12892 (
            .O(N__52986),
            .I(N__52742));
    InMux I__12891 (
            .O(N__52985),
            .I(N__52742));
    InMux I__12890 (
            .O(N__52984),
            .I(N__52742));
    InMux I__12889 (
            .O(N__52983),
            .I(N__52742));
    InMux I__12888 (
            .O(N__52982),
            .I(N__52742));
    InMux I__12887 (
            .O(N__52979),
            .I(N__52742));
    InMux I__12886 (
            .O(N__52976),
            .I(N__52742));
    InMux I__12885 (
            .O(N__52973),
            .I(N__52742));
    CascadeMux I__12884 (
            .O(N__52972),
            .I(N__52738));
    CascadeMux I__12883 (
            .O(N__52971),
            .I(N__52735));
    CascadeMux I__12882 (
            .O(N__52970),
            .I(N__52732));
    LocalMux I__12881 (
            .O(N__52967),
            .I(N__52729));
    InMux I__12880 (
            .O(N__52964),
            .I(N__52726));
    CascadeMux I__12879 (
            .O(N__52963),
            .I(N__52723));
    LocalMux I__12878 (
            .O(N__52960),
            .I(N__52720));
    InMux I__12877 (
            .O(N__52957),
            .I(N__52713));
    InMux I__12876 (
            .O(N__52954),
            .I(N__52713));
    InMux I__12875 (
            .O(N__52951),
            .I(N__52710));
    Span4Mux_v I__12874 (
            .O(N__52948),
            .I(N__52703));
    LocalMux I__12873 (
            .O(N__52945),
            .I(N__52703));
    LocalMux I__12872 (
            .O(N__52942),
            .I(N__52703));
    CascadeMux I__12871 (
            .O(N__52941),
            .I(N__52700));
    CascadeMux I__12870 (
            .O(N__52940),
            .I(N__52697));
    CascadeMux I__12869 (
            .O(N__52939),
            .I(N__52694));
    CascadeMux I__12868 (
            .O(N__52938),
            .I(N__52691));
    InMux I__12867 (
            .O(N__52937),
            .I(N__52688));
    InMux I__12866 (
            .O(N__52934),
            .I(N__52683));
    InMux I__12865 (
            .O(N__52931),
            .I(N__52683));
    LocalMux I__12864 (
            .O(N__52928),
            .I(N__52674));
    LocalMux I__12863 (
            .O(N__52925),
            .I(N__52674));
    LocalMux I__12862 (
            .O(N__52922),
            .I(N__52674));
    LocalMux I__12861 (
            .O(N__52915),
            .I(N__52674));
    InMux I__12860 (
            .O(N__52912),
            .I(N__52669));
    InMux I__12859 (
            .O(N__52909),
            .I(N__52669));
    LocalMux I__12858 (
            .O(N__52906),
            .I(N__52664));
    Span4Mux_h I__12857 (
            .O(N__52903),
            .I(N__52664));
    InMux I__12856 (
            .O(N__52900),
            .I(N__52657));
    InMux I__12855 (
            .O(N__52897),
            .I(N__52657));
    InMux I__12854 (
            .O(N__52894),
            .I(N__52657));
    InMux I__12853 (
            .O(N__52893),
            .I(N__52654));
    LocalMux I__12852 (
            .O(N__52890),
            .I(N__52647));
    LocalMux I__12851 (
            .O(N__52887),
            .I(N__52647));
    LocalMux I__12850 (
            .O(N__52884),
            .I(N__52647));
    InMux I__12849 (
            .O(N__52881),
            .I(N__52640));
    InMux I__12848 (
            .O(N__52880),
            .I(N__52640));
    InMux I__12847 (
            .O(N__52879),
            .I(N__52640));
    LocalMux I__12846 (
            .O(N__52876),
            .I(N__52633));
    LocalMux I__12845 (
            .O(N__52873),
            .I(N__52633));
    LocalMux I__12844 (
            .O(N__52870),
            .I(N__52633));
    InMux I__12843 (
            .O(N__52867),
            .I(N__52630));
    InMux I__12842 (
            .O(N__52864),
            .I(N__52625));
    InMux I__12841 (
            .O(N__52861),
            .I(N__52625));
    LocalMux I__12840 (
            .O(N__52858),
            .I(N__52620));
    LocalMux I__12839 (
            .O(N__52855),
            .I(N__52620));
    LocalMux I__12838 (
            .O(N__52848),
            .I(N__52617));
    LocalMux I__12837 (
            .O(N__52841),
            .I(N__52610));
    LocalMux I__12836 (
            .O(N__52838),
            .I(N__52610));
    LocalMux I__12835 (
            .O(N__52833),
            .I(N__52610));
    LocalMux I__12834 (
            .O(N__52830),
            .I(N__52605));
    Span4Mux_s2_v I__12833 (
            .O(N__52827),
            .I(N__52605));
    InMux I__12832 (
            .O(N__52824),
            .I(N__52602));
    LocalMux I__12831 (
            .O(N__52821),
            .I(N__52599));
    InMux I__12830 (
            .O(N__52820),
            .I(N__52593));
    InMux I__12829 (
            .O(N__52819),
            .I(N__52593));
    LocalMux I__12828 (
            .O(N__52816),
            .I(N__52586));
    LocalMux I__12827 (
            .O(N__52811),
            .I(N__52586));
    LocalMux I__12826 (
            .O(N__52808),
            .I(N__52586));
    Span4Mux_v I__12825 (
            .O(N__52803),
            .I(N__52581));
    Span4Mux_v I__12824 (
            .O(N__52800),
            .I(N__52581));
    LocalMux I__12823 (
            .O(N__52793),
            .I(N__52574));
    Span4Mux_v I__12822 (
            .O(N__52788),
            .I(N__52574));
    LocalMux I__12821 (
            .O(N__52785),
            .I(N__52574));
    Span4Mux_v I__12820 (
            .O(N__52782),
            .I(N__52567));
    LocalMux I__12819 (
            .O(N__52775),
            .I(N__52567));
    LocalMux I__12818 (
            .O(N__52766),
            .I(N__52567));
    LocalMux I__12817 (
            .O(N__52759),
            .I(N__52564));
    LocalMux I__12816 (
            .O(N__52742),
            .I(N__52561));
    InMux I__12815 (
            .O(N__52741),
            .I(N__52558));
    InMux I__12814 (
            .O(N__52738),
            .I(N__52555));
    InMux I__12813 (
            .O(N__52735),
            .I(N__52550));
    InMux I__12812 (
            .O(N__52732),
            .I(N__52550));
    Span4Mux_s3_v I__12811 (
            .O(N__52729),
            .I(N__52545));
    LocalMux I__12810 (
            .O(N__52726),
            .I(N__52545));
    InMux I__12809 (
            .O(N__52723),
            .I(N__52541));
    Span4Mux_h I__12808 (
            .O(N__52720),
            .I(N__52538));
    InMux I__12807 (
            .O(N__52719),
            .I(N__52534));
    InMux I__12806 (
            .O(N__52718),
            .I(N__52531));
    LocalMux I__12805 (
            .O(N__52713),
            .I(N__52526));
    LocalMux I__12804 (
            .O(N__52710),
            .I(N__52526));
    Span4Mux_v I__12803 (
            .O(N__52703),
            .I(N__52523));
    InMux I__12802 (
            .O(N__52700),
            .I(N__52520));
    InMux I__12801 (
            .O(N__52697),
            .I(N__52517));
    InMux I__12800 (
            .O(N__52694),
            .I(N__52512));
    InMux I__12799 (
            .O(N__52691),
            .I(N__52512));
    LocalMux I__12798 (
            .O(N__52688),
            .I(N__52509));
    LocalMux I__12797 (
            .O(N__52683),
            .I(N__52498));
    Span4Mux_s2_v I__12796 (
            .O(N__52674),
            .I(N__52498));
    LocalMux I__12795 (
            .O(N__52669),
            .I(N__52498));
    Span4Mux_h I__12794 (
            .O(N__52664),
            .I(N__52498));
    LocalMux I__12793 (
            .O(N__52657),
            .I(N__52498));
    LocalMux I__12792 (
            .O(N__52654),
            .I(N__52491));
    Span4Mux_v I__12791 (
            .O(N__52647),
            .I(N__52491));
    LocalMux I__12790 (
            .O(N__52640),
            .I(N__52491));
    Span4Mux_v I__12789 (
            .O(N__52633),
            .I(N__52486));
    LocalMux I__12788 (
            .O(N__52630),
            .I(N__52486));
    LocalMux I__12787 (
            .O(N__52625),
            .I(N__52483));
    Span4Mux_v I__12786 (
            .O(N__52620),
            .I(N__52474));
    Span4Mux_s2_v I__12785 (
            .O(N__52617),
            .I(N__52474));
    Span4Mux_s2_v I__12784 (
            .O(N__52610),
            .I(N__52474));
    Span4Mux_h I__12783 (
            .O(N__52605),
            .I(N__52474));
    LocalMux I__12782 (
            .O(N__52602),
            .I(N__52469));
    Sp12to4 I__12781 (
            .O(N__52599),
            .I(N__52469));
    CascadeMux I__12780 (
            .O(N__52598),
            .I(N__52466));
    LocalMux I__12779 (
            .O(N__52593),
            .I(N__52463));
    Span4Mux_v I__12778 (
            .O(N__52586),
            .I(N__52456));
    Span4Mux_h I__12777 (
            .O(N__52581),
            .I(N__52456));
    Span4Mux_v I__12776 (
            .O(N__52574),
            .I(N__52456));
    Span4Mux_h I__12775 (
            .O(N__52567),
            .I(N__52449));
    Span4Mux_v I__12774 (
            .O(N__52564),
            .I(N__52449));
    Span4Mux_v I__12773 (
            .O(N__52561),
            .I(N__52449));
    LocalMux I__12772 (
            .O(N__52558),
            .I(N__52444));
    LocalMux I__12771 (
            .O(N__52555),
            .I(N__52437));
    LocalMux I__12770 (
            .O(N__52550),
            .I(N__52437));
    Span4Mux_h I__12769 (
            .O(N__52545),
            .I(N__52437));
    InMux I__12768 (
            .O(N__52544),
            .I(N__52434));
    LocalMux I__12767 (
            .O(N__52541),
            .I(N__52429));
    Sp12to4 I__12766 (
            .O(N__52538),
            .I(N__52429));
    InMux I__12765 (
            .O(N__52537),
            .I(N__52426));
    LocalMux I__12764 (
            .O(N__52534),
            .I(N__52419));
    LocalMux I__12763 (
            .O(N__52531),
            .I(N__52419));
    Sp12to4 I__12762 (
            .O(N__52526),
            .I(N__52419));
    Sp12to4 I__12761 (
            .O(N__52523),
            .I(N__52416));
    LocalMux I__12760 (
            .O(N__52520),
            .I(N__52401));
    LocalMux I__12759 (
            .O(N__52517),
            .I(N__52401));
    LocalMux I__12758 (
            .O(N__52512),
            .I(N__52401));
    Span4Mux_v I__12757 (
            .O(N__52509),
            .I(N__52401));
    Span4Mux_v I__12756 (
            .O(N__52498),
            .I(N__52401));
    Span4Mux_v I__12755 (
            .O(N__52491),
            .I(N__52401));
    Span4Mux_h I__12754 (
            .O(N__52486),
            .I(N__52401));
    Span4Mux_v I__12753 (
            .O(N__52483),
            .I(N__52396));
    Span4Mux_h I__12752 (
            .O(N__52474),
            .I(N__52396));
    Span12Mux_s7_v I__12751 (
            .O(N__52469),
            .I(N__52393));
    InMux I__12750 (
            .O(N__52466),
            .I(N__52390));
    Span4Mux_h I__12749 (
            .O(N__52463),
            .I(N__52385));
    Span4Mux_h I__12748 (
            .O(N__52456),
            .I(N__52385));
    Sp12to4 I__12747 (
            .O(N__52449),
            .I(N__52382));
    InMux I__12746 (
            .O(N__52448),
            .I(N__52379));
    InMux I__12745 (
            .O(N__52447),
            .I(N__52376));
    Span4Mux_v I__12744 (
            .O(N__52444),
            .I(N__52371));
    Span4Mux_h I__12743 (
            .O(N__52437),
            .I(N__52371));
    LocalMux I__12742 (
            .O(N__52434),
            .I(N__52360));
    Span12Mux_v I__12741 (
            .O(N__52429),
            .I(N__52360));
    LocalMux I__12740 (
            .O(N__52426),
            .I(N__52360));
    Span12Mux_s6_v I__12739 (
            .O(N__52419),
            .I(N__52360));
    Span12Mux_s11_h I__12738 (
            .O(N__52416),
            .I(N__52360));
    Span4Mux_v I__12737 (
            .O(N__52401),
            .I(N__52357));
    Span4Mux_h I__12736 (
            .O(N__52396),
            .I(N__52354));
    Span12Mux_h I__12735 (
            .O(N__52393),
            .I(N__52351));
    LocalMux I__12734 (
            .O(N__52390),
            .I(N__52344));
    Sp12to4 I__12733 (
            .O(N__52385),
            .I(N__52344));
    Span12Mux_h I__12732 (
            .O(N__52382),
            .I(N__52344));
    LocalMux I__12731 (
            .O(N__52379),
            .I(opZ0Z_2));
    LocalMux I__12730 (
            .O(N__52376),
            .I(opZ0Z_2));
    Odrv4 I__12729 (
            .O(N__52371),
            .I(opZ0Z_2));
    Odrv12 I__12728 (
            .O(N__52360),
            .I(opZ0Z_2));
    Odrv4 I__12727 (
            .O(N__52357),
            .I(opZ0Z_2));
    Odrv4 I__12726 (
            .O(N__52354),
            .I(opZ0Z_2));
    Odrv12 I__12725 (
            .O(N__52351),
            .I(opZ0Z_2));
    Odrv12 I__12724 (
            .O(N__52344),
            .I(opZ0Z_2));
    InMux I__12723 (
            .O(N__52327),
            .I(N__52317));
    InMux I__12722 (
            .O(N__52326),
            .I(N__52314));
    InMux I__12721 (
            .O(N__52325),
            .I(N__52311));
    InMux I__12720 (
            .O(N__52324),
            .I(N__52303));
    InMux I__12719 (
            .O(N__52323),
            .I(N__52303));
    InMux I__12718 (
            .O(N__52322),
            .I(N__52294));
    InMux I__12717 (
            .O(N__52321),
            .I(N__52294));
    InMux I__12716 (
            .O(N__52320),
            .I(N__52290));
    LocalMux I__12715 (
            .O(N__52317),
            .I(N__52287));
    LocalMux I__12714 (
            .O(N__52314),
            .I(N__52284));
    LocalMux I__12713 (
            .O(N__52311),
            .I(N__52281));
    InMux I__12712 (
            .O(N__52310),
            .I(N__52278));
    InMux I__12711 (
            .O(N__52309),
            .I(N__52272));
    CascadeMux I__12710 (
            .O(N__52308),
            .I(N__52269));
    LocalMux I__12709 (
            .O(N__52303),
            .I(N__52266));
    InMux I__12708 (
            .O(N__52302),
            .I(N__52263));
    InMux I__12707 (
            .O(N__52301),
            .I(N__52260));
    InMux I__12706 (
            .O(N__52300),
            .I(N__52257));
    InMux I__12705 (
            .O(N__52299),
            .I(N__52250));
    LocalMux I__12704 (
            .O(N__52294),
            .I(N__52247));
    InMux I__12703 (
            .O(N__52293),
            .I(N__52244));
    LocalMux I__12702 (
            .O(N__52290),
            .I(N__52241));
    Span4Mux_v I__12701 (
            .O(N__52287),
            .I(N__52232));
    Span4Mux_v I__12700 (
            .O(N__52284),
            .I(N__52232));
    Span4Mux_h I__12699 (
            .O(N__52281),
            .I(N__52232));
    LocalMux I__12698 (
            .O(N__52278),
            .I(N__52232));
    InMux I__12697 (
            .O(N__52277),
            .I(N__52229));
    InMux I__12696 (
            .O(N__52276),
            .I(N__52223));
    InMux I__12695 (
            .O(N__52275),
            .I(N__52223));
    LocalMux I__12694 (
            .O(N__52272),
            .I(N__52218));
    InMux I__12693 (
            .O(N__52269),
            .I(N__52215));
    Span4Mux_v I__12692 (
            .O(N__52266),
            .I(N__52212));
    LocalMux I__12691 (
            .O(N__52263),
            .I(N__52205));
    LocalMux I__12690 (
            .O(N__52260),
            .I(N__52205));
    LocalMux I__12689 (
            .O(N__52257),
            .I(N__52205));
    InMux I__12688 (
            .O(N__52256),
            .I(N__52200));
    InMux I__12687 (
            .O(N__52255),
            .I(N__52200));
    CascadeMux I__12686 (
            .O(N__52254),
            .I(N__52195));
    InMux I__12685 (
            .O(N__52253),
            .I(N__52192));
    LocalMux I__12684 (
            .O(N__52250),
            .I(N__52189));
    Span4Mux_v I__12683 (
            .O(N__52247),
            .I(N__52184));
    LocalMux I__12682 (
            .O(N__52244),
            .I(N__52184));
    Span4Mux_v I__12681 (
            .O(N__52241),
            .I(N__52177));
    Span4Mux_v I__12680 (
            .O(N__52232),
            .I(N__52177));
    LocalMux I__12679 (
            .O(N__52229),
            .I(N__52177));
    CascadeMux I__12678 (
            .O(N__52228),
            .I(N__52174));
    LocalMux I__12677 (
            .O(N__52223),
            .I(N__52171));
    InMux I__12676 (
            .O(N__52222),
            .I(N__52168));
    InMux I__12675 (
            .O(N__52221),
            .I(N__52165));
    Span4Mux_v I__12674 (
            .O(N__52218),
            .I(N__52162));
    LocalMux I__12673 (
            .O(N__52215),
            .I(N__52159));
    Span4Mux_h I__12672 (
            .O(N__52212),
            .I(N__52152));
    Span4Mux_v I__12671 (
            .O(N__52205),
            .I(N__52152));
    LocalMux I__12670 (
            .O(N__52200),
            .I(N__52152));
    InMux I__12669 (
            .O(N__52199),
            .I(N__52144));
    InMux I__12668 (
            .O(N__52198),
            .I(N__52144));
    InMux I__12667 (
            .O(N__52195),
            .I(N__52144));
    LocalMux I__12666 (
            .O(N__52192),
            .I(N__52140));
    Span4Mux_s3_h I__12665 (
            .O(N__52189),
            .I(N__52136));
    Span4Mux_v I__12664 (
            .O(N__52184),
            .I(N__52131));
    Span4Mux_h I__12663 (
            .O(N__52177),
            .I(N__52131));
    InMux I__12662 (
            .O(N__52174),
            .I(N__52128));
    Span4Mux_s3_h I__12661 (
            .O(N__52171),
            .I(N__52123));
    LocalMux I__12660 (
            .O(N__52168),
            .I(N__52123));
    LocalMux I__12659 (
            .O(N__52165),
            .I(N__52118));
    Span4Mux_v I__12658 (
            .O(N__52162),
            .I(N__52111));
    Span4Mux_v I__12657 (
            .O(N__52159),
            .I(N__52111));
    Span4Mux_v I__12656 (
            .O(N__52152),
            .I(N__52111));
    InMux I__12655 (
            .O(N__52151),
            .I(N__52108));
    LocalMux I__12654 (
            .O(N__52144),
            .I(N__52105));
    InMux I__12653 (
            .O(N__52143),
            .I(N__52099));
    Span4Mux_h I__12652 (
            .O(N__52140),
            .I(N__52096));
    InMux I__12651 (
            .O(N__52139),
            .I(N__52093));
    Span4Mux_v I__12650 (
            .O(N__52136),
            .I(N__52084));
    Span4Mux_h I__12649 (
            .O(N__52131),
            .I(N__52084));
    LocalMux I__12648 (
            .O(N__52128),
            .I(N__52084));
    Span4Mux_v I__12647 (
            .O(N__52123),
            .I(N__52084));
    InMux I__12646 (
            .O(N__52122),
            .I(N__52079));
    InMux I__12645 (
            .O(N__52121),
            .I(N__52079));
    Span12Mux_v I__12644 (
            .O(N__52118),
            .I(N__52070));
    Sp12to4 I__12643 (
            .O(N__52111),
            .I(N__52070));
    LocalMux I__12642 (
            .O(N__52108),
            .I(N__52070));
    Span12Mux_s4_v I__12641 (
            .O(N__52105),
            .I(N__52070));
    InMux I__12640 (
            .O(N__52104),
            .I(N__52063));
    InMux I__12639 (
            .O(N__52103),
            .I(N__52063));
    InMux I__12638 (
            .O(N__52102),
            .I(N__52063));
    LocalMux I__12637 (
            .O(N__52099),
            .I(\ALU.a_9 ));
    Odrv4 I__12636 (
            .O(N__52096),
            .I(\ALU.a_9 ));
    LocalMux I__12635 (
            .O(N__52093),
            .I(\ALU.a_9 ));
    Odrv4 I__12634 (
            .O(N__52084),
            .I(\ALU.a_9 ));
    LocalMux I__12633 (
            .O(N__52079),
            .I(\ALU.a_9 ));
    Odrv12 I__12632 (
            .O(N__52070),
            .I(\ALU.a_9 ));
    LocalMux I__12631 (
            .O(N__52063),
            .I(\ALU.a_9 ));
    InMux I__12630 (
            .O(N__52048),
            .I(N__52045));
    LocalMux I__12629 (
            .O(N__52045),
            .I(N__52042));
    Span4Mux_v I__12628 (
            .O(N__52042),
            .I(N__52039));
    Odrv4 I__12627 (
            .O(N__52039),
            .I(\ALU.r0_12_prm_4_9_s1_c_RNOZ0 ));
    InMux I__12626 (
            .O(N__52036),
            .I(N__52030));
    CascadeMux I__12625 (
            .O(N__52035),
            .I(N__52025));
    InMux I__12624 (
            .O(N__52034),
            .I(N__52021));
    InMux I__12623 (
            .O(N__52033),
            .I(N__52018));
    LocalMux I__12622 (
            .O(N__52030),
            .I(N__52015));
    CascadeMux I__12621 (
            .O(N__52029),
            .I(N__52012));
    InMux I__12620 (
            .O(N__52028),
            .I(N__52009));
    InMux I__12619 (
            .O(N__52025),
            .I(N__52004));
    InMux I__12618 (
            .O(N__52024),
            .I(N__52004));
    LocalMux I__12617 (
            .O(N__52021),
            .I(N__51997));
    LocalMux I__12616 (
            .O(N__52018),
            .I(N__51992));
    Span4Mux_v I__12615 (
            .O(N__52015),
            .I(N__51992));
    InMux I__12614 (
            .O(N__52012),
            .I(N__51989));
    LocalMux I__12613 (
            .O(N__52009),
            .I(N__51984));
    LocalMux I__12612 (
            .O(N__52004),
            .I(N__51980));
    InMux I__12611 (
            .O(N__52003),
            .I(N__51976));
    InMux I__12610 (
            .O(N__52002),
            .I(N__51972));
    InMux I__12609 (
            .O(N__52001),
            .I(N__51969));
    InMux I__12608 (
            .O(N__52000),
            .I(N__51966));
    Span4Mux_v I__12607 (
            .O(N__51997),
            .I(N__51959));
    Span4Mux_h I__12606 (
            .O(N__51992),
            .I(N__51959));
    LocalMux I__12605 (
            .O(N__51989),
            .I(N__51959));
    InMux I__12604 (
            .O(N__51988),
            .I(N__51953));
    InMux I__12603 (
            .O(N__51987),
            .I(N__51953));
    Span4Mux_h I__12602 (
            .O(N__51984),
            .I(N__51950));
    InMux I__12601 (
            .O(N__51983),
            .I(N__51947));
    Span4Mux_h I__12600 (
            .O(N__51980),
            .I(N__51944));
    CascadeMux I__12599 (
            .O(N__51979),
            .I(N__51941));
    LocalMux I__12598 (
            .O(N__51976),
            .I(N__51936));
    InMux I__12597 (
            .O(N__51975),
            .I(N__51933));
    LocalMux I__12596 (
            .O(N__51972),
            .I(N__51928));
    LocalMux I__12595 (
            .O(N__51969),
            .I(N__51928));
    LocalMux I__12594 (
            .O(N__51966),
            .I(N__51923));
    Span4Mux_h I__12593 (
            .O(N__51959),
            .I(N__51923));
    CascadeMux I__12592 (
            .O(N__51958),
            .I(N__51920));
    LocalMux I__12591 (
            .O(N__51953),
            .I(N__51914));
    Span4Mux_h I__12590 (
            .O(N__51950),
            .I(N__51909));
    LocalMux I__12589 (
            .O(N__51947),
            .I(N__51909));
    Span4Mux_h I__12588 (
            .O(N__51944),
            .I(N__51905));
    InMux I__12587 (
            .O(N__51941),
            .I(N__51902));
    InMux I__12586 (
            .O(N__51940),
            .I(N__51899));
    InMux I__12585 (
            .O(N__51939),
            .I(N__51896));
    Span4Mux_h I__12584 (
            .O(N__51936),
            .I(N__51891));
    LocalMux I__12583 (
            .O(N__51933),
            .I(N__51891));
    Span12Mux_h I__12582 (
            .O(N__51928),
            .I(N__51888));
    Span4Mux_h I__12581 (
            .O(N__51923),
            .I(N__51885));
    InMux I__12580 (
            .O(N__51920),
            .I(N__51878));
    InMux I__12579 (
            .O(N__51919),
            .I(N__51878));
    InMux I__12578 (
            .O(N__51918),
            .I(N__51878));
    InMux I__12577 (
            .O(N__51917),
            .I(N__51875));
    Span4Mux_v I__12576 (
            .O(N__51914),
            .I(N__51870));
    Span4Mux_v I__12575 (
            .O(N__51909),
            .I(N__51870));
    InMux I__12574 (
            .O(N__51908),
            .I(N__51867));
    Span4Mux_v I__12573 (
            .O(N__51905),
            .I(N__51856));
    LocalMux I__12572 (
            .O(N__51902),
            .I(N__51856));
    LocalMux I__12571 (
            .O(N__51899),
            .I(N__51856));
    LocalMux I__12570 (
            .O(N__51896),
            .I(N__51856));
    Span4Mux_h I__12569 (
            .O(N__51891),
            .I(N__51856));
    Odrv12 I__12568 (
            .O(N__51888),
            .I(\ALU.b_10 ));
    Odrv4 I__12567 (
            .O(N__51885),
            .I(\ALU.b_10 ));
    LocalMux I__12566 (
            .O(N__51878),
            .I(\ALU.b_10 ));
    LocalMux I__12565 (
            .O(N__51875),
            .I(\ALU.b_10 ));
    Odrv4 I__12564 (
            .O(N__51870),
            .I(\ALU.b_10 ));
    LocalMux I__12563 (
            .O(N__51867),
            .I(\ALU.b_10 ));
    Odrv4 I__12562 (
            .O(N__51856),
            .I(\ALU.b_10 ));
    InMux I__12561 (
            .O(N__51841),
            .I(N__51833));
    InMux I__12560 (
            .O(N__51840),
            .I(N__51822));
    CascadeMux I__12559 (
            .O(N__51839),
            .I(N__51819));
    CascadeMux I__12558 (
            .O(N__51838),
            .I(N__51816));
    InMux I__12557 (
            .O(N__51837),
            .I(N__51812));
    InMux I__12556 (
            .O(N__51836),
            .I(N__51801));
    LocalMux I__12555 (
            .O(N__51833),
            .I(N__51798));
    InMux I__12554 (
            .O(N__51832),
            .I(N__51791));
    InMux I__12553 (
            .O(N__51831),
            .I(N__51788));
    InMux I__12552 (
            .O(N__51830),
            .I(N__51781));
    InMux I__12551 (
            .O(N__51829),
            .I(N__51781));
    InMux I__12550 (
            .O(N__51828),
            .I(N__51781));
    InMux I__12549 (
            .O(N__51827),
            .I(N__51776));
    InMux I__12548 (
            .O(N__51826),
            .I(N__51776));
    InMux I__12547 (
            .O(N__51825),
            .I(N__51773));
    LocalMux I__12546 (
            .O(N__51822),
            .I(N__51770));
    InMux I__12545 (
            .O(N__51819),
            .I(N__51767));
    InMux I__12544 (
            .O(N__51816),
            .I(N__51762));
    InMux I__12543 (
            .O(N__51815),
            .I(N__51762));
    LocalMux I__12542 (
            .O(N__51812),
            .I(N__51759));
    InMux I__12541 (
            .O(N__51811),
            .I(N__51756));
    InMux I__12540 (
            .O(N__51810),
            .I(N__51751));
    InMux I__12539 (
            .O(N__51809),
            .I(N__51751));
    InMux I__12538 (
            .O(N__51808),
            .I(N__51748));
    CascadeMux I__12537 (
            .O(N__51807),
            .I(N__51744));
    CascadeMux I__12536 (
            .O(N__51806),
            .I(N__51739));
    InMux I__12535 (
            .O(N__51805),
            .I(N__51736));
    InMux I__12534 (
            .O(N__51804),
            .I(N__51733));
    LocalMux I__12533 (
            .O(N__51801),
            .I(N__51729));
    Span4Mux_v I__12532 (
            .O(N__51798),
            .I(N__51726));
    InMux I__12531 (
            .O(N__51797),
            .I(N__51723));
    InMux I__12530 (
            .O(N__51796),
            .I(N__51720));
    InMux I__12529 (
            .O(N__51795),
            .I(N__51717));
    InMux I__12528 (
            .O(N__51794),
            .I(N__51713));
    LocalMux I__12527 (
            .O(N__51791),
            .I(N__51702));
    LocalMux I__12526 (
            .O(N__51788),
            .I(N__51702));
    LocalMux I__12525 (
            .O(N__51781),
            .I(N__51702));
    LocalMux I__12524 (
            .O(N__51776),
            .I(N__51702));
    LocalMux I__12523 (
            .O(N__51773),
            .I(N__51702));
    Span4Mux_v I__12522 (
            .O(N__51770),
            .I(N__51699));
    LocalMux I__12521 (
            .O(N__51767),
            .I(N__51696));
    LocalMux I__12520 (
            .O(N__51762),
            .I(N__51691));
    Span4Mux_v I__12519 (
            .O(N__51759),
            .I(N__51691));
    LocalMux I__12518 (
            .O(N__51756),
            .I(N__51688));
    LocalMux I__12517 (
            .O(N__51751),
            .I(N__51683));
    LocalMux I__12516 (
            .O(N__51748),
            .I(N__51683));
    InMux I__12515 (
            .O(N__51747),
            .I(N__51680));
    InMux I__12514 (
            .O(N__51744),
            .I(N__51677));
    InMux I__12513 (
            .O(N__51743),
            .I(N__51672));
    InMux I__12512 (
            .O(N__51742),
            .I(N__51672));
    InMux I__12511 (
            .O(N__51739),
            .I(N__51669));
    LocalMux I__12510 (
            .O(N__51736),
            .I(N__51666));
    LocalMux I__12509 (
            .O(N__51733),
            .I(N__51663));
    InMux I__12508 (
            .O(N__51732),
            .I(N__51660));
    Span12Mux_s4_h I__12507 (
            .O(N__51729),
            .I(N__51653));
    Sp12to4 I__12506 (
            .O(N__51726),
            .I(N__51653));
    LocalMux I__12505 (
            .O(N__51723),
            .I(N__51653));
    LocalMux I__12504 (
            .O(N__51720),
            .I(N__51649));
    LocalMux I__12503 (
            .O(N__51717),
            .I(N__51646));
    InMux I__12502 (
            .O(N__51716),
            .I(N__51643));
    LocalMux I__12501 (
            .O(N__51713),
            .I(N__51638));
    Span4Mux_v I__12500 (
            .O(N__51702),
            .I(N__51638));
    Span4Mux_h I__12499 (
            .O(N__51699),
            .I(N__51631));
    Span4Mux_v I__12498 (
            .O(N__51696),
            .I(N__51631));
    Span4Mux_h I__12497 (
            .O(N__51691),
            .I(N__51631));
    Span4Mux_v I__12496 (
            .O(N__51688),
            .I(N__51626));
    Span4Mux_v I__12495 (
            .O(N__51683),
            .I(N__51626));
    LocalMux I__12494 (
            .O(N__51680),
            .I(N__51623));
    LocalMux I__12493 (
            .O(N__51677),
            .I(N__51620));
    LocalMux I__12492 (
            .O(N__51672),
            .I(N__51617));
    LocalMux I__12491 (
            .O(N__51669),
            .I(N__51614));
    Span4Mux_v I__12490 (
            .O(N__51666),
            .I(N__51607));
    Span4Mux_h I__12489 (
            .O(N__51663),
            .I(N__51607));
    LocalMux I__12488 (
            .O(N__51660),
            .I(N__51607));
    Span12Mux_h I__12487 (
            .O(N__51653),
            .I(N__51604));
    InMux I__12486 (
            .O(N__51652),
            .I(N__51601));
    Sp12to4 I__12485 (
            .O(N__51649),
            .I(N__51594));
    Span12Mux_s9_v I__12484 (
            .O(N__51646),
            .I(N__51594));
    LocalMux I__12483 (
            .O(N__51643),
            .I(N__51594));
    Span4Mux_h I__12482 (
            .O(N__51638),
            .I(N__51587));
    Span4Mux_h I__12481 (
            .O(N__51631),
            .I(N__51587));
    Span4Mux_h I__12480 (
            .O(N__51626),
            .I(N__51587));
    Span4Mux_h I__12479 (
            .O(N__51623),
            .I(N__51582));
    Span4Mux_v I__12478 (
            .O(N__51620),
            .I(N__51582));
    Span4Mux_h I__12477 (
            .O(N__51617),
            .I(N__51575));
    Span4Mux_v I__12476 (
            .O(N__51614),
            .I(N__51575));
    Span4Mux_h I__12475 (
            .O(N__51607),
            .I(N__51575));
    Odrv12 I__12474 (
            .O(N__51604),
            .I(\ALU.a_10 ));
    LocalMux I__12473 (
            .O(N__51601),
            .I(\ALU.a_10 ));
    Odrv12 I__12472 (
            .O(N__51594),
            .I(\ALU.a_10 ));
    Odrv4 I__12471 (
            .O(N__51587),
            .I(\ALU.a_10 ));
    Odrv4 I__12470 (
            .O(N__51582),
            .I(\ALU.a_10 ));
    Odrv4 I__12469 (
            .O(N__51575),
            .I(\ALU.a_10 ));
    CascadeMux I__12468 (
            .O(N__51562),
            .I(N__51559));
    InMux I__12467 (
            .O(N__51559),
            .I(N__51556));
    LocalMux I__12466 (
            .O(N__51556),
            .I(N__51553));
    Span4Mux_h I__12465 (
            .O(N__51553),
            .I(N__51550));
    Span4Mux_h I__12464 (
            .O(N__51550),
            .I(N__51547));
    Span4Mux_h I__12463 (
            .O(N__51547),
            .I(N__51544));
    Odrv4 I__12462 (
            .O(N__51544),
            .I(\ALU.r0_12_prm_7_10_s0_c_RNOZ0 ));
    CascadeMux I__12461 (
            .O(N__51541),
            .I(N__51538));
    InMux I__12460 (
            .O(N__51538),
            .I(N__51534));
    CascadeMux I__12459 (
            .O(N__51537),
            .I(N__51524));
    LocalMux I__12458 (
            .O(N__51534),
            .I(N__51515));
    CascadeMux I__12457 (
            .O(N__51533),
            .I(N__51510));
    CascadeMux I__12456 (
            .O(N__51532),
            .I(N__51504));
    CascadeMux I__12455 (
            .O(N__51531),
            .I(N__51501));
    CascadeMux I__12454 (
            .O(N__51530),
            .I(N__51495));
    CascadeMux I__12453 (
            .O(N__51529),
            .I(N__51492));
    CascadeMux I__12452 (
            .O(N__51528),
            .I(N__51488));
    CascadeMux I__12451 (
            .O(N__51527),
            .I(N__51485));
    InMux I__12450 (
            .O(N__51524),
            .I(N__51479));
    InMux I__12449 (
            .O(N__51523),
            .I(N__51476));
    CascadeMux I__12448 (
            .O(N__51522),
            .I(N__51469));
    CascadeMux I__12447 (
            .O(N__51521),
            .I(N__51466));
    CascadeMux I__12446 (
            .O(N__51520),
            .I(N__51462));
    InMux I__12445 (
            .O(N__51519),
            .I(N__51457));
    InMux I__12444 (
            .O(N__51518),
            .I(N__51457));
    Span4Mux_v I__12443 (
            .O(N__51515),
            .I(N__51454));
    InMux I__12442 (
            .O(N__51514),
            .I(N__51447));
    InMux I__12441 (
            .O(N__51513),
            .I(N__51447));
    InMux I__12440 (
            .O(N__51510),
            .I(N__51447));
    InMux I__12439 (
            .O(N__51509),
            .I(N__51443));
    InMux I__12438 (
            .O(N__51508),
            .I(N__51438));
    InMux I__12437 (
            .O(N__51507),
            .I(N__51435));
    InMux I__12436 (
            .O(N__51504),
            .I(N__51430));
    InMux I__12435 (
            .O(N__51501),
            .I(N__51430));
    CascadeMux I__12434 (
            .O(N__51500),
            .I(N__51427));
    CascadeMux I__12433 (
            .O(N__51499),
            .I(N__51424));
    InMux I__12432 (
            .O(N__51498),
            .I(N__51420));
    InMux I__12431 (
            .O(N__51495),
            .I(N__51415));
    InMux I__12430 (
            .O(N__51492),
            .I(N__51415));
    CascadeMux I__12429 (
            .O(N__51491),
            .I(N__51411));
    InMux I__12428 (
            .O(N__51488),
            .I(N__51406));
    InMux I__12427 (
            .O(N__51485),
            .I(N__51406));
    CascadeMux I__12426 (
            .O(N__51484),
            .I(N__51403));
    CascadeMux I__12425 (
            .O(N__51483),
            .I(N__51400));
    CascadeMux I__12424 (
            .O(N__51482),
            .I(N__51397));
    LocalMux I__12423 (
            .O(N__51479),
            .I(N__51392));
    LocalMux I__12422 (
            .O(N__51476),
            .I(N__51392));
    InMux I__12421 (
            .O(N__51475),
            .I(N__51389));
    InMux I__12420 (
            .O(N__51474),
            .I(N__51386));
    InMux I__12419 (
            .O(N__51473),
            .I(N__51381));
    InMux I__12418 (
            .O(N__51472),
            .I(N__51381));
    InMux I__12417 (
            .O(N__51469),
            .I(N__51378));
    InMux I__12416 (
            .O(N__51466),
            .I(N__51371));
    InMux I__12415 (
            .O(N__51465),
            .I(N__51371));
    InMux I__12414 (
            .O(N__51462),
            .I(N__51371));
    LocalMux I__12413 (
            .O(N__51457),
            .I(N__51368));
    Span4Mux_h I__12412 (
            .O(N__51454),
            .I(N__51363));
    LocalMux I__12411 (
            .O(N__51447),
            .I(N__51363));
    CascadeMux I__12410 (
            .O(N__51446),
            .I(N__51360));
    LocalMux I__12409 (
            .O(N__51443),
            .I(N__51356));
    InMux I__12408 (
            .O(N__51442),
            .I(N__51353));
    InMux I__12407 (
            .O(N__51441),
            .I(N__51350));
    LocalMux I__12406 (
            .O(N__51438),
            .I(N__51347));
    LocalMux I__12405 (
            .O(N__51435),
            .I(N__51342));
    LocalMux I__12404 (
            .O(N__51430),
            .I(N__51342));
    InMux I__12403 (
            .O(N__51427),
            .I(N__51337));
    InMux I__12402 (
            .O(N__51424),
            .I(N__51337));
    InMux I__12401 (
            .O(N__51423),
            .I(N__51334));
    LocalMux I__12400 (
            .O(N__51420),
            .I(N__51329));
    LocalMux I__12399 (
            .O(N__51415),
            .I(N__51329));
    InMux I__12398 (
            .O(N__51414),
            .I(N__51326));
    InMux I__12397 (
            .O(N__51411),
            .I(N__51323));
    LocalMux I__12396 (
            .O(N__51406),
            .I(N__51320));
    InMux I__12395 (
            .O(N__51403),
            .I(N__51315));
    InMux I__12394 (
            .O(N__51400),
            .I(N__51315));
    InMux I__12393 (
            .O(N__51397),
            .I(N__51312));
    Span4Mux_v I__12392 (
            .O(N__51392),
            .I(N__51305));
    LocalMux I__12391 (
            .O(N__51389),
            .I(N__51305));
    LocalMux I__12390 (
            .O(N__51386),
            .I(N__51305));
    LocalMux I__12389 (
            .O(N__51381),
            .I(N__51297));
    LocalMux I__12388 (
            .O(N__51378),
            .I(N__51291));
    LocalMux I__12387 (
            .O(N__51371),
            .I(N__51291));
    Span4Mux_v I__12386 (
            .O(N__51368),
            .I(N__51286));
    Span4Mux_v I__12385 (
            .O(N__51363),
            .I(N__51286));
    InMux I__12384 (
            .O(N__51360),
            .I(N__51281));
    InMux I__12383 (
            .O(N__51359),
            .I(N__51281));
    Span4Mux_s3_v I__12382 (
            .O(N__51356),
            .I(N__51276));
    LocalMux I__12381 (
            .O(N__51353),
            .I(N__51276));
    LocalMux I__12380 (
            .O(N__51350),
            .I(N__51269));
    Span4Mux_h I__12379 (
            .O(N__51347),
            .I(N__51269));
    Span4Mux_h I__12378 (
            .O(N__51342),
            .I(N__51269));
    LocalMux I__12377 (
            .O(N__51337),
            .I(N__51265));
    LocalMux I__12376 (
            .O(N__51334),
            .I(N__51258));
    Span4Mux_h I__12375 (
            .O(N__51329),
            .I(N__51258));
    LocalMux I__12374 (
            .O(N__51326),
            .I(N__51258));
    LocalMux I__12373 (
            .O(N__51323),
            .I(N__51247));
    Span4Mux_h I__12372 (
            .O(N__51320),
            .I(N__51247));
    LocalMux I__12371 (
            .O(N__51315),
            .I(N__51247));
    LocalMux I__12370 (
            .O(N__51312),
            .I(N__51247));
    Span4Mux_v I__12369 (
            .O(N__51305),
            .I(N__51247));
    CascadeMux I__12368 (
            .O(N__51304),
            .I(N__51241));
    InMux I__12367 (
            .O(N__51303),
            .I(N__51238));
    CascadeMux I__12366 (
            .O(N__51302),
            .I(N__51235));
    CascadeMux I__12365 (
            .O(N__51301),
            .I(N__51232));
    InMux I__12364 (
            .O(N__51300),
            .I(N__51228));
    Span4Mux_h I__12363 (
            .O(N__51297),
            .I(N__51225));
    CascadeMux I__12362 (
            .O(N__51296),
            .I(N__51218));
    Span4Mux_v I__12361 (
            .O(N__51291),
            .I(N__51213));
    Span4Mux_v I__12360 (
            .O(N__51286),
            .I(N__51213));
    LocalMux I__12359 (
            .O(N__51281),
            .I(N__51205));
    Span4Mux_h I__12358 (
            .O(N__51276),
            .I(N__51205));
    Span4Mux_v I__12357 (
            .O(N__51269),
            .I(N__51205));
    InMux I__12356 (
            .O(N__51268),
            .I(N__51202));
    Span4Mux_v I__12355 (
            .O(N__51265),
            .I(N__51199));
    Span4Mux_v I__12354 (
            .O(N__51258),
            .I(N__51196));
    Span4Mux_v I__12353 (
            .O(N__51247),
            .I(N__51193));
    InMux I__12352 (
            .O(N__51246),
            .I(N__51190));
    InMux I__12351 (
            .O(N__51245),
            .I(N__51185));
    InMux I__12350 (
            .O(N__51244),
            .I(N__51185));
    InMux I__12349 (
            .O(N__51241),
            .I(N__51182));
    LocalMux I__12348 (
            .O(N__51238),
            .I(N__51179));
    InMux I__12347 (
            .O(N__51235),
            .I(N__51172));
    InMux I__12346 (
            .O(N__51232),
            .I(N__51172));
    InMux I__12345 (
            .O(N__51231),
            .I(N__51172));
    LocalMux I__12344 (
            .O(N__51228),
            .I(N__51167));
    Span4Mux_h I__12343 (
            .O(N__51225),
            .I(N__51167));
    InMux I__12342 (
            .O(N__51224),
            .I(N__51164));
    InMux I__12341 (
            .O(N__51223),
            .I(N__51159));
    InMux I__12340 (
            .O(N__51222),
            .I(N__51159));
    InMux I__12339 (
            .O(N__51221),
            .I(N__51154));
    InMux I__12338 (
            .O(N__51218),
            .I(N__51154));
    Span4Mux_v I__12337 (
            .O(N__51213),
            .I(N__51151));
    InMux I__12336 (
            .O(N__51212),
            .I(N__51148));
    Span4Mux_v I__12335 (
            .O(N__51205),
            .I(N__51143));
    LocalMux I__12334 (
            .O(N__51202),
            .I(N__51143));
    Span4Mux_s0_v I__12333 (
            .O(N__51199),
            .I(N__51136));
    Span4Mux_s0_v I__12332 (
            .O(N__51196),
            .I(N__51136));
    Span4Mux_s0_v I__12331 (
            .O(N__51193),
            .I(N__51136));
    LocalMux I__12330 (
            .O(N__51190),
            .I(N__51123));
    LocalMux I__12329 (
            .O(N__51185),
            .I(N__51123));
    LocalMux I__12328 (
            .O(N__51182),
            .I(N__51123));
    Span12Mux_v I__12327 (
            .O(N__51179),
            .I(N__51123));
    LocalMux I__12326 (
            .O(N__51172),
            .I(N__51123));
    Sp12to4 I__12325 (
            .O(N__51167),
            .I(N__51123));
    LocalMux I__12324 (
            .O(N__51164),
            .I(paramsZ0Z_3));
    LocalMux I__12323 (
            .O(N__51159),
            .I(paramsZ0Z_3));
    LocalMux I__12322 (
            .O(N__51154),
            .I(paramsZ0Z_3));
    Odrv4 I__12321 (
            .O(N__51151),
            .I(paramsZ0Z_3));
    LocalMux I__12320 (
            .O(N__51148),
            .I(paramsZ0Z_3));
    Odrv4 I__12319 (
            .O(N__51143),
            .I(paramsZ0Z_3));
    Odrv4 I__12318 (
            .O(N__51136),
            .I(paramsZ0Z_3));
    Odrv12 I__12317 (
            .O(N__51123),
            .I(paramsZ0Z_3));
    InMux I__12316 (
            .O(N__51106),
            .I(N__51093));
    InMux I__12315 (
            .O(N__51105),
            .I(N__51093));
    InMux I__12314 (
            .O(N__51104),
            .I(N__51090));
    InMux I__12313 (
            .O(N__51103),
            .I(N__51084));
    InMux I__12312 (
            .O(N__51102),
            .I(N__51081));
    InMux I__12311 (
            .O(N__51101),
            .I(N__51075));
    InMux I__12310 (
            .O(N__51100),
            .I(N__51075));
    InMux I__12309 (
            .O(N__51099),
            .I(N__51071));
    InMux I__12308 (
            .O(N__51098),
            .I(N__51068));
    LocalMux I__12307 (
            .O(N__51093),
            .I(N__51065));
    LocalMux I__12306 (
            .O(N__51090),
            .I(N__51062));
    InMux I__12305 (
            .O(N__51089),
            .I(N__51059));
    CascadeMux I__12304 (
            .O(N__51088),
            .I(N__51055));
    CascadeMux I__12303 (
            .O(N__51087),
            .I(N__51051));
    LocalMux I__12302 (
            .O(N__51084),
            .I(N__51048));
    LocalMux I__12301 (
            .O(N__51081),
            .I(N__51044));
    InMux I__12300 (
            .O(N__51080),
            .I(N__51041));
    LocalMux I__12299 (
            .O(N__51075),
            .I(N__51034));
    CascadeMux I__12298 (
            .O(N__51074),
            .I(N__51029));
    LocalMux I__12297 (
            .O(N__51071),
            .I(N__51021));
    LocalMux I__12296 (
            .O(N__51068),
            .I(N__51016));
    Span4Mux_h I__12295 (
            .O(N__51065),
            .I(N__51016));
    Span4Mux_v I__12294 (
            .O(N__51062),
            .I(N__51011));
    LocalMux I__12293 (
            .O(N__51059),
            .I(N__51011));
    InMux I__12292 (
            .O(N__51058),
            .I(N__51004));
    InMux I__12291 (
            .O(N__51055),
            .I(N__51004));
    InMux I__12290 (
            .O(N__51054),
            .I(N__51004));
    InMux I__12289 (
            .O(N__51051),
            .I(N__50996));
    Span4Mux_v I__12288 (
            .O(N__51048),
            .I(N__50989));
    InMux I__12287 (
            .O(N__51047),
            .I(N__50986));
    Span4Mux_v I__12286 (
            .O(N__51044),
            .I(N__50979));
    LocalMux I__12285 (
            .O(N__51041),
            .I(N__50979));
    InMux I__12284 (
            .O(N__51040),
            .I(N__50974));
    InMux I__12283 (
            .O(N__51039),
            .I(N__50974));
    InMux I__12282 (
            .O(N__51038),
            .I(N__50971));
    InMux I__12281 (
            .O(N__51037),
            .I(N__50968));
    Span4Mux_h I__12280 (
            .O(N__51034),
            .I(N__50965));
    InMux I__12279 (
            .O(N__51033),
            .I(N__50962));
    InMux I__12278 (
            .O(N__51032),
            .I(N__50958));
    InMux I__12277 (
            .O(N__51029),
            .I(N__50955));
    InMux I__12276 (
            .O(N__51028),
            .I(N__50952));
    InMux I__12275 (
            .O(N__51027),
            .I(N__50949));
    InMux I__12274 (
            .O(N__51026),
            .I(N__50942));
    InMux I__12273 (
            .O(N__51025),
            .I(N__50942));
    InMux I__12272 (
            .O(N__51024),
            .I(N__50942));
    Span4Mux_v I__12271 (
            .O(N__51021),
            .I(N__50933));
    Span4Mux_h I__12270 (
            .O(N__51016),
            .I(N__50933));
    Span4Mux_h I__12269 (
            .O(N__51011),
            .I(N__50933));
    LocalMux I__12268 (
            .O(N__51004),
            .I(N__50933));
    InMux I__12267 (
            .O(N__51003),
            .I(N__50926));
    InMux I__12266 (
            .O(N__51002),
            .I(N__50926));
    InMux I__12265 (
            .O(N__51001),
            .I(N__50921));
    InMux I__12264 (
            .O(N__51000),
            .I(N__50921));
    InMux I__12263 (
            .O(N__50999),
            .I(N__50918));
    LocalMux I__12262 (
            .O(N__50996),
            .I(N__50915));
    InMux I__12261 (
            .O(N__50995),
            .I(N__50912));
    InMux I__12260 (
            .O(N__50994),
            .I(N__50909));
    InMux I__12259 (
            .O(N__50993),
            .I(N__50904));
    InMux I__12258 (
            .O(N__50992),
            .I(N__50904));
    Span4Mux_h I__12257 (
            .O(N__50989),
            .I(N__50899));
    LocalMux I__12256 (
            .O(N__50986),
            .I(N__50899));
    InMux I__12255 (
            .O(N__50985),
            .I(N__50894));
    InMux I__12254 (
            .O(N__50984),
            .I(N__50894));
    Span4Mux_v I__12253 (
            .O(N__50979),
            .I(N__50889));
    LocalMux I__12252 (
            .O(N__50974),
            .I(N__50889));
    LocalMux I__12251 (
            .O(N__50971),
            .I(N__50882));
    LocalMux I__12250 (
            .O(N__50968),
            .I(N__50882));
    Span4Mux_h I__12249 (
            .O(N__50965),
            .I(N__50882));
    LocalMux I__12248 (
            .O(N__50962),
            .I(N__50879));
    CascadeMux I__12247 (
            .O(N__50961),
            .I(N__50875));
    LocalMux I__12246 (
            .O(N__50958),
            .I(N__50860));
    LocalMux I__12245 (
            .O(N__50955),
            .I(N__50860));
    LocalMux I__12244 (
            .O(N__50952),
            .I(N__50860));
    LocalMux I__12243 (
            .O(N__50949),
            .I(N__50860));
    LocalMux I__12242 (
            .O(N__50942),
            .I(N__50860));
    Span4Mux_v I__12241 (
            .O(N__50933),
            .I(N__50860));
    CascadeMux I__12240 (
            .O(N__50932),
            .I(N__50857));
    CascadeMux I__12239 (
            .O(N__50931),
            .I(N__50853));
    LocalMux I__12238 (
            .O(N__50926),
            .I(N__50850));
    LocalMux I__12237 (
            .O(N__50921),
            .I(N__50845));
    LocalMux I__12236 (
            .O(N__50918),
            .I(N__50845));
    Span4Mux_h I__12235 (
            .O(N__50915),
            .I(N__50834));
    LocalMux I__12234 (
            .O(N__50912),
            .I(N__50834));
    LocalMux I__12233 (
            .O(N__50909),
            .I(N__50834));
    LocalMux I__12232 (
            .O(N__50904),
            .I(N__50834));
    Span4Mux_v I__12231 (
            .O(N__50899),
            .I(N__50834));
    LocalMux I__12230 (
            .O(N__50894),
            .I(N__50825));
    Sp12to4 I__12229 (
            .O(N__50889),
            .I(N__50825));
    Sp12to4 I__12228 (
            .O(N__50882),
            .I(N__50825));
    Span12Mux_h I__12227 (
            .O(N__50879),
            .I(N__50825));
    InMux I__12226 (
            .O(N__50878),
            .I(N__50822));
    InMux I__12225 (
            .O(N__50875),
            .I(N__50819));
    InMux I__12224 (
            .O(N__50874),
            .I(N__50816));
    InMux I__12223 (
            .O(N__50873),
            .I(N__50813));
    Span4Mux_v I__12222 (
            .O(N__50860),
            .I(N__50810));
    InMux I__12221 (
            .O(N__50857),
            .I(N__50803));
    InMux I__12220 (
            .O(N__50856),
            .I(N__50803));
    InMux I__12219 (
            .O(N__50853),
            .I(N__50803));
    Span4Mux_h I__12218 (
            .O(N__50850),
            .I(N__50800));
    Span4Mux_v I__12217 (
            .O(N__50845),
            .I(N__50795));
    Span4Mux_v I__12216 (
            .O(N__50834),
            .I(N__50795));
    Span12Mux_v I__12215 (
            .O(N__50825),
            .I(N__50792));
    LocalMux I__12214 (
            .O(N__50822),
            .I(paramsZ0Z_2));
    LocalMux I__12213 (
            .O(N__50819),
            .I(paramsZ0Z_2));
    LocalMux I__12212 (
            .O(N__50816),
            .I(paramsZ0Z_2));
    LocalMux I__12211 (
            .O(N__50813),
            .I(paramsZ0Z_2));
    Odrv4 I__12210 (
            .O(N__50810),
            .I(paramsZ0Z_2));
    LocalMux I__12209 (
            .O(N__50803),
            .I(paramsZ0Z_2));
    Odrv4 I__12208 (
            .O(N__50800),
            .I(paramsZ0Z_2));
    Odrv4 I__12207 (
            .O(N__50795),
            .I(paramsZ0Z_2));
    Odrv12 I__12206 (
            .O(N__50792),
            .I(paramsZ0Z_2));
    InMux I__12205 (
            .O(N__50773),
            .I(N__50769));
    InMux I__12204 (
            .O(N__50772),
            .I(N__50766));
    LocalMux I__12203 (
            .O(N__50769),
            .I(N__50762));
    LocalMux I__12202 (
            .O(N__50766),
            .I(N__50759));
    InMux I__12201 (
            .O(N__50765),
            .I(N__50756));
    Span4Mux_v I__12200 (
            .O(N__50762),
            .I(N__50753));
    Span4Mux_h I__12199 (
            .O(N__50759),
            .I(N__50749));
    LocalMux I__12198 (
            .O(N__50756),
            .I(N__50744));
    Span4Mux_v I__12197 (
            .O(N__50753),
            .I(N__50744));
    InMux I__12196 (
            .O(N__50752),
            .I(N__50741));
    Span4Mux_h I__12195 (
            .O(N__50749),
            .I(N__50737));
    Span4Mux_h I__12194 (
            .O(N__50744),
            .I(N__50734));
    LocalMux I__12193 (
            .O(N__50741),
            .I(N__50731));
    InMux I__12192 (
            .O(N__50740),
            .I(N__50728));
    Odrv4 I__12191 (
            .O(N__50737),
            .I(\ALU.r4_RNII2A0LZ0Z_1 ));
    Odrv4 I__12190 (
            .O(N__50734),
            .I(\ALU.r4_RNII2A0LZ0Z_1 ));
    Odrv4 I__12189 (
            .O(N__50731),
            .I(\ALU.r4_RNII2A0LZ0Z_1 ));
    LocalMux I__12188 (
            .O(N__50728),
            .I(\ALU.r4_RNII2A0LZ0Z_1 ));
    CascadeMux I__12187 (
            .O(N__50719),
            .I(N__50716));
    InMux I__12186 (
            .O(N__50716),
            .I(N__50713));
    LocalMux I__12185 (
            .O(N__50713),
            .I(N__50710));
    Odrv12 I__12184 (
            .O(N__50710),
            .I(\ALU.lshift_3 ));
    CascadeMux I__12183 (
            .O(N__50707),
            .I(N__50702));
    InMux I__12182 (
            .O(N__50706),
            .I(N__50697));
    InMux I__12181 (
            .O(N__50705),
            .I(N__50694));
    InMux I__12180 (
            .O(N__50702),
            .I(N__50691));
    InMux I__12179 (
            .O(N__50701),
            .I(N__50686));
    InMux I__12178 (
            .O(N__50700),
            .I(N__50686));
    LocalMux I__12177 (
            .O(N__50697),
            .I(N__50683));
    LocalMux I__12176 (
            .O(N__50694),
            .I(N__50680));
    LocalMux I__12175 (
            .O(N__50691),
            .I(N__50676));
    LocalMux I__12174 (
            .O(N__50686),
            .I(N__50673));
    Span4Mux_v I__12173 (
            .O(N__50683),
            .I(N__50670));
    Span4Mux_h I__12172 (
            .O(N__50680),
            .I(N__50666));
    CascadeMux I__12171 (
            .O(N__50679),
            .I(N__50663));
    Span12Mux_h I__12170 (
            .O(N__50676),
            .I(N__50660));
    Span4Mux_v I__12169 (
            .O(N__50673),
            .I(N__50657));
    Span4Mux_v I__12168 (
            .O(N__50670),
            .I(N__50654));
    CascadeMux I__12167 (
            .O(N__50669),
            .I(N__50651));
    Span4Mux_v I__12166 (
            .O(N__50666),
            .I(N__50648));
    InMux I__12165 (
            .O(N__50663),
            .I(N__50645));
    Span12Mux_v I__12164 (
            .O(N__50660),
            .I(N__50642));
    Span4Mux_v I__12163 (
            .O(N__50657),
            .I(N__50637));
    Span4Mux_v I__12162 (
            .O(N__50654),
            .I(N__50637));
    InMux I__12161 (
            .O(N__50651),
            .I(N__50634));
    Odrv4 I__12160 (
            .O(N__50648),
            .I(\ALU.lshift63Z0Z_2 ));
    LocalMux I__12159 (
            .O(N__50645),
            .I(\ALU.lshift63Z0Z_2 ));
    Odrv12 I__12158 (
            .O(N__50642),
            .I(\ALU.lshift63Z0Z_2 ));
    Odrv4 I__12157 (
            .O(N__50637),
            .I(\ALU.lshift63Z0Z_2 ));
    LocalMux I__12156 (
            .O(N__50634),
            .I(\ALU.lshift63Z0Z_2 ));
    InMux I__12155 (
            .O(N__50623),
            .I(N__50618));
    InMux I__12154 (
            .O(N__50622),
            .I(N__50615));
    InMux I__12153 (
            .O(N__50621),
            .I(N__50612));
    LocalMux I__12152 (
            .O(N__50618),
            .I(N__50607));
    LocalMux I__12151 (
            .O(N__50615),
            .I(N__50604));
    LocalMux I__12150 (
            .O(N__50612),
            .I(N__50601));
    InMux I__12149 (
            .O(N__50611),
            .I(N__50596));
    InMux I__12148 (
            .O(N__50610),
            .I(N__50596));
    Span4Mux_v I__12147 (
            .O(N__50607),
            .I(N__50593));
    Span4Mux_v I__12146 (
            .O(N__50604),
            .I(N__50590));
    Span4Mux_v I__12145 (
            .O(N__50601),
            .I(N__50587));
    LocalMux I__12144 (
            .O(N__50596),
            .I(N__50584));
    Span4Mux_h I__12143 (
            .O(N__50593),
            .I(N__50581));
    Span4Mux_h I__12142 (
            .O(N__50590),
            .I(N__50578));
    Sp12to4 I__12141 (
            .O(N__50587),
            .I(N__50573));
    Sp12to4 I__12140 (
            .O(N__50584),
            .I(N__50573));
    Sp12to4 I__12139 (
            .O(N__50581),
            .I(N__50568));
    Sp12to4 I__12138 (
            .O(N__50578),
            .I(N__50568));
    Span12Mux_h I__12137 (
            .O(N__50573),
            .I(N__50565));
    Odrv12 I__12136 (
            .O(N__50568),
            .I(\ALU.r5_RNIAG9A9Z0Z_15 ));
    Odrv12 I__12135 (
            .O(N__50565),
            .I(\ALU.r5_RNIAG9A9Z0Z_15 ));
    InMux I__12134 (
            .O(N__50560),
            .I(N__50557));
    LocalMux I__12133 (
            .O(N__50557),
            .I(\ALU.r0_12_prm_8_14_s1_c_RNOZ0Z_1 ));
    InMux I__12132 (
            .O(N__50554),
            .I(N__50551));
    LocalMux I__12131 (
            .O(N__50551),
            .I(op_i_0));
    InMux I__12130 (
            .O(N__50548),
            .I(N__50544));
    InMux I__12129 (
            .O(N__50547),
            .I(N__50541));
    LocalMux I__12128 (
            .O(N__50544),
            .I(N__50538));
    LocalMux I__12127 (
            .O(N__50541),
            .I(N__50533));
    Span4Mux_h I__12126 (
            .O(N__50538),
            .I(N__50533));
    Span4Mux_v I__12125 (
            .O(N__50533),
            .I(N__50530));
    Span4Mux_h I__12124 (
            .O(N__50530),
            .I(N__50527));
    Odrv4 I__12123 (
            .O(N__50527),
            .I(\ALU.un2_addsub_cry_0_c_RNIJPSHDZ0 ));
    CascadeMux I__12122 (
            .O(N__50524),
            .I(N__50521));
    InMux I__12121 (
            .O(N__50521),
            .I(N__50518));
    LocalMux I__12120 (
            .O(N__50518),
            .I(N__50515));
    Span4Mux_h I__12119 (
            .O(N__50515),
            .I(N__50512));
    Odrv4 I__12118 (
            .O(N__50512),
            .I(\ALU.r0_12_prm_2_1_c_RNOZ0 ));
    InMux I__12117 (
            .O(N__50509),
            .I(op_1_cry_1));
    InMux I__12116 (
            .O(N__50506),
            .I(op_1_cry_2));
    InMux I__12115 (
            .O(N__50503),
            .I(op_1_cry_3));
    CascadeMux I__12114 (
            .O(N__50500),
            .I(N__50494));
    CascadeMux I__12113 (
            .O(N__50499),
            .I(N__50490));
    CascadeMux I__12112 (
            .O(N__50498),
            .I(N__50486));
    InMux I__12111 (
            .O(N__50497),
            .I(N__50467));
    InMux I__12110 (
            .O(N__50494),
            .I(N__50467));
    InMux I__12109 (
            .O(N__50493),
            .I(N__50467));
    InMux I__12108 (
            .O(N__50490),
            .I(N__50467));
    InMux I__12107 (
            .O(N__50489),
            .I(N__50467));
    InMux I__12106 (
            .O(N__50486),
            .I(N__50467));
    InMux I__12105 (
            .O(N__50485),
            .I(N__50467));
    InMux I__12104 (
            .O(N__50484),
            .I(N__50467));
    LocalMux I__12103 (
            .O(N__50467),
            .I(N__50463));
    InMux I__12102 (
            .O(N__50466),
            .I(N__50458));
    Span4Mux_v I__12101 (
            .O(N__50463),
            .I(N__50455));
    InMux I__12100 (
            .O(N__50462),
            .I(N__50450));
    InMux I__12099 (
            .O(N__50461),
            .I(N__50450));
    LocalMux I__12098 (
            .O(N__50458),
            .I(yZ0Z_0));
    Odrv4 I__12097 (
            .O(N__50455),
            .I(yZ0Z_0));
    LocalMux I__12096 (
            .O(N__50450),
            .I(yZ0Z_0));
    InMux I__12095 (
            .O(N__50443),
            .I(N__50419));
    InMux I__12094 (
            .O(N__50442),
            .I(N__50419));
    InMux I__12093 (
            .O(N__50441),
            .I(N__50419));
    InMux I__12092 (
            .O(N__50440),
            .I(N__50419));
    InMux I__12091 (
            .O(N__50439),
            .I(N__50419));
    InMux I__12090 (
            .O(N__50438),
            .I(N__50419));
    InMux I__12089 (
            .O(N__50437),
            .I(N__50419));
    InMux I__12088 (
            .O(N__50436),
            .I(N__50419));
    LocalMux I__12087 (
            .O(N__50419),
            .I(N__50416));
    Span4Mux_v I__12086 (
            .O(N__50416),
            .I(N__50413));
    Span4Mux_v I__12085 (
            .O(N__50413),
            .I(N__50408));
    InMux I__12084 (
            .O(N__50412),
            .I(N__50403));
    InMux I__12083 (
            .O(N__50411),
            .I(N__50403));
    Odrv4 I__12082 (
            .O(N__50408),
            .I(yZ0Z_1));
    LocalMux I__12081 (
            .O(N__50403),
            .I(yZ0Z_1));
    InMux I__12080 (
            .O(N__50398),
            .I(N__50395));
    LocalMux I__12079 (
            .O(N__50395),
            .I(N__50392));
    Odrv4 I__12078 (
            .O(N__50392),
            .I(TXbufferZ0Z_7));
    InMux I__12077 (
            .O(N__50389),
            .I(N__50386));
    LocalMux I__12076 (
            .O(N__50386),
            .I(N__50383));
    Span4Mux_v I__12075 (
            .O(N__50383),
            .I(N__50380));
    Span4Mux_h I__12074 (
            .O(N__50380),
            .I(N__50377));
    Span4Mux_h I__12073 (
            .O(N__50377),
            .I(N__50374));
    Odrv4 I__12072 (
            .O(N__50374),
            .I(TXbufferZ0Z_1));
    InMux I__12071 (
            .O(N__50371),
            .I(N__50368));
    LocalMux I__12070 (
            .O(N__50368),
            .I(N__50365));
    Span4Mux_h I__12069 (
            .O(N__50365),
            .I(N__50362));
    Span4Mux_h I__12068 (
            .O(N__50362),
            .I(N__50359));
    Span4Mux_h I__12067 (
            .O(N__50359),
            .I(N__50356));
    Span4Mux_v I__12066 (
            .O(N__50356),
            .I(N__50353));
    Odrv4 I__12065 (
            .O(N__50353),
            .I(TXbufferZ0Z_2));
    InMux I__12064 (
            .O(N__50350),
            .I(N__50347));
    LocalMux I__12063 (
            .O(N__50347),
            .I(\FTDI.TXshiftZ0Z_2 ));
    InMux I__12062 (
            .O(N__50344),
            .I(N__50341));
    LocalMux I__12061 (
            .O(N__50341),
            .I(N__50338));
    Sp12to4 I__12060 (
            .O(N__50338),
            .I(N__50335));
    Span12Mux_s11_v I__12059 (
            .O(N__50335),
            .I(N__50332));
    Span12Mux_h I__12058 (
            .O(N__50332),
            .I(N__50329));
    Odrv12 I__12057 (
            .O(N__50329),
            .I(TXbufferZ0Z_4));
    InMux I__12056 (
            .O(N__50326),
            .I(N__50323));
    LocalMux I__12055 (
            .O(N__50323),
            .I(\FTDI.TXshiftZ0Z_4 ));
    InMux I__12054 (
            .O(N__50320),
            .I(N__50317));
    LocalMux I__12053 (
            .O(N__50317),
            .I(N__50314));
    Span12Mux_h I__12052 (
            .O(N__50314),
            .I(N__50311));
    Span12Mux_v I__12051 (
            .O(N__50311),
            .I(N__50308));
    Span12Mux_h I__12050 (
            .O(N__50308),
            .I(N__50305));
    Odrv12 I__12049 (
            .O(N__50305),
            .I(TXbufferZ0Z_3));
    InMux I__12048 (
            .O(N__50302),
            .I(N__50299));
    LocalMux I__12047 (
            .O(N__50299),
            .I(\FTDI.TXshiftZ0Z_3 ));
    InMux I__12046 (
            .O(N__50296),
            .I(N__50293));
    LocalMux I__12045 (
            .O(N__50293),
            .I(N__50290));
    Odrv4 I__12044 (
            .O(N__50290),
            .I(\FTDI.TXshiftZ0Z_7 ));
    InMux I__12043 (
            .O(N__50287),
            .I(N__50284));
    LocalMux I__12042 (
            .O(N__50284),
            .I(N__50281));
    Span12Mux_v I__12041 (
            .O(N__50281),
            .I(N__50278));
    Span12Mux_h I__12040 (
            .O(N__50278),
            .I(N__50275));
    Odrv12 I__12039 (
            .O(N__50275),
            .I(TXbufferZ0Z_6));
    InMux I__12038 (
            .O(N__50272),
            .I(N__50269));
    LocalMux I__12037 (
            .O(N__50269),
            .I(\FTDI.TXshiftZ0Z_6 ));
    InMux I__12036 (
            .O(N__50266),
            .I(N__50263));
    LocalMux I__12035 (
            .O(N__50263),
            .I(N__50260));
    Span4Mux_v I__12034 (
            .O(N__50260),
            .I(N__50257));
    Span4Mux_h I__12033 (
            .O(N__50257),
            .I(N__50254));
    Span4Mux_h I__12032 (
            .O(N__50254),
            .I(N__50251));
    Odrv4 I__12031 (
            .O(N__50251),
            .I(TXbufferZ0Z_5));
    InMux I__12030 (
            .O(N__50248),
            .I(N__50245));
    LocalMux I__12029 (
            .O(N__50245),
            .I(\FTDI.TXshiftZ0Z_5 ));
    InMux I__12028 (
            .O(N__50242),
            .I(N__50239));
    LocalMux I__12027 (
            .O(N__50239),
            .I(\ALU.r0_12_prm_1_3_c_RNOZ0 ));
    CascadeMux I__12026 (
            .O(N__50236),
            .I(N__50233));
    InMux I__12025 (
            .O(N__50233),
            .I(N__50229));
    InMux I__12024 (
            .O(N__50232),
            .I(N__50226));
    LocalMux I__12023 (
            .O(N__50229),
            .I(N__50223));
    LocalMux I__12022 (
            .O(N__50226),
            .I(N__50220));
    Span4Mux_v I__12021 (
            .O(N__50223),
            .I(N__50217));
    Span4Mux_v I__12020 (
            .O(N__50220),
            .I(N__50214));
    Span4Mux_h I__12019 (
            .O(N__50217),
            .I(N__50211));
    Span4Mux_h I__12018 (
            .O(N__50214),
            .I(N__50208));
    Odrv4 I__12017 (
            .O(N__50211),
            .I(\ALU.un9_addsub_cry_2_c_RNIOR8AJZ0 ));
    Odrv4 I__12016 (
            .O(N__50208),
            .I(\ALU.un9_addsub_cry_2_c_RNIOR8AJZ0 ));
    InMux I__12015 (
            .O(N__50203),
            .I(\ALU.r0_12_3 ));
    InMux I__12014 (
            .O(N__50200),
            .I(N__50196));
    InMux I__12013 (
            .O(N__50199),
            .I(N__50193));
    LocalMux I__12012 (
            .O(N__50196),
            .I(N__50189));
    LocalMux I__12011 (
            .O(N__50193),
            .I(N__50185));
    InMux I__12010 (
            .O(N__50192),
            .I(N__50182));
    Span4Mux_h I__12009 (
            .O(N__50189),
            .I(N__50179));
    InMux I__12008 (
            .O(N__50188),
            .I(N__50176));
    Span4Mux_v I__12007 (
            .O(N__50185),
            .I(N__50172));
    LocalMux I__12006 (
            .O(N__50182),
            .I(N__50168));
    Span4Mux_h I__12005 (
            .O(N__50179),
            .I(N__50163));
    LocalMux I__12004 (
            .O(N__50176),
            .I(N__50163));
    InMux I__12003 (
            .O(N__50175),
            .I(N__50160));
    Span4Mux_h I__12002 (
            .O(N__50172),
            .I(N__50156));
    InMux I__12001 (
            .O(N__50171),
            .I(N__50153));
    Span4Mux_h I__12000 (
            .O(N__50168),
            .I(N__50150));
    Span4Mux_v I__11999 (
            .O(N__50163),
            .I(N__50145));
    LocalMux I__11998 (
            .O(N__50160),
            .I(N__50145));
    InMux I__11997 (
            .O(N__50159),
            .I(N__50142));
    Span4Mux_h I__11996 (
            .O(N__50156),
            .I(N__50137));
    LocalMux I__11995 (
            .O(N__50153),
            .I(N__50137));
    Span4Mux_h I__11994 (
            .O(N__50150),
            .I(N__50129));
    Span4Mux_h I__11993 (
            .O(N__50145),
            .I(N__50129));
    LocalMux I__11992 (
            .O(N__50142),
            .I(N__50129));
    Span4Mux_h I__11991 (
            .O(N__50137),
            .I(N__50126));
    InMux I__11990 (
            .O(N__50136),
            .I(N__50123));
    Span4Mux_h I__11989 (
            .O(N__50129),
            .I(N__50120));
    Sp12to4 I__11988 (
            .O(N__50126),
            .I(N__50115));
    LocalMux I__11987 (
            .O(N__50123),
            .I(N__50115));
    Odrv4 I__11986 (
            .O(N__50120),
            .I(\ALU.r0_12_3_THRU_CO ));
    Odrv12 I__11985 (
            .O(N__50115),
            .I(\ALU.r0_12_3_THRU_CO ));
    CascadeMux I__11984 (
            .O(N__50110),
            .I(N__50107));
    InMux I__11983 (
            .O(N__50107),
            .I(N__50104));
    LocalMux I__11982 (
            .O(N__50104),
            .I(N__50100));
    InMux I__11981 (
            .O(N__50103),
            .I(N__50097));
    Span4Mux_h I__11980 (
            .O(N__50100),
            .I(N__50094));
    LocalMux I__11979 (
            .O(N__50097),
            .I(N__50091));
    Span4Mux_h I__11978 (
            .O(N__50094),
            .I(N__50088));
    Span4Mux_h I__11977 (
            .O(N__50091),
            .I(N__50085));
    Span4Mux_h I__11976 (
            .O(N__50088),
            .I(N__50082));
    Span4Mux_h I__11975 (
            .O(N__50085),
            .I(N__50079));
    Odrv4 I__11974 (
            .O(N__50082),
            .I(\ALU.un2_addsub_cry_2_c_RNI3K9SGZ0 ));
    Odrv4 I__11973 (
            .O(N__50079),
            .I(\ALU.un2_addsub_cry_2_c_RNI3K9SGZ0 ));
    InMux I__11972 (
            .O(N__50074),
            .I(N__50071));
    LocalMux I__11971 (
            .O(N__50071),
            .I(\ALU.r0_12_prm_2_3_c_RNOZ0 ));
    InMux I__11970 (
            .O(N__50068),
            .I(N__50065));
    LocalMux I__11969 (
            .O(N__50065),
            .I(\ALU.r0_12_prm_3_3_c_RNOZ0 ));
    InMux I__11968 (
            .O(N__50062),
            .I(N__50056));
    InMux I__11967 (
            .O(N__50061),
            .I(N__50056));
    LocalMux I__11966 (
            .O(N__50056),
            .I(N__50053));
    Span4Mux_h I__11965 (
            .O(N__50053),
            .I(N__50049));
    InMux I__11964 (
            .O(N__50052),
            .I(N__50046));
    Span4Mux_h I__11963 (
            .O(N__50049),
            .I(N__50041));
    LocalMux I__11962 (
            .O(N__50046),
            .I(N__50041));
    Span4Mux_h I__11961 (
            .O(N__50041),
            .I(N__50038));
    Odrv4 I__11960 (
            .O(N__50038),
            .I(\ALU.madd_axb_2 ));
    CascadeMux I__11959 (
            .O(N__50035),
            .I(N__50032));
    InMux I__11958 (
            .O(N__50032),
            .I(N__50026));
    InMux I__11957 (
            .O(N__50031),
            .I(N__50026));
    LocalMux I__11956 (
            .O(N__50026),
            .I(N__50023));
    Span4Mux_h I__11955 (
            .O(N__50023),
            .I(N__50020));
    Span4Mux_h I__11954 (
            .O(N__50020),
            .I(N__50017));
    Span4Mux_h I__11953 (
            .O(N__50017),
            .I(N__50014));
    Odrv4 I__11952 (
            .O(N__50014),
            .I(\ALU.madd_cry_1_THRU_CO ));
    CascadeMux I__11951 (
            .O(N__50011),
            .I(N__50008));
    InMux I__11950 (
            .O(N__50008),
            .I(N__50005));
    LocalMux I__11949 (
            .O(N__50005),
            .I(\ALU.mult_3 ));
    InMux I__11948 (
            .O(N__50002),
            .I(N__49999));
    LocalMux I__11947 (
            .O(N__49999),
            .I(N__49996));
    Span12Mux_v I__11946 (
            .O(N__49996),
            .I(N__49993));
    Span12Mux_h I__11945 (
            .O(N__49993),
            .I(N__49990));
    Odrv12 I__11944 (
            .O(N__49990),
            .I(TXbuffer_RNO_1Z0Z_7));
    InMux I__11943 (
            .O(N__49987),
            .I(N__49984));
    LocalMux I__11942 (
            .O(N__49984),
            .I(N__49981));
    Odrv12 I__11941 (
            .O(N__49981),
            .I(TXbuffer_RNO_0Z0Z_7));
    CascadeMux I__11940 (
            .O(N__49978),
            .I(N__49975));
    InMux I__11939 (
            .O(N__49975),
            .I(N__49971));
    CascadeMux I__11938 (
            .O(N__49974),
            .I(N__49964));
    LocalMux I__11937 (
            .O(N__49971),
            .I(N__49961));
    InMux I__11936 (
            .O(N__49970),
            .I(N__49958));
    InMux I__11935 (
            .O(N__49969),
            .I(N__49955));
    InMux I__11934 (
            .O(N__49968),
            .I(N__49952));
    CascadeMux I__11933 (
            .O(N__49967),
            .I(N__49949));
    InMux I__11932 (
            .O(N__49964),
            .I(N__49946));
    Span4Mux_v I__11931 (
            .O(N__49961),
            .I(N__49941));
    LocalMux I__11930 (
            .O(N__49958),
            .I(N__49941));
    LocalMux I__11929 (
            .O(N__49955),
            .I(N__49933));
    LocalMux I__11928 (
            .O(N__49952),
            .I(N__49929));
    InMux I__11927 (
            .O(N__49949),
            .I(N__49926));
    LocalMux I__11926 (
            .O(N__49946),
            .I(N__49922));
    Span4Mux_v I__11925 (
            .O(N__49941),
            .I(N__49919));
    InMux I__11924 (
            .O(N__49940),
            .I(N__49916));
    InMux I__11923 (
            .O(N__49939),
            .I(N__49911));
    InMux I__11922 (
            .O(N__49938),
            .I(N__49911));
    InMux I__11921 (
            .O(N__49937),
            .I(N__49906));
    InMux I__11920 (
            .O(N__49936),
            .I(N__49906));
    Span4Mux_v I__11919 (
            .O(N__49933),
            .I(N__49903));
    InMux I__11918 (
            .O(N__49932),
            .I(N__49899));
    Span4Mux_v I__11917 (
            .O(N__49929),
            .I(N__49896));
    LocalMux I__11916 (
            .O(N__49926),
            .I(N__49893));
    InMux I__11915 (
            .O(N__49925),
            .I(N__49890));
    Span12Mux_h I__11914 (
            .O(N__49922),
            .I(N__49881));
    Sp12to4 I__11913 (
            .O(N__49919),
            .I(N__49881));
    LocalMux I__11912 (
            .O(N__49916),
            .I(N__49881));
    LocalMux I__11911 (
            .O(N__49911),
            .I(N__49874));
    LocalMux I__11910 (
            .O(N__49906),
            .I(N__49874));
    Span4Mux_h I__11909 (
            .O(N__49903),
            .I(N__49874));
    InMux I__11908 (
            .O(N__49902),
            .I(N__49871));
    LocalMux I__11907 (
            .O(N__49899),
            .I(N__49868));
    Span4Mux_h I__11906 (
            .O(N__49896),
            .I(N__49865));
    Span4Mux_h I__11905 (
            .O(N__49893),
            .I(N__49860));
    LocalMux I__11904 (
            .O(N__49890),
            .I(N__49860));
    InMux I__11903 (
            .O(N__49889),
            .I(N__49857));
    InMux I__11902 (
            .O(N__49888),
            .I(N__49854));
    Span12Mux_h I__11901 (
            .O(N__49881),
            .I(N__49850));
    Span4Mux_v I__11900 (
            .O(N__49874),
            .I(N__49847));
    LocalMux I__11899 (
            .O(N__49871),
            .I(N__49842));
    Span4Mux_v I__11898 (
            .O(N__49868),
            .I(N__49842));
    Span4Mux_v I__11897 (
            .O(N__49865),
            .I(N__49837));
    Span4Mux_h I__11896 (
            .O(N__49860),
            .I(N__49837));
    LocalMux I__11895 (
            .O(N__49857),
            .I(N__49832));
    LocalMux I__11894 (
            .O(N__49854),
            .I(N__49832));
    InMux I__11893 (
            .O(N__49853),
            .I(N__49829));
    Odrv12 I__11892 (
            .O(N__49850),
            .I(clkdivZ0Z_4));
    Odrv4 I__11891 (
            .O(N__49847),
            .I(clkdivZ0Z_4));
    Odrv4 I__11890 (
            .O(N__49842),
            .I(clkdivZ0Z_4));
    Odrv4 I__11889 (
            .O(N__49837),
            .I(clkdivZ0Z_4));
    Odrv4 I__11888 (
            .O(N__49832),
            .I(clkdivZ0Z_4));
    LocalMux I__11887 (
            .O(N__49829),
            .I(clkdivZ0Z_4));
    InMux I__11886 (
            .O(N__49816),
            .I(N__49813));
    LocalMux I__11885 (
            .O(N__49813),
            .I(N__49810));
    Odrv12 I__11884 (
            .O(N__49810),
            .I(TXbuffer_18_15_ns_1_7));
    CascadeMux I__11883 (
            .O(N__49807),
            .I(N__49804));
    InMux I__11882 (
            .O(N__49804),
            .I(N__49797));
    CascadeMux I__11881 (
            .O(N__49803),
            .I(N__49792));
    CascadeMux I__11880 (
            .O(N__49802),
            .I(N__49788));
    CascadeMux I__11879 (
            .O(N__49801),
            .I(N__49784));
    CascadeMux I__11878 (
            .O(N__49800),
            .I(N__49781));
    LocalMux I__11877 (
            .O(N__49797),
            .I(N__49778));
    InMux I__11876 (
            .O(N__49796),
            .I(N__49761));
    InMux I__11875 (
            .O(N__49795),
            .I(N__49761));
    InMux I__11874 (
            .O(N__49792),
            .I(N__49761));
    InMux I__11873 (
            .O(N__49791),
            .I(N__49761));
    InMux I__11872 (
            .O(N__49788),
            .I(N__49761));
    InMux I__11871 (
            .O(N__49787),
            .I(N__49761));
    InMux I__11870 (
            .O(N__49784),
            .I(N__49761));
    InMux I__11869 (
            .O(N__49781),
            .I(N__49761));
    Odrv4 I__11868 (
            .O(N__49778),
            .I(yZ0Z_2));
    LocalMux I__11867 (
            .O(N__49761),
            .I(yZ0Z_2));
    CEMux I__11866 (
            .O(N__49756),
            .I(N__49753));
    LocalMux I__11865 (
            .O(N__49753),
            .I(N__49750));
    Span4Mux_v I__11864 (
            .O(N__49750),
            .I(N__49747));
    Span4Mux_h I__11863 (
            .O(N__49747),
            .I(N__49743));
    CEMux I__11862 (
            .O(N__49746),
            .I(N__49740));
    Span4Mux_h I__11861 (
            .O(N__49743),
            .I(N__49734));
    LocalMux I__11860 (
            .O(N__49740),
            .I(N__49734));
    CEMux I__11859 (
            .O(N__49739),
            .I(N__49727));
    Span4Mux_v I__11858 (
            .O(N__49734),
            .I(N__49723));
    CEMux I__11857 (
            .O(N__49733),
            .I(N__49720));
    CEMux I__11856 (
            .O(N__49732),
            .I(N__49713));
    CEMux I__11855 (
            .O(N__49731),
            .I(N__49710));
    CEMux I__11854 (
            .O(N__49730),
            .I(N__49707));
    LocalMux I__11853 (
            .O(N__49727),
            .I(N__49704));
    CEMux I__11852 (
            .O(N__49726),
            .I(N__49701));
    Span4Mux_h I__11851 (
            .O(N__49723),
            .I(N__49698));
    LocalMux I__11850 (
            .O(N__49720),
            .I(N__49695));
    CEMux I__11849 (
            .O(N__49719),
            .I(N__49692));
    CEMux I__11848 (
            .O(N__49718),
            .I(N__49689));
    CEMux I__11847 (
            .O(N__49717),
            .I(N__49686));
    CEMux I__11846 (
            .O(N__49716),
            .I(N__49682));
    LocalMux I__11845 (
            .O(N__49713),
            .I(N__49679));
    LocalMux I__11844 (
            .O(N__49710),
            .I(N__49676));
    LocalMux I__11843 (
            .O(N__49707),
            .I(N__49673));
    Span4Mux_v I__11842 (
            .O(N__49704),
            .I(N__49670));
    LocalMux I__11841 (
            .O(N__49701),
            .I(N__49667));
    Span4Mux_s0_h I__11840 (
            .O(N__49698),
            .I(N__49664));
    Span4Mux_h I__11839 (
            .O(N__49695),
            .I(N__49661));
    LocalMux I__11838 (
            .O(N__49692),
            .I(N__49658));
    LocalMux I__11837 (
            .O(N__49689),
            .I(N__49655));
    LocalMux I__11836 (
            .O(N__49686),
            .I(N__49652));
    CEMux I__11835 (
            .O(N__49685),
            .I(N__49649));
    LocalMux I__11834 (
            .O(N__49682),
            .I(N__49646));
    Span4Mux_v I__11833 (
            .O(N__49679),
            .I(N__49643));
    Span4Mux_v I__11832 (
            .O(N__49676),
            .I(N__49640));
    Span4Mux_h I__11831 (
            .O(N__49673),
            .I(N__49637));
    Span4Mux_s3_h I__11830 (
            .O(N__49670),
            .I(N__49634));
    Span4Mux_h I__11829 (
            .O(N__49667),
            .I(N__49631));
    Span4Mux_v I__11828 (
            .O(N__49664),
            .I(N__49626));
    Span4Mux_s0_h I__11827 (
            .O(N__49661),
            .I(N__49626));
    Span4Mux_v I__11826 (
            .O(N__49658),
            .I(N__49619));
    Span4Mux_v I__11825 (
            .O(N__49655),
            .I(N__49619));
    Span4Mux_h I__11824 (
            .O(N__49652),
            .I(N__49619));
    LocalMux I__11823 (
            .O(N__49649),
            .I(N__49616));
    Span4Mux_v I__11822 (
            .O(N__49646),
            .I(N__49609));
    Span4Mux_h I__11821 (
            .O(N__49643),
            .I(N__49609));
    Span4Mux_h I__11820 (
            .O(N__49640),
            .I(N__49609));
    Span4Mux_h I__11819 (
            .O(N__49637),
            .I(N__49606));
    Span4Mux_h I__11818 (
            .O(N__49634),
            .I(N__49603));
    Span4Mux_h I__11817 (
            .O(N__49631),
            .I(N__49600));
    Span4Mux_v I__11816 (
            .O(N__49626),
            .I(N__49597));
    Span4Mux_h I__11815 (
            .O(N__49619),
            .I(N__49594));
    Span4Mux_h I__11814 (
            .O(N__49616),
            .I(N__49591));
    Span4Mux_h I__11813 (
            .O(N__49609),
            .I(N__49588));
    Span4Mux_v I__11812 (
            .O(N__49606),
            .I(N__49583));
    Span4Mux_h I__11811 (
            .O(N__49603),
            .I(N__49583));
    Sp12to4 I__11810 (
            .O(N__49600),
            .I(N__49580));
    Sp12to4 I__11809 (
            .O(N__49597),
            .I(N__49577));
    Span4Mux_h I__11808 (
            .O(N__49594),
            .I(N__49574));
    Span4Mux_h I__11807 (
            .O(N__49591),
            .I(N__49569));
    Span4Mux_h I__11806 (
            .O(N__49588),
            .I(N__49569));
    Span4Mux_h I__11805 (
            .O(N__49583),
            .I(N__49566));
    Span12Mux_v I__11804 (
            .O(N__49580),
            .I(N__49561));
    Span12Mux_s11_h I__11803 (
            .O(N__49577),
            .I(N__49561));
    Span4Mux_v I__11802 (
            .O(N__49574),
            .I(N__49558));
    Odrv4 I__11801 (
            .O(N__49569),
            .I(\ALU.un1_yindexZ0Z_8 ));
    Odrv4 I__11800 (
            .O(N__49566),
            .I(\ALU.un1_yindexZ0Z_8 ));
    Odrv12 I__11799 (
            .O(N__49561),
            .I(\ALU.un1_yindexZ0Z_8 ));
    Odrv4 I__11798 (
            .O(N__49558),
            .I(\ALU.un1_yindexZ0Z_8 ));
    CascadeMux I__11797 (
            .O(N__49549),
            .I(N__49546));
    InMux I__11796 (
            .O(N__49546),
            .I(N__49542));
    InMux I__11795 (
            .O(N__49545),
            .I(N__49539));
    LocalMux I__11794 (
            .O(N__49542),
            .I(\ALU.rshift_3 ));
    LocalMux I__11793 (
            .O(N__49539),
            .I(\ALU.rshift_3 ));
    InMux I__11792 (
            .O(N__49534),
            .I(N__49531));
    LocalMux I__11791 (
            .O(N__49531),
            .I(N__49528));
    Span4Mux_h I__11790 (
            .O(N__49528),
            .I(N__49525));
    Odrv4 I__11789 (
            .O(N__49525),
            .I(\ALU.r0_12_prm_8_3_c_RNOZ0 ));
    InMux I__11788 (
            .O(N__49522),
            .I(N__49519));
    LocalMux I__11787 (
            .O(N__49519),
            .I(\ALU.r0_12_prm_7_3_c_RNOZ0 ));
    CascadeMux I__11786 (
            .O(N__49516),
            .I(N__49513));
    InMux I__11785 (
            .O(N__49513),
            .I(N__49509));
    InMux I__11784 (
            .O(N__49512),
            .I(N__49506));
    LocalMux I__11783 (
            .O(N__49509),
            .I(N__49501));
    LocalMux I__11782 (
            .O(N__49506),
            .I(N__49501));
    Span4Mux_v I__11781 (
            .O(N__49501),
            .I(N__49498));
    Span4Mux_h I__11780 (
            .O(N__49498),
            .I(N__49495));
    Odrv4 I__11779 (
            .O(N__49495),
            .I(\ALU.a3_b_3 ));
    InMux I__11778 (
            .O(N__49492),
            .I(N__49489));
    LocalMux I__11777 (
            .O(N__49489),
            .I(N__49486));
    Span12Mux_h I__11776 (
            .O(N__49486),
            .I(N__49483));
    Odrv12 I__11775 (
            .O(N__49483),
            .I(\ALU.un14_log_0_i_3 ));
    CascadeMux I__11774 (
            .O(N__49480),
            .I(N__49477));
    InMux I__11773 (
            .O(N__49477),
            .I(N__49474));
    LocalMux I__11772 (
            .O(N__49474),
            .I(N__49471));
    Span12Mux_h I__11771 (
            .O(N__49471),
            .I(N__49468));
    Odrv12 I__11770 (
            .O(N__49468),
            .I(\ALU.r0_12_prm_6_3_c_RNOZ0 ));
    InMux I__11769 (
            .O(N__49465),
            .I(N__49462));
    LocalMux I__11768 (
            .O(N__49462),
            .I(\ALU.r0_12_prm_5_3_c_RNOZ0 ));
    CascadeMux I__11767 (
            .O(N__49459),
            .I(N__49456));
    InMux I__11766 (
            .O(N__49456),
            .I(N__49453));
    LocalMux I__11765 (
            .O(N__49453),
            .I(N__49450));
    Span4Mux_h I__11764 (
            .O(N__49450),
            .I(N__49447));
    Odrv4 I__11763 (
            .O(N__49447),
            .I(\ALU.r0_12_prm_5_3_c_RNOZ0Z_0 ));
    InMux I__11762 (
            .O(N__49444),
            .I(N__49441));
    LocalMux I__11761 (
            .O(N__49441),
            .I(N__49438));
    Span4Mux_v I__11760 (
            .O(N__49438),
            .I(N__49435));
    Span4Mux_v I__11759 (
            .O(N__49435),
            .I(N__49432));
    Span4Mux_h I__11758 (
            .O(N__49432),
            .I(N__49429));
    Odrv4 I__11757 (
            .O(N__49429),
            .I(\ALU.r4_RNIUH636Z0Z_3 ));
    InMux I__11756 (
            .O(N__49426),
            .I(N__49420));
    InMux I__11755 (
            .O(N__49425),
            .I(N__49413));
    InMux I__11754 (
            .O(N__49424),
            .I(N__49409));
    InMux I__11753 (
            .O(N__49423),
            .I(N__49405));
    LocalMux I__11752 (
            .O(N__49420),
            .I(N__49402));
    InMux I__11751 (
            .O(N__49419),
            .I(N__49399));
    InMux I__11750 (
            .O(N__49418),
            .I(N__49394));
    InMux I__11749 (
            .O(N__49417),
            .I(N__49390));
    InMux I__11748 (
            .O(N__49416),
            .I(N__49387));
    LocalMux I__11747 (
            .O(N__49413),
            .I(N__49384));
    InMux I__11746 (
            .O(N__49412),
            .I(N__49381));
    LocalMux I__11745 (
            .O(N__49409),
            .I(N__49378));
    InMux I__11744 (
            .O(N__49408),
            .I(N__49375));
    LocalMux I__11743 (
            .O(N__49405),
            .I(N__49372));
    Span4Mux_h I__11742 (
            .O(N__49402),
            .I(N__49367));
    LocalMux I__11741 (
            .O(N__49399),
            .I(N__49367));
    InMux I__11740 (
            .O(N__49398),
            .I(N__49357));
    InMux I__11739 (
            .O(N__49397),
            .I(N__49354));
    LocalMux I__11738 (
            .O(N__49394),
            .I(N__49345));
    InMux I__11737 (
            .O(N__49393),
            .I(N__49342));
    LocalMux I__11736 (
            .O(N__49390),
            .I(N__49338));
    LocalMux I__11735 (
            .O(N__49387),
            .I(N__49335));
    Span4Mux_v I__11734 (
            .O(N__49384),
            .I(N__49326));
    LocalMux I__11733 (
            .O(N__49381),
            .I(N__49326));
    Span4Mux_h I__11732 (
            .O(N__49378),
            .I(N__49326));
    LocalMux I__11731 (
            .O(N__49375),
            .I(N__49326));
    Span4Mux_h I__11730 (
            .O(N__49372),
            .I(N__49319));
    Span4Mux_v I__11729 (
            .O(N__49367),
            .I(N__49319));
    InMux I__11728 (
            .O(N__49366),
            .I(N__49316));
    InMux I__11727 (
            .O(N__49365),
            .I(N__49309));
    InMux I__11726 (
            .O(N__49364),
            .I(N__49309));
    InMux I__11725 (
            .O(N__49363),
            .I(N__49309));
    InMux I__11724 (
            .O(N__49362),
            .I(N__49306));
    InMux I__11723 (
            .O(N__49361),
            .I(N__49303));
    InMux I__11722 (
            .O(N__49360),
            .I(N__49300));
    LocalMux I__11721 (
            .O(N__49357),
            .I(N__49297));
    LocalMux I__11720 (
            .O(N__49354),
            .I(N__49294));
    InMux I__11719 (
            .O(N__49353),
            .I(N__49289));
    InMux I__11718 (
            .O(N__49352),
            .I(N__49289));
    InMux I__11717 (
            .O(N__49351),
            .I(N__49283));
    InMux I__11716 (
            .O(N__49350),
            .I(N__49283));
    InMux I__11715 (
            .O(N__49349),
            .I(N__49278));
    InMux I__11714 (
            .O(N__49348),
            .I(N__49278));
    Span4Mux_v I__11713 (
            .O(N__49345),
            .I(N__49274));
    LocalMux I__11712 (
            .O(N__49342),
            .I(N__49271));
    InMux I__11711 (
            .O(N__49341),
            .I(N__49268));
    Span4Mux_v I__11710 (
            .O(N__49338),
            .I(N__49265));
    Span4Mux_h I__11709 (
            .O(N__49335),
            .I(N__49260));
    Span4Mux_v I__11708 (
            .O(N__49326),
            .I(N__49260));
    InMux I__11707 (
            .O(N__49325),
            .I(N__49255));
    InMux I__11706 (
            .O(N__49324),
            .I(N__49255));
    Span4Mux_h I__11705 (
            .O(N__49319),
            .I(N__49250));
    LocalMux I__11704 (
            .O(N__49316),
            .I(N__49247));
    LocalMux I__11703 (
            .O(N__49309),
            .I(N__49242));
    LocalMux I__11702 (
            .O(N__49306),
            .I(N__49242));
    LocalMux I__11701 (
            .O(N__49303),
            .I(N__49239));
    LocalMux I__11700 (
            .O(N__49300),
            .I(N__49227));
    Span4Mux_s0_v I__11699 (
            .O(N__49297),
            .I(N__49227));
    Span4Mux_v I__11698 (
            .O(N__49294),
            .I(N__49227));
    LocalMux I__11697 (
            .O(N__49289),
            .I(N__49227));
    InMux I__11696 (
            .O(N__49288),
            .I(N__49224));
    LocalMux I__11695 (
            .O(N__49283),
            .I(N__49219));
    LocalMux I__11694 (
            .O(N__49278),
            .I(N__49219));
    InMux I__11693 (
            .O(N__49277),
            .I(N__49216));
    Span4Mux_h I__11692 (
            .O(N__49274),
            .I(N__49213));
    Span12Mux_v I__11691 (
            .O(N__49271),
            .I(N__49202));
    LocalMux I__11690 (
            .O(N__49268),
            .I(N__49202));
    Sp12to4 I__11689 (
            .O(N__49265),
            .I(N__49202));
    Sp12to4 I__11688 (
            .O(N__49260),
            .I(N__49202));
    LocalMux I__11687 (
            .O(N__49255),
            .I(N__49202));
    InMux I__11686 (
            .O(N__49254),
            .I(N__49197));
    InMux I__11685 (
            .O(N__49253),
            .I(N__49197));
    Span4Mux_v I__11684 (
            .O(N__49250),
            .I(N__49192));
    Span4Mux_h I__11683 (
            .O(N__49247),
            .I(N__49192));
    Span4Mux_v I__11682 (
            .O(N__49242),
            .I(N__49187));
    Span4Mux_s3_v I__11681 (
            .O(N__49239),
            .I(N__49187));
    InMux I__11680 (
            .O(N__49238),
            .I(N__49184));
    InMux I__11679 (
            .O(N__49237),
            .I(N__49179));
    InMux I__11678 (
            .O(N__49236),
            .I(N__49179));
    Span4Mux_h I__11677 (
            .O(N__49227),
            .I(N__49170));
    LocalMux I__11676 (
            .O(N__49224),
            .I(N__49170));
    Span4Mux_h I__11675 (
            .O(N__49219),
            .I(N__49170));
    LocalMux I__11674 (
            .O(N__49216),
            .I(N__49170));
    Odrv4 I__11673 (
            .O(N__49213),
            .I(\ALU.a_3 ));
    Odrv12 I__11672 (
            .O(N__49202),
            .I(\ALU.a_3 ));
    LocalMux I__11671 (
            .O(N__49197),
            .I(\ALU.a_3 ));
    Odrv4 I__11670 (
            .O(N__49192),
            .I(\ALU.a_3 ));
    Odrv4 I__11669 (
            .O(N__49187),
            .I(\ALU.a_3 ));
    LocalMux I__11668 (
            .O(N__49184),
            .I(\ALU.a_3 ));
    LocalMux I__11667 (
            .O(N__49179),
            .I(\ALU.a_3 ));
    Odrv4 I__11666 (
            .O(N__49170),
            .I(\ALU.a_3 ));
    CascadeMux I__11665 (
            .O(N__49153),
            .I(N__49150));
    InMux I__11664 (
            .O(N__49150),
            .I(N__49147));
    LocalMux I__11663 (
            .O(N__49147),
            .I(N__49144));
    Odrv4 I__11662 (
            .O(N__49144),
            .I(\ALU.a_i_3 ));
    InMux I__11661 (
            .O(N__49141),
            .I(N__49137));
    InMux I__11660 (
            .O(N__49140),
            .I(N__49133));
    LocalMux I__11659 (
            .O(N__49137),
            .I(N__49129));
    InMux I__11658 (
            .O(N__49136),
            .I(N__49126));
    LocalMux I__11657 (
            .O(N__49133),
            .I(N__49123));
    InMux I__11656 (
            .O(N__49132),
            .I(N__49120));
    Span4Mux_h I__11655 (
            .O(N__49129),
            .I(N__49115));
    LocalMux I__11654 (
            .O(N__49126),
            .I(N__49115));
    Span4Mux_h I__11653 (
            .O(N__49123),
            .I(N__49108));
    LocalMux I__11652 (
            .O(N__49120),
            .I(N__49108));
    Span4Mux_h I__11651 (
            .O(N__49115),
            .I(N__49108));
    Odrv4 I__11650 (
            .O(N__49108),
            .I(\ALU.un2_addsub_cry_13_c_RNIR5I0EZ0 ));
    CascadeMux I__11649 (
            .O(N__49105),
            .I(N__49102));
    InMux I__11648 (
            .O(N__49102),
            .I(N__49099));
    LocalMux I__11647 (
            .O(N__49099),
            .I(\ALU.r0_12_prm_2_14_s1_c_RNOZ0 ));
    InMux I__11646 (
            .O(N__49096),
            .I(N__49093));
    LocalMux I__11645 (
            .O(N__49093),
            .I(N__49090));
    Span4Mux_v I__11644 (
            .O(N__49090),
            .I(N__49087));
    Odrv4 I__11643 (
            .O(N__49087),
            .I(\ALU.r0_12_prm_1_14_s1_c_RNOZ0 ));
    CascadeMux I__11642 (
            .O(N__49084),
            .I(N__49080));
    InMux I__11641 (
            .O(N__49083),
            .I(N__49077));
    InMux I__11640 (
            .O(N__49080),
            .I(N__49074));
    LocalMux I__11639 (
            .O(N__49077),
            .I(N__49070));
    LocalMux I__11638 (
            .O(N__49074),
            .I(N__49067));
    InMux I__11637 (
            .O(N__49073),
            .I(N__49064));
    Span4Mux_v I__11636 (
            .O(N__49070),
            .I(N__49061));
    Span4Mux_v I__11635 (
            .O(N__49067),
            .I(N__49058));
    LocalMux I__11634 (
            .O(N__49064),
            .I(N__49055));
    Span4Mux_h I__11633 (
            .O(N__49061),
            .I(N__49049));
    Span4Mux_h I__11632 (
            .O(N__49058),
            .I(N__49049));
    Span4Mux_v I__11631 (
            .O(N__49055),
            .I(N__49046));
    InMux I__11630 (
            .O(N__49054),
            .I(N__49043));
    Odrv4 I__11629 (
            .O(N__49049),
            .I(\ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9 ));
    Odrv4 I__11628 (
            .O(N__49046),
            .I(\ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9 ));
    LocalMux I__11627 (
            .O(N__49043),
            .I(\ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9 ));
    InMux I__11626 (
            .O(N__49036),
            .I(\ALU.r0_12_s1_14 ));
    InMux I__11625 (
            .O(N__49033),
            .I(N__49030));
    LocalMux I__11624 (
            .O(N__49030),
            .I(N__49027));
    Span4Mux_h I__11623 (
            .O(N__49027),
            .I(N__49024));
    Span4Mux_h I__11622 (
            .O(N__49024),
            .I(N__49021));
    Odrv4 I__11621 (
            .O(N__49021),
            .I(\ALU.r0_12_s1_14_THRU_CO ));
    CascadeMux I__11620 (
            .O(N__49018),
            .I(N__49009));
    InMux I__11619 (
            .O(N__49017),
            .I(N__49005));
    InMux I__11618 (
            .O(N__49016),
            .I(N__48995));
    InMux I__11617 (
            .O(N__49015),
            .I(N__48990));
    InMux I__11616 (
            .O(N__49014),
            .I(N__48990));
    InMux I__11615 (
            .O(N__49013),
            .I(N__48984));
    InMux I__11614 (
            .O(N__49012),
            .I(N__48980));
    InMux I__11613 (
            .O(N__49009),
            .I(N__48977));
    InMux I__11612 (
            .O(N__49008),
            .I(N__48974));
    LocalMux I__11611 (
            .O(N__49005),
            .I(N__48971));
    InMux I__11610 (
            .O(N__49004),
            .I(N__48968));
    InMux I__11609 (
            .O(N__49003),
            .I(N__48965));
    InMux I__11608 (
            .O(N__49002),
            .I(N__48962));
    InMux I__11607 (
            .O(N__49001),
            .I(N__48959));
    InMux I__11606 (
            .O(N__49000),
            .I(N__48956));
    InMux I__11605 (
            .O(N__48999),
            .I(N__48950));
    InMux I__11604 (
            .O(N__48998),
            .I(N__48950));
    LocalMux I__11603 (
            .O(N__48995),
            .I(N__48946));
    LocalMux I__11602 (
            .O(N__48990),
            .I(N__48940));
    InMux I__11601 (
            .O(N__48989),
            .I(N__48937));
    CascadeMux I__11600 (
            .O(N__48988),
            .I(N__48929));
    CascadeMux I__11599 (
            .O(N__48987),
            .I(N__48923));
    LocalMux I__11598 (
            .O(N__48984),
            .I(N__48917));
    InMux I__11597 (
            .O(N__48983),
            .I(N__48904));
    LocalMux I__11596 (
            .O(N__48980),
            .I(N__48901));
    LocalMux I__11595 (
            .O(N__48977),
            .I(N__48894));
    LocalMux I__11594 (
            .O(N__48974),
            .I(N__48894));
    Span4Mux_v I__11593 (
            .O(N__48971),
            .I(N__48894));
    LocalMux I__11592 (
            .O(N__48968),
            .I(N__48891));
    LocalMux I__11591 (
            .O(N__48965),
            .I(N__48888));
    LocalMux I__11590 (
            .O(N__48962),
            .I(N__48885));
    LocalMux I__11589 (
            .O(N__48959),
            .I(N__48880));
    LocalMux I__11588 (
            .O(N__48956),
            .I(N__48880));
    InMux I__11587 (
            .O(N__48955),
            .I(N__48877));
    LocalMux I__11586 (
            .O(N__48950),
            .I(N__48874));
    InMux I__11585 (
            .O(N__48949),
            .I(N__48871));
    Span4Mux_v I__11584 (
            .O(N__48946),
            .I(N__48867));
    InMux I__11583 (
            .O(N__48945),
            .I(N__48860));
    InMux I__11582 (
            .O(N__48944),
            .I(N__48860));
    InMux I__11581 (
            .O(N__48943),
            .I(N__48860));
    Span4Mux_s2_v I__11580 (
            .O(N__48940),
            .I(N__48855));
    LocalMux I__11579 (
            .O(N__48937),
            .I(N__48855));
    InMux I__11578 (
            .O(N__48936),
            .I(N__48846));
    InMux I__11577 (
            .O(N__48935),
            .I(N__48846));
    InMux I__11576 (
            .O(N__48934),
            .I(N__48846));
    InMux I__11575 (
            .O(N__48933),
            .I(N__48846));
    InMux I__11574 (
            .O(N__48932),
            .I(N__48839));
    InMux I__11573 (
            .O(N__48929),
            .I(N__48839));
    InMux I__11572 (
            .O(N__48928),
            .I(N__48839));
    InMux I__11571 (
            .O(N__48927),
            .I(N__48834));
    InMux I__11570 (
            .O(N__48926),
            .I(N__48834));
    InMux I__11569 (
            .O(N__48923),
            .I(N__48831));
    InMux I__11568 (
            .O(N__48922),
            .I(N__48827));
    InMux I__11567 (
            .O(N__48921),
            .I(N__48822));
    InMux I__11566 (
            .O(N__48920),
            .I(N__48822));
    Span4Mux_s3_h I__11565 (
            .O(N__48917),
            .I(N__48819));
    InMux I__11564 (
            .O(N__48916),
            .I(N__48816));
    InMux I__11563 (
            .O(N__48915),
            .I(N__48809));
    InMux I__11562 (
            .O(N__48914),
            .I(N__48809));
    InMux I__11561 (
            .O(N__48913),
            .I(N__48809));
    InMux I__11560 (
            .O(N__48912),
            .I(N__48802));
    InMux I__11559 (
            .O(N__48911),
            .I(N__48802));
    InMux I__11558 (
            .O(N__48910),
            .I(N__48802));
    InMux I__11557 (
            .O(N__48909),
            .I(N__48799));
    InMux I__11556 (
            .O(N__48908),
            .I(N__48794));
    InMux I__11555 (
            .O(N__48907),
            .I(N__48794));
    LocalMux I__11554 (
            .O(N__48904),
            .I(N__48785));
    Span4Mux_h I__11553 (
            .O(N__48901),
            .I(N__48785));
    Span4Mux_v I__11552 (
            .O(N__48894),
            .I(N__48785));
    Span4Mux_s2_h I__11551 (
            .O(N__48891),
            .I(N__48782));
    Span4Mux_s1_v I__11550 (
            .O(N__48888),
            .I(N__48779));
    Span4Mux_s1_v I__11549 (
            .O(N__48885),
            .I(N__48770));
    Span4Mux_h I__11548 (
            .O(N__48880),
            .I(N__48770));
    LocalMux I__11547 (
            .O(N__48877),
            .I(N__48770));
    Span4Mux_v I__11546 (
            .O(N__48874),
            .I(N__48770));
    LocalMux I__11545 (
            .O(N__48871),
            .I(N__48767));
    InMux I__11544 (
            .O(N__48870),
            .I(N__48764));
    Span4Mux_h I__11543 (
            .O(N__48867),
            .I(N__48750));
    LocalMux I__11542 (
            .O(N__48860),
            .I(N__48750));
    Span4Mux_v I__11541 (
            .O(N__48855),
            .I(N__48750));
    LocalMux I__11540 (
            .O(N__48846),
            .I(N__48750));
    LocalMux I__11539 (
            .O(N__48839),
            .I(N__48747));
    LocalMux I__11538 (
            .O(N__48834),
            .I(N__48742));
    LocalMux I__11537 (
            .O(N__48831),
            .I(N__48742));
    InMux I__11536 (
            .O(N__48830),
            .I(N__48739));
    LocalMux I__11535 (
            .O(N__48827),
            .I(N__48736));
    LocalMux I__11534 (
            .O(N__48822),
            .I(N__48727));
    Span4Mux_v I__11533 (
            .O(N__48819),
            .I(N__48727));
    LocalMux I__11532 (
            .O(N__48816),
            .I(N__48727));
    LocalMux I__11531 (
            .O(N__48809),
            .I(N__48727));
    LocalMux I__11530 (
            .O(N__48802),
            .I(N__48724));
    LocalMux I__11529 (
            .O(N__48799),
            .I(N__48719));
    LocalMux I__11528 (
            .O(N__48794),
            .I(N__48719));
    InMux I__11527 (
            .O(N__48793),
            .I(N__48716));
    InMux I__11526 (
            .O(N__48792),
            .I(N__48713));
    Span4Mux_h I__11525 (
            .O(N__48785),
            .I(N__48708));
    Span4Mux_h I__11524 (
            .O(N__48782),
            .I(N__48708));
    Span4Mux_h I__11523 (
            .O(N__48779),
            .I(N__48699));
    Span4Mux_h I__11522 (
            .O(N__48770),
            .I(N__48699));
    Span4Mux_s1_v I__11521 (
            .O(N__48767),
            .I(N__48699));
    LocalMux I__11520 (
            .O(N__48764),
            .I(N__48699));
    InMux I__11519 (
            .O(N__48763),
            .I(N__48690));
    InMux I__11518 (
            .O(N__48762),
            .I(N__48690));
    InMux I__11517 (
            .O(N__48761),
            .I(N__48690));
    InMux I__11516 (
            .O(N__48760),
            .I(N__48690));
    InMux I__11515 (
            .O(N__48759),
            .I(N__48687));
    Span4Mux_h I__11514 (
            .O(N__48750),
            .I(N__48674));
    Span4Mux_s3_h I__11513 (
            .O(N__48747),
            .I(N__48674));
    Span4Mux_s2_v I__11512 (
            .O(N__48742),
            .I(N__48674));
    LocalMux I__11511 (
            .O(N__48739),
            .I(N__48674));
    Span4Mux_s2_v I__11510 (
            .O(N__48736),
            .I(N__48674));
    Span4Mux_v I__11509 (
            .O(N__48727),
            .I(N__48674));
    Odrv4 I__11508 (
            .O(N__48724),
            .I(\ALU.aZ0Z_0 ));
    Odrv12 I__11507 (
            .O(N__48719),
            .I(\ALU.aZ0Z_0 ));
    LocalMux I__11506 (
            .O(N__48716),
            .I(\ALU.aZ0Z_0 ));
    LocalMux I__11505 (
            .O(N__48713),
            .I(\ALU.aZ0Z_0 ));
    Odrv4 I__11504 (
            .O(N__48708),
            .I(\ALU.aZ0Z_0 ));
    Odrv4 I__11503 (
            .O(N__48699),
            .I(\ALU.aZ0Z_0 ));
    LocalMux I__11502 (
            .O(N__48690),
            .I(\ALU.aZ0Z_0 ));
    LocalMux I__11501 (
            .O(N__48687),
            .I(\ALU.aZ0Z_0 ));
    Odrv4 I__11500 (
            .O(N__48674),
            .I(\ALU.aZ0Z_0 ));
    InMux I__11499 (
            .O(N__48655),
            .I(N__48649));
    InMux I__11498 (
            .O(N__48654),
            .I(N__48644));
    InMux I__11497 (
            .O(N__48653),
            .I(N__48641));
    InMux I__11496 (
            .O(N__48652),
            .I(N__48635));
    LocalMux I__11495 (
            .O(N__48649),
            .I(N__48632));
    InMux I__11494 (
            .O(N__48648),
            .I(N__48629));
    InMux I__11493 (
            .O(N__48647),
            .I(N__48626));
    LocalMux I__11492 (
            .O(N__48644),
            .I(N__48621));
    LocalMux I__11491 (
            .O(N__48641),
            .I(N__48621));
    InMux I__11490 (
            .O(N__48640),
            .I(N__48618));
    InMux I__11489 (
            .O(N__48639),
            .I(N__48605));
    InMux I__11488 (
            .O(N__48638),
            .I(N__48602));
    LocalMux I__11487 (
            .O(N__48635),
            .I(N__48597));
    Span4Mux_v I__11486 (
            .O(N__48632),
            .I(N__48597));
    LocalMux I__11485 (
            .O(N__48629),
            .I(N__48594));
    LocalMux I__11484 (
            .O(N__48626),
            .I(N__48587));
    Span4Mux_v I__11483 (
            .O(N__48621),
            .I(N__48587));
    LocalMux I__11482 (
            .O(N__48618),
            .I(N__48587));
    InMux I__11481 (
            .O(N__48617),
            .I(N__48582));
    InMux I__11480 (
            .O(N__48616),
            .I(N__48582));
    InMux I__11479 (
            .O(N__48615),
            .I(N__48577));
    InMux I__11478 (
            .O(N__48614),
            .I(N__48577));
    InMux I__11477 (
            .O(N__48613),
            .I(N__48572));
    InMux I__11476 (
            .O(N__48612),
            .I(N__48564));
    InMux I__11475 (
            .O(N__48611),
            .I(N__48561));
    InMux I__11474 (
            .O(N__48610),
            .I(N__48554));
    InMux I__11473 (
            .O(N__48609),
            .I(N__48554));
    InMux I__11472 (
            .O(N__48608),
            .I(N__48554));
    LocalMux I__11471 (
            .O(N__48605),
            .I(N__48550));
    LocalMux I__11470 (
            .O(N__48602),
            .I(N__48545));
    Span4Mux_v I__11469 (
            .O(N__48597),
            .I(N__48545));
    Span4Mux_h I__11468 (
            .O(N__48594),
            .I(N__48536));
    Span4Mux_v I__11467 (
            .O(N__48587),
            .I(N__48536));
    LocalMux I__11466 (
            .O(N__48582),
            .I(N__48536));
    LocalMux I__11465 (
            .O(N__48577),
            .I(N__48536));
    InMux I__11464 (
            .O(N__48576),
            .I(N__48531));
    InMux I__11463 (
            .O(N__48575),
            .I(N__48531));
    LocalMux I__11462 (
            .O(N__48572),
            .I(N__48528));
    InMux I__11461 (
            .O(N__48571),
            .I(N__48521));
    InMux I__11460 (
            .O(N__48570),
            .I(N__48521));
    InMux I__11459 (
            .O(N__48569),
            .I(N__48521));
    InMux I__11458 (
            .O(N__48568),
            .I(N__48516));
    InMux I__11457 (
            .O(N__48567),
            .I(N__48516));
    LocalMux I__11456 (
            .O(N__48564),
            .I(N__48506));
    LocalMux I__11455 (
            .O(N__48561),
            .I(N__48500));
    LocalMux I__11454 (
            .O(N__48554),
            .I(N__48500));
    InMux I__11453 (
            .O(N__48553),
            .I(N__48497));
    Span4Mux_s3_v I__11452 (
            .O(N__48550),
            .I(N__48490));
    Span4Mux_v I__11451 (
            .O(N__48545),
            .I(N__48490));
    Span4Mux_h I__11450 (
            .O(N__48536),
            .I(N__48490));
    LocalMux I__11449 (
            .O(N__48531),
            .I(N__48487));
    Span4Mux_h I__11448 (
            .O(N__48528),
            .I(N__48484));
    LocalMux I__11447 (
            .O(N__48521),
            .I(N__48479));
    LocalMux I__11446 (
            .O(N__48516),
            .I(N__48479));
    InMux I__11445 (
            .O(N__48515),
            .I(N__48474));
    InMux I__11444 (
            .O(N__48514),
            .I(N__48474));
    InMux I__11443 (
            .O(N__48513),
            .I(N__48469));
    InMux I__11442 (
            .O(N__48512),
            .I(N__48464));
    InMux I__11441 (
            .O(N__48511),
            .I(N__48464));
    InMux I__11440 (
            .O(N__48510),
            .I(N__48461));
    InMux I__11439 (
            .O(N__48509),
            .I(N__48458));
    Span4Mux_s3_v I__11438 (
            .O(N__48506),
            .I(N__48455));
    InMux I__11437 (
            .O(N__48505),
            .I(N__48452));
    Span4Mux_v I__11436 (
            .O(N__48500),
            .I(N__48443));
    LocalMux I__11435 (
            .O(N__48497),
            .I(N__48443));
    Span4Mux_h I__11434 (
            .O(N__48490),
            .I(N__48443));
    Span4Mux_s3_v I__11433 (
            .O(N__48487),
            .I(N__48443));
    Span4Mux_v I__11432 (
            .O(N__48484),
            .I(N__48436));
    Span4Mux_h I__11431 (
            .O(N__48479),
            .I(N__48436));
    LocalMux I__11430 (
            .O(N__48474),
            .I(N__48436));
    InMux I__11429 (
            .O(N__48473),
            .I(N__48431));
    InMux I__11428 (
            .O(N__48472),
            .I(N__48431));
    LocalMux I__11427 (
            .O(N__48469),
            .I(N__48426));
    LocalMux I__11426 (
            .O(N__48464),
            .I(N__48426));
    LocalMux I__11425 (
            .O(N__48461),
            .I(\ALU.a_1 ));
    LocalMux I__11424 (
            .O(N__48458),
            .I(\ALU.a_1 ));
    Odrv4 I__11423 (
            .O(N__48455),
            .I(\ALU.a_1 ));
    LocalMux I__11422 (
            .O(N__48452),
            .I(\ALU.a_1 ));
    Odrv4 I__11421 (
            .O(N__48443),
            .I(\ALU.a_1 ));
    Odrv4 I__11420 (
            .O(N__48436),
            .I(\ALU.a_1 ));
    LocalMux I__11419 (
            .O(N__48431),
            .I(\ALU.a_1 ));
    Odrv4 I__11418 (
            .O(N__48426),
            .I(\ALU.a_1 ));
    CascadeMux I__11417 (
            .O(N__48409),
            .I(N__48396));
    InMux I__11416 (
            .O(N__48408),
            .I(N__48392));
    InMux I__11415 (
            .O(N__48407),
            .I(N__48387));
    InMux I__11414 (
            .O(N__48406),
            .I(N__48384));
    InMux I__11413 (
            .O(N__48405),
            .I(N__48381));
    InMux I__11412 (
            .O(N__48404),
            .I(N__48378));
    InMux I__11411 (
            .O(N__48403),
            .I(N__48373));
    InMux I__11410 (
            .O(N__48402),
            .I(N__48373));
    InMux I__11409 (
            .O(N__48401),
            .I(N__48370));
    InMux I__11408 (
            .O(N__48400),
            .I(N__48367));
    InMux I__11407 (
            .O(N__48399),
            .I(N__48358));
    InMux I__11406 (
            .O(N__48396),
            .I(N__48355));
    InMux I__11405 (
            .O(N__48395),
            .I(N__48352));
    LocalMux I__11404 (
            .O(N__48392),
            .I(N__48348));
    InMux I__11403 (
            .O(N__48391),
            .I(N__48343));
    InMux I__11402 (
            .O(N__48390),
            .I(N__48343));
    LocalMux I__11401 (
            .O(N__48387),
            .I(N__48339));
    LocalMux I__11400 (
            .O(N__48384),
            .I(N__48336));
    LocalMux I__11399 (
            .O(N__48381),
            .I(N__48330));
    LocalMux I__11398 (
            .O(N__48378),
            .I(N__48330));
    LocalMux I__11397 (
            .O(N__48373),
            .I(N__48327));
    LocalMux I__11396 (
            .O(N__48370),
            .I(N__48324));
    LocalMux I__11395 (
            .O(N__48367),
            .I(N__48320));
    InMux I__11394 (
            .O(N__48366),
            .I(N__48315));
    InMux I__11393 (
            .O(N__48365),
            .I(N__48315));
    InMux I__11392 (
            .O(N__48364),
            .I(N__48308));
    InMux I__11391 (
            .O(N__48363),
            .I(N__48308));
    InMux I__11390 (
            .O(N__48362),
            .I(N__48308));
    InMux I__11389 (
            .O(N__48361),
            .I(N__48304));
    LocalMux I__11388 (
            .O(N__48358),
            .I(N__48301));
    LocalMux I__11387 (
            .O(N__48355),
            .I(N__48296));
    LocalMux I__11386 (
            .O(N__48352),
            .I(N__48296));
    InMux I__11385 (
            .O(N__48351),
            .I(N__48293));
    Span4Mux_v I__11384 (
            .O(N__48348),
            .I(N__48285));
    LocalMux I__11383 (
            .O(N__48343),
            .I(N__48282));
    InMux I__11382 (
            .O(N__48342),
            .I(N__48279));
    Span4Mux_s3_v I__11381 (
            .O(N__48339),
            .I(N__48274));
    Span4Mux_s3_v I__11380 (
            .O(N__48336),
            .I(N__48274));
    InMux I__11379 (
            .O(N__48335),
            .I(N__48271));
    Span4Mux_s3_v I__11378 (
            .O(N__48330),
            .I(N__48264));
    Span4Mux_s3_v I__11377 (
            .O(N__48327),
            .I(N__48264));
    Span4Mux_v I__11376 (
            .O(N__48324),
            .I(N__48264));
    InMux I__11375 (
            .O(N__48323),
            .I(N__48261));
    Span4Mux_v I__11374 (
            .O(N__48320),
            .I(N__48258));
    LocalMux I__11373 (
            .O(N__48315),
            .I(N__48253));
    LocalMux I__11372 (
            .O(N__48308),
            .I(N__48253));
    InMux I__11371 (
            .O(N__48307),
            .I(N__48250));
    LocalMux I__11370 (
            .O(N__48304),
            .I(N__48247));
    Span4Mux_s3_v I__11369 (
            .O(N__48301),
            .I(N__48242));
    Span4Mux_v I__11368 (
            .O(N__48296),
            .I(N__48242));
    LocalMux I__11367 (
            .O(N__48293),
            .I(N__48239));
    CascadeMux I__11366 (
            .O(N__48292),
            .I(N__48236));
    InMux I__11365 (
            .O(N__48291),
            .I(N__48230));
    InMux I__11364 (
            .O(N__48290),
            .I(N__48230));
    InMux I__11363 (
            .O(N__48289),
            .I(N__48225));
    InMux I__11362 (
            .O(N__48288),
            .I(N__48225));
    Span4Mux_h I__11361 (
            .O(N__48285),
            .I(N__48222));
    Span4Mux_v I__11360 (
            .O(N__48282),
            .I(N__48217));
    LocalMux I__11359 (
            .O(N__48279),
            .I(N__48217));
    Sp12to4 I__11358 (
            .O(N__48274),
            .I(N__48206));
    LocalMux I__11357 (
            .O(N__48271),
            .I(N__48206));
    Sp12to4 I__11356 (
            .O(N__48264),
            .I(N__48206));
    LocalMux I__11355 (
            .O(N__48261),
            .I(N__48206));
    Sp12to4 I__11354 (
            .O(N__48258),
            .I(N__48206));
    Span4Mux_v I__11353 (
            .O(N__48253),
            .I(N__48195));
    LocalMux I__11352 (
            .O(N__48250),
            .I(N__48195));
    Span4Mux_s3_v I__11351 (
            .O(N__48247),
            .I(N__48195));
    Span4Mux_h I__11350 (
            .O(N__48242),
            .I(N__48195));
    Span4Mux_s3_v I__11349 (
            .O(N__48239),
            .I(N__48195));
    InMux I__11348 (
            .O(N__48236),
            .I(N__48190));
    InMux I__11347 (
            .O(N__48235),
            .I(N__48190));
    LocalMux I__11346 (
            .O(N__48230),
            .I(N__48185));
    LocalMux I__11345 (
            .O(N__48225),
            .I(N__48185));
    Span4Mux_v I__11344 (
            .O(N__48222),
            .I(N__48180));
    Span4Mux_h I__11343 (
            .O(N__48217),
            .I(N__48180));
    Odrv12 I__11342 (
            .O(N__48206),
            .I(\ALU.a_2 ));
    Odrv4 I__11341 (
            .O(N__48195),
            .I(\ALU.a_2 ));
    LocalMux I__11340 (
            .O(N__48190),
            .I(\ALU.a_2 ));
    Odrv4 I__11339 (
            .O(N__48185),
            .I(\ALU.a_2 ));
    Odrv4 I__11338 (
            .O(N__48180),
            .I(\ALU.a_2 ));
    CascadeMux I__11337 (
            .O(N__48169),
            .I(\ALU.rshift_3_ns_1_0_cascade_ ));
    InMux I__11336 (
            .O(N__48166),
            .I(N__48163));
    LocalMux I__11335 (
            .O(N__48163),
            .I(N__48160));
    Span4Mux_s3_v I__11334 (
            .O(N__48160),
            .I(N__48157));
    Span4Mux_h I__11333 (
            .O(N__48157),
            .I(N__48154));
    Odrv4 I__11332 (
            .O(N__48154),
            .I(\ALU.r4_RNII2A0LZ0Z_2 ));
    InMux I__11331 (
            .O(N__48151),
            .I(N__48147));
    CascadeMux I__11330 (
            .O(N__48150),
            .I(N__48144));
    LocalMux I__11329 (
            .O(N__48147),
            .I(N__48141));
    InMux I__11328 (
            .O(N__48144),
            .I(N__48138));
    Span4Mux_h I__11327 (
            .O(N__48141),
            .I(N__48131));
    LocalMux I__11326 (
            .O(N__48138),
            .I(N__48131));
    InMux I__11325 (
            .O(N__48137),
            .I(N__48128));
    InMux I__11324 (
            .O(N__48136),
            .I(N__48125));
    Odrv4 I__11323 (
            .O(N__48131),
            .I(\ALU.lshift_5 ));
    LocalMux I__11322 (
            .O(N__48128),
            .I(\ALU.lshift_5 ));
    LocalMux I__11321 (
            .O(N__48125),
            .I(\ALU.lshift_5 ));
    CascadeMux I__11320 (
            .O(N__48118),
            .I(N__48115));
    InMux I__11319 (
            .O(N__48115),
            .I(N__48112));
    LocalMux I__11318 (
            .O(N__48112),
            .I(N__48109));
    Span4Mux_h I__11317 (
            .O(N__48109),
            .I(N__48106));
    Span4Mux_v I__11316 (
            .O(N__48106),
            .I(N__48103));
    Odrv4 I__11315 (
            .O(N__48103),
            .I(\ALU.r0_12_prm_8_5_s0_c_RNOZ0 ));
    CascadeMux I__11314 (
            .O(N__48100),
            .I(N__48097));
    InMux I__11313 (
            .O(N__48097),
            .I(N__48094));
    LocalMux I__11312 (
            .O(N__48094),
            .I(N__48091));
    Span4Mux_v I__11311 (
            .O(N__48091),
            .I(N__48088));
    Span4Mux_h I__11310 (
            .O(N__48088),
            .I(N__48085));
    Span4Mux_h I__11309 (
            .O(N__48085),
            .I(N__48082));
    Odrv4 I__11308 (
            .O(N__48082),
            .I(\ALU.r4_RNI0C236Z0Z_9 ));
    InMux I__11307 (
            .O(N__48079),
            .I(N__48073));
    InMux I__11306 (
            .O(N__48078),
            .I(N__48070));
    InMux I__11305 (
            .O(N__48077),
            .I(N__48065));
    InMux I__11304 (
            .O(N__48076),
            .I(N__48065));
    LocalMux I__11303 (
            .O(N__48073),
            .I(N__48062));
    LocalMux I__11302 (
            .O(N__48070),
            .I(N__48058));
    LocalMux I__11301 (
            .O(N__48065),
            .I(N__48055));
    Span4Mux_h I__11300 (
            .O(N__48062),
            .I(N__48052));
    CascadeMux I__11299 (
            .O(N__48061),
            .I(N__48049));
    Span4Mux_v I__11298 (
            .O(N__48058),
            .I(N__48046));
    Span4Mux_v I__11297 (
            .O(N__48055),
            .I(N__48043));
    Span4Mux_h I__11296 (
            .O(N__48052),
            .I(N__48040));
    InMux I__11295 (
            .O(N__48049),
            .I(N__48037));
    Span4Mux_h I__11294 (
            .O(N__48046),
            .I(N__48034));
    Span4Mux_h I__11293 (
            .O(N__48043),
            .I(N__48031));
    Span4Mux_h I__11292 (
            .O(N__48040),
            .I(N__48026));
    LocalMux I__11291 (
            .O(N__48037),
            .I(N__48026));
    Span4Mux_h I__11290 (
            .O(N__48034),
            .I(N__48021));
    Span4Mux_h I__11289 (
            .O(N__48031),
            .I(N__48021));
    Span4Mux_v I__11288 (
            .O(N__48026),
            .I(N__48018));
    Span4Mux_v I__11287 (
            .O(N__48021),
            .I(N__48015));
    Span4Mux_s2_h I__11286 (
            .O(N__48018),
            .I(N__48012));
    Span4Mux_h I__11285 (
            .O(N__48015),
            .I(N__48009));
    Odrv4 I__11284 (
            .O(N__48012),
            .I(\ALU.a7_b_7 ));
    Odrv4 I__11283 (
            .O(N__48009),
            .I(\ALU.a7_b_7 ));
    CascadeMux I__11282 (
            .O(N__48004),
            .I(N__48001));
    InMux I__11281 (
            .O(N__48001),
            .I(N__47998));
    LocalMux I__11280 (
            .O(N__47998),
            .I(N__47995));
    Span4Mux_h I__11279 (
            .O(N__47995),
            .I(N__47992));
    Span4Mux_v I__11278 (
            .O(N__47992),
            .I(N__47989));
    Odrv4 I__11277 (
            .O(N__47989),
            .I(\ALU.r0_12_prm_7_7_s0_c_RNOZ0 ));
    InMux I__11276 (
            .O(N__47986),
            .I(N__47983));
    LocalMux I__11275 (
            .O(N__47983),
            .I(\ALU.r0_12_prm_8_14_s1_c_RNOZ0 ));
    InMux I__11274 (
            .O(N__47980),
            .I(N__47977));
    LocalMux I__11273 (
            .O(N__47977),
            .I(N__47973));
    CascadeMux I__11272 (
            .O(N__47976),
            .I(N__47970));
    Span4Mux_h I__11271 (
            .O(N__47973),
            .I(N__47966));
    InMux I__11270 (
            .O(N__47970),
            .I(N__47963));
    InMux I__11269 (
            .O(N__47969),
            .I(N__47960));
    Span4Mux_h I__11268 (
            .O(N__47966),
            .I(N__47956));
    LocalMux I__11267 (
            .O(N__47963),
            .I(N__47953));
    LocalMux I__11266 (
            .O(N__47960),
            .I(N__47950));
    InMux I__11265 (
            .O(N__47959),
            .I(N__47947));
    Odrv4 I__11264 (
            .O(N__47956),
            .I(\ALU.lshift_14 ));
    Odrv4 I__11263 (
            .O(N__47953),
            .I(\ALU.lshift_14 ));
    Odrv4 I__11262 (
            .O(N__47950),
            .I(\ALU.lshift_14 ));
    LocalMux I__11261 (
            .O(N__47947),
            .I(\ALU.lshift_14 ));
    InMux I__11260 (
            .O(N__47938),
            .I(N__47935));
    LocalMux I__11259 (
            .O(N__47935),
            .I(N__47932));
    Odrv4 I__11258 (
            .O(N__47932),
            .I(\ALU.r0_12_prm_7_14_s1_c_RNOZ0 ));
    CascadeMux I__11257 (
            .O(N__47929),
            .I(N__47925));
    InMux I__11256 (
            .O(N__47928),
            .I(N__47922));
    InMux I__11255 (
            .O(N__47925),
            .I(N__47919));
    LocalMux I__11254 (
            .O(N__47922),
            .I(N__47916));
    LocalMux I__11253 (
            .O(N__47919),
            .I(N__47913));
    Odrv12 I__11252 (
            .O(N__47916),
            .I(\ALU.r2_RNINPPC9_0Z0Z_14 ));
    Odrv4 I__11251 (
            .O(N__47913),
            .I(\ALU.r2_RNINPPC9_0Z0Z_14 ));
    InMux I__11250 (
            .O(N__47908),
            .I(N__47905));
    LocalMux I__11249 (
            .O(N__47905),
            .I(N__47902));
    Span4Mux_h I__11248 (
            .O(N__47902),
            .I(N__47899));
    Odrv4 I__11247 (
            .O(N__47899),
            .I(\ALU.r0_12_prm_6_14_s1_c_RNOZ0 ));
    CascadeMux I__11246 (
            .O(N__47896),
            .I(N__47892));
    InMux I__11245 (
            .O(N__47895),
            .I(N__47889));
    InMux I__11244 (
            .O(N__47892),
            .I(N__47886));
    LocalMux I__11243 (
            .O(N__47889),
            .I(N__47883));
    LocalMux I__11242 (
            .O(N__47886),
            .I(N__47880));
    Span4Mux_h I__11241 (
            .O(N__47883),
            .I(N__47875));
    Span4Mux_h I__11240 (
            .O(N__47880),
            .I(N__47875));
    Odrv4 I__11239 (
            .O(N__47875),
            .I(\ALU.un14_log_0_i_14 ));
    InMux I__11238 (
            .O(N__47872),
            .I(N__47869));
    LocalMux I__11237 (
            .O(N__47869),
            .I(\ALU.r0_12_prm_5_14_s1_c_RNOZ0 ));
    CascadeMux I__11236 (
            .O(N__47866),
            .I(N__47863));
    InMux I__11235 (
            .O(N__47863),
            .I(N__47860));
    LocalMux I__11234 (
            .O(N__47860),
            .I(N__47856));
    CascadeMux I__11233 (
            .O(N__47859),
            .I(N__47853));
    Span4Mux_h I__11232 (
            .O(N__47856),
            .I(N__47850));
    InMux I__11231 (
            .O(N__47853),
            .I(N__47847));
    Odrv4 I__11230 (
            .O(N__47850),
            .I(\ALU.r2_RNINPPC9_1Z0Z_14 ));
    LocalMux I__11229 (
            .O(N__47847),
            .I(\ALU.r2_RNINPPC9_1Z0Z_14 ));
    InMux I__11228 (
            .O(N__47842),
            .I(N__47839));
    LocalMux I__11227 (
            .O(N__47839),
            .I(N__47836));
    Odrv4 I__11226 (
            .O(N__47836),
            .I(\ALU.r0_12_prm_4_14_s1_c_RNOZ0 ));
    CascadeMux I__11225 (
            .O(N__47833),
            .I(N__47830));
    InMux I__11224 (
            .O(N__47830),
            .I(N__47827));
    LocalMux I__11223 (
            .O(N__47827),
            .I(N__47824));
    Span4Mux_h I__11222 (
            .O(N__47824),
            .I(N__47820));
    InMux I__11221 (
            .O(N__47823),
            .I(N__47817));
    Span4Mux_h I__11220 (
            .O(N__47820),
            .I(N__47814));
    LocalMux I__11219 (
            .O(N__47817),
            .I(\ALU.a_i_14 ));
    Odrv4 I__11218 (
            .O(N__47814),
            .I(\ALU.a_i_14 ));
    CEMux I__11217 (
            .O(N__47809),
            .I(N__47806));
    LocalMux I__11216 (
            .O(N__47806),
            .I(N__47803));
    Span4Mux_v I__11215 (
            .O(N__47803),
            .I(N__47799));
    CEMux I__11214 (
            .O(N__47802),
            .I(N__47796));
    Span4Mux_h I__11213 (
            .O(N__47799),
            .I(N__47791));
    LocalMux I__11212 (
            .O(N__47796),
            .I(N__47791));
    Span4Mux_v I__11211 (
            .O(N__47791),
            .I(N__47788));
    Span4Mux_h I__11210 (
            .O(N__47788),
            .I(N__47784));
    CEMux I__11209 (
            .O(N__47787),
            .I(N__47781));
    Span4Mux_h I__11208 (
            .O(N__47784),
            .I(N__47778));
    LocalMux I__11207 (
            .O(N__47781),
            .I(N__47775));
    Span4Mux_h I__11206 (
            .O(N__47778),
            .I(N__47772));
    Sp12to4 I__11205 (
            .O(N__47775),
            .I(N__47769));
    Odrv4 I__11204 (
            .O(N__47772),
            .I(\ALU.un1_yindexZ0Z_4 ));
    Odrv12 I__11203 (
            .O(N__47769),
            .I(\ALU.un1_yindexZ0Z_4 ));
    CEMux I__11202 (
            .O(N__47764),
            .I(N__47759));
    CEMux I__11201 (
            .O(N__47763),
            .I(N__47756));
    CEMux I__11200 (
            .O(N__47762),
            .I(N__47752));
    LocalMux I__11199 (
            .O(N__47759),
            .I(N__47749));
    LocalMux I__11198 (
            .O(N__47756),
            .I(N__47746));
    CEMux I__11197 (
            .O(N__47755),
            .I(N__47743));
    LocalMux I__11196 (
            .O(N__47752),
            .I(N__47736));
    Span4Mux_v I__11195 (
            .O(N__47749),
            .I(N__47736));
    Span4Mux_v I__11194 (
            .O(N__47746),
            .I(N__47736));
    LocalMux I__11193 (
            .O(N__47743),
            .I(N__47733));
    Span4Mux_h I__11192 (
            .O(N__47736),
            .I(N__47730));
    Sp12to4 I__11191 (
            .O(N__47733),
            .I(N__47727));
    Sp12to4 I__11190 (
            .O(N__47730),
            .I(N__47724));
    Span12Mux_s5_h I__11189 (
            .O(N__47727),
            .I(N__47719));
    Span12Mux_v I__11188 (
            .O(N__47724),
            .I(N__47719));
    Odrv12 I__11187 (
            .O(N__47719),
            .I(\ALU.un1_yindexZ0Z_5 ));
    CEMux I__11186 (
            .O(N__47716),
            .I(N__47713));
    LocalMux I__11185 (
            .O(N__47713),
            .I(N__47709));
    CEMux I__11184 (
            .O(N__47712),
            .I(N__47703));
    IoSpan4Mux I__11183 (
            .O(N__47709),
            .I(N__47700));
    CEMux I__11182 (
            .O(N__47708),
            .I(N__47697));
    CEMux I__11181 (
            .O(N__47707),
            .I(N__47694));
    CEMux I__11180 (
            .O(N__47706),
            .I(N__47691));
    LocalMux I__11179 (
            .O(N__47703),
            .I(N__47687));
    Span4Mux_s1_h I__11178 (
            .O(N__47700),
            .I(N__47681));
    LocalMux I__11177 (
            .O(N__47697),
            .I(N__47681));
    LocalMux I__11176 (
            .O(N__47694),
            .I(N__47678));
    LocalMux I__11175 (
            .O(N__47691),
            .I(N__47675));
    CEMux I__11174 (
            .O(N__47690),
            .I(N__47672));
    Span4Mux_s2_h I__11173 (
            .O(N__47687),
            .I(N__47668));
    CEMux I__11172 (
            .O(N__47686),
            .I(N__47665));
    Span4Mux_h I__11171 (
            .O(N__47681),
            .I(N__47661));
    Span4Mux_s3_h I__11170 (
            .O(N__47678),
            .I(N__47656));
    Span4Mux_s3_h I__11169 (
            .O(N__47675),
            .I(N__47656));
    LocalMux I__11168 (
            .O(N__47672),
            .I(N__47653));
    CEMux I__11167 (
            .O(N__47671),
            .I(N__47650));
    Span4Mux_v I__11166 (
            .O(N__47668),
            .I(N__47645));
    LocalMux I__11165 (
            .O(N__47665),
            .I(N__47645));
    CEMux I__11164 (
            .O(N__47664),
            .I(N__47642));
    Span4Mux_h I__11163 (
            .O(N__47661),
            .I(N__47639));
    Span4Mux_h I__11162 (
            .O(N__47656),
            .I(N__47634));
    Span4Mux_h I__11161 (
            .O(N__47653),
            .I(N__47634));
    LocalMux I__11160 (
            .O(N__47650),
            .I(N__47631));
    Span4Mux_h I__11159 (
            .O(N__47645),
            .I(N__47628));
    LocalMux I__11158 (
            .O(N__47642),
            .I(N__47625));
    Span4Mux_v I__11157 (
            .O(N__47639),
            .I(N__47622));
    Span4Mux_v I__11156 (
            .O(N__47634),
            .I(N__47619));
    Span4Mux_h I__11155 (
            .O(N__47631),
            .I(N__47616));
    Span4Mux_v I__11154 (
            .O(N__47628),
            .I(N__47611));
    Span4Mux_v I__11153 (
            .O(N__47625),
            .I(N__47611));
    Sp12to4 I__11152 (
            .O(N__47622),
            .I(N__47608));
    Span4Mux_h I__11151 (
            .O(N__47619),
            .I(N__47605));
    Span4Mux_h I__11150 (
            .O(N__47616),
            .I(N__47602));
    Span4Mux_h I__11149 (
            .O(N__47611),
            .I(N__47599));
    Span12Mux_h I__11148 (
            .O(N__47608),
            .I(N__47596));
    Span4Mux_h I__11147 (
            .O(N__47605),
            .I(N__47593));
    Span4Mux_v I__11146 (
            .O(N__47602),
            .I(N__47588));
    Span4Mux_h I__11145 (
            .O(N__47599),
            .I(N__47588));
    Odrv12 I__11144 (
            .O(N__47596),
            .I(\ALU.un1_yindexZ0Z_6 ));
    Odrv4 I__11143 (
            .O(N__47593),
            .I(\ALU.un1_yindexZ0Z_6 ));
    Odrv4 I__11142 (
            .O(N__47588),
            .I(\ALU.un1_yindexZ0Z_6 ));
    CEMux I__11141 (
            .O(N__47581),
            .I(N__47578));
    LocalMux I__11140 (
            .O(N__47578),
            .I(N__47573));
    CEMux I__11139 (
            .O(N__47577),
            .I(N__47570));
    CEMux I__11138 (
            .O(N__47576),
            .I(N__47566));
    Span4Mux_h I__11137 (
            .O(N__47573),
            .I(N__47561));
    LocalMux I__11136 (
            .O(N__47570),
            .I(N__47561));
    CEMux I__11135 (
            .O(N__47569),
            .I(N__47556));
    LocalMux I__11134 (
            .O(N__47566),
            .I(N__47553));
    Span4Mux_v I__11133 (
            .O(N__47561),
            .I(N__47550));
    CEMux I__11132 (
            .O(N__47560),
            .I(N__47547));
    CEMux I__11131 (
            .O(N__47559),
            .I(N__47544));
    LocalMux I__11130 (
            .O(N__47556),
            .I(N__47540));
    Span4Mux_h I__11129 (
            .O(N__47553),
            .I(N__47537));
    Span4Mux_h I__11128 (
            .O(N__47550),
            .I(N__47534));
    LocalMux I__11127 (
            .O(N__47547),
            .I(N__47531));
    LocalMux I__11126 (
            .O(N__47544),
            .I(N__47528));
    CEMux I__11125 (
            .O(N__47543),
            .I(N__47525));
    Span4Mux_h I__11124 (
            .O(N__47540),
            .I(N__47522));
    Span4Mux_h I__11123 (
            .O(N__47537),
            .I(N__47519));
    Sp12to4 I__11122 (
            .O(N__47534),
            .I(N__47516));
    Span4Mux_h I__11121 (
            .O(N__47531),
            .I(N__47513));
    Span4Mux_h I__11120 (
            .O(N__47528),
            .I(N__47508));
    LocalMux I__11119 (
            .O(N__47525),
            .I(N__47508));
    Span4Mux_h I__11118 (
            .O(N__47522),
            .I(N__47505));
    Span4Mux_v I__11117 (
            .O(N__47519),
            .I(N__47502));
    Span12Mux_h I__11116 (
            .O(N__47516),
            .I(N__47499));
    Span4Mux_h I__11115 (
            .O(N__47513),
            .I(N__47496));
    Span4Mux_v I__11114 (
            .O(N__47508),
            .I(N__47493));
    Odrv4 I__11113 (
            .O(N__47505),
            .I(\ALU.un1_yindexZ0Z_7 ));
    Odrv4 I__11112 (
            .O(N__47502),
            .I(\ALU.un1_yindexZ0Z_7 ));
    Odrv12 I__11111 (
            .O(N__47499),
            .I(\ALU.un1_yindexZ0Z_7 ));
    Odrv4 I__11110 (
            .O(N__47496),
            .I(\ALU.un1_yindexZ0Z_7 ));
    Odrv4 I__11109 (
            .O(N__47493),
            .I(\ALU.un1_yindexZ0Z_7 ));
    InMux I__11108 (
            .O(N__47482),
            .I(N__47479));
    LocalMux I__11107 (
            .O(N__47479),
            .I(N__47467));
    InMux I__11106 (
            .O(N__47478),
            .I(N__47464));
    InMux I__11105 (
            .O(N__47477),
            .I(N__47461));
    InMux I__11104 (
            .O(N__47476),
            .I(N__47458));
    CascadeMux I__11103 (
            .O(N__47475),
            .I(N__47452));
    InMux I__11102 (
            .O(N__47474),
            .I(N__47449));
    InMux I__11101 (
            .O(N__47473),
            .I(N__47446));
    InMux I__11100 (
            .O(N__47472),
            .I(N__47443));
    InMux I__11099 (
            .O(N__47471),
            .I(N__47440));
    InMux I__11098 (
            .O(N__47470),
            .I(N__47437));
    Span4Mux_h I__11097 (
            .O(N__47467),
            .I(N__47426));
    LocalMux I__11096 (
            .O(N__47464),
            .I(N__47426));
    LocalMux I__11095 (
            .O(N__47461),
            .I(N__47426));
    LocalMux I__11094 (
            .O(N__47458),
            .I(N__47426));
    CascadeMux I__11093 (
            .O(N__47457),
            .I(N__47420));
    CascadeMux I__11092 (
            .O(N__47456),
            .I(N__47417));
    CascadeMux I__11091 (
            .O(N__47455),
            .I(N__47414));
    InMux I__11090 (
            .O(N__47452),
            .I(N__47410));
    LocalMux I__11089 (
            .O(N__47449),
            .I(N__47407));
    LocalMux I__11088 (
            .O(N__47446),
            .I(N__47398));
    LocalMux I__11087 (
            .O(N__47443),
            .I(N__47398));
    LocalMux I__11086 (
            .O(N__47440),
            .I(N__47398));
    LocalMux I__11085 (
            .O(N__47437),
            .I(N__47398));
    InMux I__11084 (
            .O(N__47436),
            .I(N__47395));
    CascadeMux I__11083 (
            .O(N__47435),
            .I(N__47391));
    Span4Mux_h I__11082 (
            .O(N__47426),
            .I(N__47388));
    InMux I__11081 (
            .O(N__47425),
            .I(N__47385));
    InMux I__11080 (
            .O(N__47424),
            .I(N__47382));
    InMux I__11079 (
            .O(N__47423),
            .I(N__47377));
    InMux I__11078 (
            .O(N__47420),
            .I(N__47377));
    InMux I__11077 (
            .O(N__47417),
            .I(N__47374));
    InMux I__11076 (
            .O(N__47414),
            .I(N__47369));
    InMux I__11075 (
            .O(N__47413),
            .I(N__47369));
    LocalMux I__11074 (
            .O(N__47410),
            .I(N__47366));
    Span4Mux_v I__11073 (
            .O(N__47407),
            .I(N__47361));
    Span4Mux_v I__11072 (
            .O(N__47398),
            .I(N__47361));
    LocalMux I__11071 (
            .O(N__47395),
            .I(N__47358));
    InMux I__11070 (
            .O(N__47394),
            .I(N__47353));
    InMux I__11069 (
            .O(N__47391),
            .I(N__47353));
    Span4Mux_h I__11068 (
            .O(N__47388),
            .I(N__47349));
    LocalMux I__11067 (
            .O(N__47385),
            .I(N__47346));
    LocalMux I__11066 (
            .O(N__47382),
            .I(N__47343));
    LocalMux I__11065 (
            .O(N__47377),
            .I(N__47335));
    LocalMux I__11064 (
            .O(N__47374),
            .I(N__47335));
    LocalMux I__11063 (
            .O(N__47369),
            .I(N__47335));
    Span4Mux_v I__11062 (
            .O(N__47366),
            .I(N__47330));
    Span4Mux_h I__11061 (
            .O(N__47361),
            .I(N__47330));
    Span4Mux_v I__11060 (
            .O(N__47358),
            .I(N__47325));
    LocalMux I__11059 (
            .O(N__47353),
            .I(N__47325));
    InMux I__11058 (
            .O(N__47352),
            .I(N__47322));
    Span4Mux_v I__11057 (
            .O(N__47349),
            .I(N__47317));
    Span4Mux_v I__11056 (
            .O(N__47346),
            .I(N__47317));
    Span4Mux_s3_v I__11055 (
            .O(N__47343),
            .I(N__47314));
    InMux I__11054 (
            .O(N__47342),
            .I(N__47311));
    Span4Mux_v I__11053 (
            .O(N__47335),
            .I(N__47308));
    Sp12to4 I__11052 (
            .O(N__47330),
            .I(N__47305));
    Span4Mux_h I__11051 (
            .O(N__47325),
            .I(N__47302));
    LocalMux I__11050 (
            .O(N__47322),
            .I(\ALU.b_9 ));
    Odrv4 I__11049 (
            .O(N__47317),
            .I(\ALU.b_9 ));
    Odrv4 I__11048 (
            .O(N__47314),
            .I(\ALU.b_9 ));
    LocalMux I__11047 (
            .O(N__47311),
            .I(\ALU.b_9 ));
    Odrv4 I__11046 (
            .O(N__47308),
            .I(\ALU.b_9 ));
    Odrv12 I__11045 (
            .O(N__47305),
            .I(\ALU.b_9 ));
    Odrv4 I__11044 (
            .O(N__47302),
            .I(\ALU.b_9 ));
    CascadeMux I__11043 (
            .O(N__47287),
            .I(N__47284));
    InMux I__11042 (
            .O(N__47284),
            .I(N__47281));
    LocalMux I__11041 (
            .O(N__47281),
            .I(N__47278));
    Span4Mux_h I__11040 (
            .O(N__47278),
            .I(N__47275));
    Span4Mux_h I__11039 (
            .O(N__47275),
            .I(N__47272));
    Odrv4 I__11038 (
            .O(N__47272),
            .I(\ALU.r4_RNISU5D9_2Z0Z_9 ));
    CascadeMux I__11037 (
            .O(N__47269),
            .I(N__47262));
    CascadeMux I__11036 (
            .O(N__47268),
            .I(N__47259));
    InMux I__11035 (
            .O(N__47267),
            .I(N__47256));
    InMux I__11034 (
            .O(N__47266),
            .I(N__47252));
    InMux I__11033 (
            .O(N__47265),
            .I(N__47249));
    InMux I__11032 (
            .O(N__47262),
            .I(N__47244));
    InMux I__11031 (
            .O(N__47259),
            .I(N__47244));
    LocalMux I__11030 (
            .O(N__47256),
            .I(N__47241));
    InMux I__11029 (
            .O(N__47255),
            .I(N__47238));
    LocalMux I__11028 (
            .O(N__47252),
            .I(N__47233));
    LocalMux I__11027 (
            .O(N__47249),
            .I(N__47233));
    LocalMux I__11026 (
            .O(N__47244),
            .I(N__47230));
    Span12Mux_h I__11025 (
            .O(N__47241),
            .I(N__47227));
    LocalMux I__11024 (
            .O(N__47238),
            .I(N__47224));
    Span12Mux_v I__11023 (
            .O(N__47233),
            .I(N__47221));
    Span4Mux_s2_v I__11022 (
            .O(N__47230),
            .I(N__47218));
    Odrv12 I__11021 (
            .O(N__47227),
            .I(\ALU.a5_b_5 ));
    Odrv4 I__11020 (
            .O(N__47224),
            .I(\ALU.a5_b_5 ));
    Odrv12 I__11019 (
            .O(N__47221),
            .I(\ALU.a5_b_5 ));
    Odrv4 I__11018 (
            .O(N__47218),
            .I(\ALU.a5_b_5 ));
    CascadeMux I__11017 (
            .O(N__47209),
            .I(N__47206));
    InMux I__11016 (
            .O(N__47206),
            .I(N__47203));
    LocalMux I__11015 (
            .O(N__47203),
            .I(N__47200));
    Odrv12 I__11014 (
            .O(N__47200),
            .I(\ALU.r0_12_prm_7_5_s1_c_RNOZ0 ));
    InMux I__11013 (
            .O(N__47197),
            .I(N__47191));
    InMux I__11012 (
            .O(N__47196),
            .I(N__47186));
    InMux I__11011 (
            .O(N__47195),
            .I(N__47186));
    InMux I__11010 (
            .O(N__47194),
            .I(N__47179));
    LocalMux I__11009 (
            .O(N__47191),
            .I(N__47176));
    LocalMux I__11008 (
            .O(N__47186),
            .I(N__47173));
    InMux I__11007 (
            .O(N__47185),
            .I(N__47166));
    InMux I__11006 (
            .O(N__47184),
            .I(N__47166));
    InMux I__11005 (
            .O(N__47183),
            .I(N__47166));
    CascadeMux I__11004 (
            .O(N__47182),
            .I(N__47163));
    LocalMux I__11003 (
            .O(N__47179),
            .I(N__47160));
    Span4Mux_v I__11002 (
            .O(N__47176),
            .I(N__47153));
    Span4Mux_h I__11001 (
            .O(N__47173),
            .I(N__47153));
    LocalMux I__11000 (
            .O(N__47166),
            .I(N__47153));
    InMux I__10999 (
            .O(N__47163),
            .I(N__47150));
    Span4Mux_h I__10998 (
            .O(N__47160),
            .I(N__47145));
    Span4Mux_v I__10997 (
            .O(N__47153),
            .I(N__47140));
    LocalMux I__10996 (
            .O(N__47150),
            .I(N__47140));
    InMux I__10995 (
            .O(N__47149),
            .I(N__47136));
    InMux I__10994 (
            .O(N__47148),
            .I(N__47133));
    Span4Mux_v I__10993 (
            .O(N__47145),
            .I(N__47128));
    Span4Mux_h I__10992 (
            .O(N__47140),
            .I(N__47128));
    CascadeMux I__10991 (
            .O(N__47139),
            .I(N__47125));
    LocalMux I__10990 (
            .O(N__47136),
            .I(N__47122));
    LocalMux I__10989 (
            .O(N__47133),
            .I(N__47119));
    Span4Mux_h I__10988 (
            .O(N__47128),
            .I(N__47116));
    InMux I__10987 (
            .O(N__47125),
            .I(N__47113));
    Span4Mux_v I__10986 (
            .O(N__47122),
            .I(N__47107));
    Span4Mux_v I__10985 (
            .O(N__47119),
            .I(N__47107));
    Span4Mux_h I__10984 (
            .O(N__47116),
            .I(N__47102));
    LocalMux I__10983 (
            .O(N__47113),
            .I(N__47102));
    InMux I__10982 (
            .O(N__47112),
            .I(N__47099));
    Span4Mux_h I__10981 (
            .O(N__47107),
            .I(N__47096));
    Span4Mux_v I__10980 (
            .O(N__47102),
            .I(N__47093));
    LocalMux I__10979 (
            .O(N__47099),
            .I(N__47090));
    Span4Mux_h I__10978 (
            .O(N__47096),
            .I(N__47087));
    IoSpan4Mux I__10977 (
            .O(N__47093),
            .I(N__47084));
    Span4Mux_v I__10976 (
            .O(N__47090),
            .I(N__47081));
    Span4Mux_h I__10975 (
            .O(N__47087),
            .I(N__47076));
    Span4Mux_s2_h I__10974 (
            .O(N__47084),
            .I(N__47076));
    Odrv4 I__10973 (
            .O(N__47081),
            .I(\ALU.b_14 ));
    Odrv4 I__10972 (
            .O(N__47076),
            .I(\ALU.b_14 ));
    CascadeMux I__10971 (
            .O(N__47071),
            .I(N__47067));
    CascadeMux I__10970 (
            .O(N__47070),
            .I(N__47063));
    InMux I__10969 (
            .O(N__47067),
            .I(N__47060));
    InMux I__10968 (
            .O(N__47066),
            .I(N__47057));
    InMux I__10967 (
            .O(N__47063),
            .I(N__47053));
    LocalMux I__10966 (
            .O(N__47060),
            .I(N__47047));
    LocalMux I__10965 (
            .O(N__47057),
            .I(N__47042));
    InMux I__10964 (
            .O(N__47056),
            .I(N__47037));
    LocalMux I__10963 (
            .O(N__47053),
            .I(N__47034));
    InMux I__10962 (
            .O(N__47052),
            .I(N__47027));
    InMux I__10961 (
            .O(N__47051),
            .I(N__47024));
    InMux I__10960 (
            .O(N__47050),
            .I(N__47021));
    Span4Mux_v I__10959 (
            .O(N__47047),
            .I(N__47018));
    InMux I__10958 (
            .O(N__47046),
            .I(N__47015));
    InMux I__10957 (
            .O(N__47045),
            .I(N__47012));
    Span4Mux_h I__10956 (
            .O(N__47042),
            .I(N__47004));
    CascadeMux I__10955 (
            .O(N__47041),
            .I(N__46998));
    InMux I__10954 (
            .O(N__47040),
            .I(N__46995));
    LocalMux I__10953 (
            .O(N__47037),
            .I(N__46992));
    Span4Mux_v I__10952 (
            .O(N__47034),
            .I(N__46989));
    InMux I__10951 (
            .O(N__47033),
            .I(N__46985));
    InMux I__10950 (
            .O(N__47032),
            .I(N__46982));
    InMux I__10949 (
            .O(N__47031),
            .I(N__46977));
    InMux I__10948 (
            .O(N__47030),
            .I(N__46977));
    LocalMux I__10947 (
            .O(N__47027),
            .I(N__46974));
    LocalMux I__10946 (
            .O(N__47024),
            .I(N__46969));
    LocalMux I__10945 (
            .O(N__47021),
            .I(N__46969));
    Span4Mux_v I__10944 (
            .O(N__47018),
            .I(N__46966));
    LocalMux I__10943 (
            .O(N__47015),
            .I(N__46963));
    LocalMux I__10942 (
            .O(N__47012),
            .I(N__46960));
    InMux I__10941 (
            .O(N__47011),
            .I(N__46956));
    InMux I__10940 (
            .O(N__47010),
            .I(N__46949));
    InMux I__10939 (
            .O(N__47009),
            .I(N__46949));
    InMux I__10938 (
            .O(N__47008),
            .I(N__46949));
    InMux I__10937 (
            .O(N__47007),
            .I(N__46946));
    Span4Mux_h I__10936 (
            .O(N__47004),
            .I(N__46943));
    InMux I__10935 (
            .O(N__47003),
            .I(N__46940));
    InMux I__10934 (
            .O(N__47002),
            .I(N__46933));
    InMux I__10933 (
            .O(N__47001),
            .I(N__46933));
    InMux I__10932 (
            .O(N__46998),
            .I(N__46933));
    LocalMux I__10931 (
            .O(N__46995),
            .I(N__46930));
    Span4Mux_h I__10930 (
            .O(N__46992),
            .I(N__46925));
    Span4Mux_v I__10929 (
            .O(N__46989),
            .I(N__46925));
    InMux I__10928 (
            .O(N__46988),
            .I(N__46922));
    LocalMux I__10927 (
            .O(N__46985),
            .I(N__46919));
    LocalMux I__10926 (
            .O(N__46982),
            .I(N__46910));
    LocalMux I__10925 (
            .O(N__46977),
            .I(N__46910));
    Span4Mux_v I__10924 (
            .O(N__46974),
            .I(N__46910));
    Span4Mux_v I__10923 (
            .O(N__46969),
            .I(N__46910));
    Span4Mux_v I__10922 (
            .O(N__46966),
            .I(N__46907));
    Span4Mux_s2_h I__10921 (
            .O(N__46963),
            .I(N__46904));
    Span4Mux_v I__10920 (
            .O(N__46960),
            .I(N__46901));
    InMux I__10919 (
            .O(N__46959),
            .I(N__46898));
    LocalMux I__10918 (
            .O(N__46956),
            .I(N__46891));
    LocalMux I__10917 (
            .O(N__46949),
            .I(N__46891));
    LocalMux I__10916 (
            .O(N__46946),
            .I(N__46891));
    Span4Mux_h I__10915 (
            .O(N__46943),
            .I(N__46886));
    LocalMux I__10914 (
            .O(N__46940),
            .I(N__46886));
    LocalMux I__10913 (
            .O(N__46933),
            .I(N__46883));
    Span4Mux_v I__10912 (
            .O(N__46930),
            .I(N__46870));
    Span4Mux_v I__10911 (
            .O(N__46925),
            .I(N__46870));
    LocalMux I__10910 (
            .O(N__46922),
            .I(N__46870));
    Span4Mux_h I__10909 (
            .O(N__46919),
            .I(N__46870));
    Span4Mux_h I__10908 (
            .O(N__46910),
            .I(N__46870));
    Span4Mux_h I__10907 (
            .O(N__46907),
            .I(N__46870));
    Span4Mux_h I__10906 (
            .O(N__46904),
            .I(N__46867));
    Odrv4 I__10905 (
            .O(N__46901),
            .I(\ALU.a_14 ));
    LocalMux I__10904 (
            .O(N__46898),
            .I(\ALU.a_14 ));
    Odrv12 I__10903 (
            .O(N__46891),
            .I(\ALU.a_14 ));
    Odrv4 I__10902 (
            .O(N__46886),
            .I(\ALU.a_14 ));
    Odrv12 I__10901 (
            .O(N__46883),
            .I(\ALU.a_14 ));
    Odrv4 I__10900 (
            .O(N__46870),
            .I(\ALU.a_14 ));
    Odrv4 I__10899 (
            .O(N__46867),
            .I(\ALU.a_14 ));
    CascadeMux I__10898 (
            .O(N__46852),
            .I(N__46849));
    InMux I__10897 (
            .O(N__46849),
            .I(N__46846));
    LocalMux I__10896 (
            .O(N__46846),
            .I(N__46843));
    Span12Mux_s3_v I__10895 (
            .O(N__46843),
            .I(N__46840));
    Odrv12 I__10894 (
            .O(N__46840),
            .I(\ALU.r0_12_prm_7_7_s1_c_RNOZ0 ));
    InMux I__10893 (
            .O(N__46837),
            .I(N__46834));
    LocalMux I__10892 (
            .O(N__46834),
            .I(N__46828));
    InMux I__10891 (
            .O(N__46833),
            .I(N__46825));
    CascadeMux I__10890 (
            .O(N__46832),
            .I(N__46819));
    InMux I__10889 (
            .O(N__46831),
            .I(N__46816));
    Span4Mux_v I__10888 (
            .O(N__46828),
            .I(N__46811));
    LocalMux I__10887 (
            .O(N__46825),
            .I(N__46811));
    InMux I__10886 (
            .O(N__46824),
            .I(N__46808));
    CascadeMux I__10885 (
            .O(N__46823),
            .I(N__46802));
    InMux I__10884 (
            .O(N__46822),
            .I(N__46799));
    InMux I__10883 (
            .O(N__46819),
            .I(N__46790));
    LocalMux I__10882 (
            .O(N__46816),
            .I(N__46782));
    Span4Mux_h I__10881 (
            .O(N__46811),
            .I(N__46782));
    LocalMux I__10880 (
            .O(N__46808),
            .I(N__46782));
    InMux I__10879 (
            .O(N__46807),
            .I(N__46772));
    InMux I__10878 (
            .O(N__46806),
            .I(N__46767));
    InMux I__10877 (
            .O(N__46805),
            .I(N__46767));
    InMux I__10876 (
            .O(N__46802),
            .I(N__46764));
    LocalMux I__10875 (
            .O(N__46799),
            .I(N__46761));
    InMux I__10874 (
            .O(N__46798),
            .I(N__46758));
    InMux I__10873 (
            .O(N__46797),
            .I(N__46755));
    InMux I__10872 (
            .O(N__46796),
            .I(N__46751));
    InMux I__10871 (
            .O(N__46795),
            .I(N__46737));
    InMux I__10870 (
            .O(N__46794),
            .I(N__46737));
    InMux I__10869 (
            .O(N__46793),
            .I(N__46737));
    LocalMux I__10868 (
            .O(N__46790),
            .I(N__46734));
    InMux I__10867 (
            .O(N__46789),
            .I(N__46731));
    Span4Mux_h I__10866 (
            .O(N__46782),
            .I(N__46728));
    InMux I__10865 (
            .O(N__46781),
            .I(N__46723));
    InMux I__10864 (
            .O(N__46780),
            .I(N__46723));
    InMux I__10863 (
            .O(N__46779),
            .I(N__46714));
    InMux I__10862 (
            .O(N__46778),
            .I(N__46714));
    InMux I__10861 (
            .O(N__46777),
            .I(N__46714));
    InMux I__10860 (
            .O(N__46776),
            .I(N__46714));
    CascadeMux I__10859 (
            .O(N__46775),
            .I(N__46711));
    LocalMux I__10858 (
            .O(N__46772),
            .I(N__46705));
    LocalMux I__10857 (
            .O(N__46767),
            .I(N__46705));
    LocalMux I__10856 (
            .O(N__46764),
            .I(N__46702));
    Span4Mux_v I__10855 (
            .O(N__46761),
            .I(N__46699));
    LocalMux I__10854 (
            .O(N__46758),
            .I(N__46694));
    LocalMux I__10853 (
            .O(N__46755),
            .I(N__46694));
    CascadeMux I__10852 (
            .O(N__46754),
            .I(N__46690));
    LocalMux I__10851 (
            .O(N__46751),
            .I(N__46687));
    InMux I__10850 (
            .O(N__46750),
            .I(N__46684));
    InMux I__10849 (
            .O(N__46749),
            .I(N__46681));
    InMux I__10848 (
            .O(N__46748),
            .I(N__46673));
    InMux I__10847 (
            .O(N__46747),
            .I(N__46673));
    InMux I__10846 (
            .O(N__46746),
            .I(N__46663));
    InMux I__10845 (
            .O(N__46745),
            .I(N__46663));
    InMux I__10844 (
            .O(N__46744),
            .I(N__46663));
    LocalMux I__10843 (
            .O(N__46737),
            .I(N__46660));
    Span4Mux_v I__10842 (
            .O(N__46734),
            .I(N__46655));
    LocalMux I__10841 (
            .O(N__46731),
            .I(N__46655));
    Span4Mux_v I__10840 (
            .O(N__46728),
            .I(N__46652));
    LocalMux I__10839 (
            .O(N__46723),
            .I(N__46647));
    LocalMux I__10838 (
            .O(N__46714),
            .I(N__46647));
    InMux I__10837 (
            .O(N__46711),
            .I(N__46644));
    InMux I__10836 (
            .O(N__46710),
            .I(N__46641));
    Span4Mux_v I__10835 (
            .O(N__46705),
            .I(N__46638));
    Span4Mux_h I__10834 (
            .O(N__46702),
            .I(N__46631));
    Span4Mux_h I__10833 (
            .O(N__46699),
            .I(N__46631));
    Span4Mux_s2_v I__10832 (
            .O(N__46694),
            .I(N__46631));
    InMux I__10831 (
            .O(N__46693),
            .I(N__46626));
    InMux I__10830 (
            .O(N__46690),
            .I(N__46626));
    Span4Mux_s1_h I__10829 (
            .O(N__46687),
            .I(N__46621));
    LocalMux I__10828 (
            .O(N__46684),
            .I(N__46621));
    LocalMux I__10827 (
            .O(N__46681),
            .I(N__46618));
    InMux I__10826 (
            .O(N__46680),
            .I(N__46615));
    InMux I__10825 (
            .O(N__46679),
            .I(N__46612));
    InMux I__10824 (
            .O(N__46678),
            .I(N__46609));
    LocalMux I__10823 (
            .O(N__46673),
            .I(N__46606));
    InMux I__10822 (
            .O(N__46672),
            .I(N__46603));
    InMux I__10821 (
            .O(N__46671),
            .I(N__46598));
    InMux I__10820 (
            .O(N__46670),
            .I(N__46598));
    LocalMux I__10819 (
            .O(N__46663),
            .I(N__46595));
    Span4Mux_s3_h I__10818 (
            .O(N__46660),
            .I(N__46586));
    Span4Mux_s3_h I__10817 (
            .O(N__46655),
            .I(N__46586));
    Span4Mux_v I__10816 (
            .O(N__46652),
            .I(N__46586));
    Span4Mux_v I__10815 (
            .O(N__46647),
            .I(N__46586));
    LocalMux I__10814 (
            .O(N__46644),
            .I(N__46575));
    LocalMux I__10813 (
            .O(N__46641),
            .I(N__46575));
    Span4Mux_h I__10812 (
            .O(N__46638),
            .I(N__46575));
    Span4Mux_h I__10811 (
            .O(N__46631),
            .I(N__46575));
    LocalMux I__10810 (
            .O(N__46626),
            .I(N__46575));
    Span4Mux_h I__10809 (
            .O(N__46621),
            .I(N__46572));
    Odrv12 I__10808 (
            .O(N__46618),
            .I(\ALU.b_1 ));
    LocalMux I__10807 (
            .O(N__46615),
            .I(\ALU.b_1 ));
    LocalMux I__10806 (
            .O(N__46612),
            .I(\ALU.b_1 ));
    LocalMux I__10805 (
            .O(N__46609),
            .I(\ALU.b_1 ));
    Odrv4 I__10804 (
            .O(N__46606),
            .I(\ALU.b_1 ));
    LocalMux I__10803 (
            .O(N__46603),
            .I(\ALU.b_1 ));
    LocalMux I__10802 (
            .O(N__46598),
            .I(\ALU.b_1 ));
    Odrv4 I__10801 (
            .O(N__46595),
            .I(\ALU.b_1 ));
    Odrv4 I__10800 (
            .O(N__46586),
            .I(\ALU.b_1 ));
    Odrv4 I__10799 (
            .O(N__46575),
            .I(\ALU.b_1 ));
    Odrv4 I__10798 (
            .O(N__46572),
            .I(\ALU.b_1 ));
    CascadeMux I__10797 (
            .O(N__46549),
            .I(N__46546));
    InMux I__10796 (
            .O(N__46546),
            .I(N__46543));
    LocalMux I__10795 (
            .O(N__46543),
            .I(N__46540));
    Span4Mux_h I__10794 (
            .O(N__46540),
            .I(N__46537));
    Odrv4 I__10793 (
            .O(N__46537),
            .I(\ALU.un14_log_0_i_1 ));
    CascadeMux I__10792 (
            .O(N__46534),
            .I(N__46531));
    InMux I__10791 (
            .O(N__46531),
            .I(N__46528));
    LocalMux I__10790 (
            .O(N__46528),
            .I(\ALU.r0_12_prm_5_1_c_RNOZ0Z_0 ));
    InMux I__10789 (
            .O(N__46525),
            .I(N__46522));
    LocalMux I__10788 (
            .O(N__46522),
            .I(N__46519));
    Span4Mux_v I__10787 (
            .O(N__46519),
            .I(N__46516));
    Span4Mux_h I__10786 (
            .O(N__46516),
            .I(N__46513));
    Odrv4 I__10785 (
            .O(N__46513),
            .I(\ALU.rshift_14 ));
    InMux I__10784 (
            .O(N__46510),
            .I(N__46506));
    InMux I__10783 (
            .O(N__46509),
            .I(N__46503));
    LocalMux I__10782 (
            .O(N__46506),
            .I(N__46497));
    LocalMux I__10781 (
            .O(N__46503),
            .I(N__46497));
    InMux I__10780 (
            .O(N__46502),
            .I(N__46494));
    Span4Mux_v I__10779 (
            .O(N__46497),
            .I(N__46488));
    LocalMux I__10778 (
            .O(N__46494),
            .I(N__46488));
    InMux I__10777 (
            .O(N__46493),
            .I(N__46485));
    Span4Mux_v I__10776 (
            .O(N__46488),
            .I(N__46482));
    LocalMux I__10775 (
            .O(N__46485),
            .I(N__46479));
    Span4Mux_h I__10774 (
            .O(N__46482),
            .I(N__46474));
    Span4Mux_v I__10773 (
            .O(N__46479),
            .I(N__46474));
    Odrv4 I__10772 (
            .O(N__46474),
            .I(\ALU.N_622_1 ));
    InMux I__10771 (
            .O(N__46471),
            .I(N__46468));
    LocalMux I__10770 (
            .O(N__46468),
            .I(\ALU.r0_12_prm_8_1_c_RNOZ0 ));
    InMux I__10769 (
            .O(N__46465),
            .I(N__46457));
    InMux I__10768 (
            .O(N__46464),
            .I(N__46453));
    InMux I__10767 (
            .O(N__46463),
            .I(N__46450));
    InMux I__10766 (
            .O(N__46462),
            .I(N__46447));
    CascadeMux I__10765 (
            .O(N__46461),
            .I(N__46443));
    InMux I__10764 (
            .O(N__46460),
            .I(N__46440));
    LocalMux I__10763 (
            .O(N__46457),
            .I(N__46437));
    InMux I__10762 (
            .O(N__46456),
            .I(N__46434));
    LocalMux I__10761 (
            .O(N__46453),
            .I(N__46426));
    LocalMux I__10760 (
            .O(N__46450),
            .I(N__46426));
    LocalMux I__10759 (
            .O(N__46447),
            .I(N__46423));
    CascadeMux I__10758 (
            .O(N__46446),
            .I(N__46419));
    InMux I__10757 (
            .O(N__46443),
            .I(N__46416));
    LocalMux I__10756 (
            .O(N__46440),
            .I(N__46413));
    Span4Mux_h I__10755 (
            .O(N__46437),
            .I(N__46409));
    LocalMux I__10754 (
            .O(N__46434),
            .I(N__46406));
    InMux I__10753 (
            .O(N__46433),
            .I(N__46403));
    InMux I__10752 (
            .O(N__46432),
            .I(N__46400));
    CascadeMux I__10751 (
            .O(N__46431),
            .I(N__46397));
    Span4Mux_v I__10750 (
            .O(N__46426),
            .I(N__46392));
    Span4Mux_v I__10749 (
            .O(N__46423),
            .I(N__46392));
    InMux I__10748 (
            .O(N__46422),
            .I(N__46387));
    InMux I__10747 (
            .O(N__46419),
            .I(N__46387));
    LocalMux I__10746 (
            .O(N__46416),
            .I(N__46384));
    Span4Mux_v I__10745 (
            .O(N__46413),
            .I(N__46379));
    InMux I__10744 (
            .O(N__46412),
            .I(N__46376));
    Span4Mux_h I__10743 (
            .O(N__46409),
            .I(N__46372));
    Span4Mux_v I__10742 (
            .O(N__46406),
            .I(N__46367));
    LocalMux I__10741 (
            .O(N__46403),
            .I(N__46367));
    LocalMux I__10740 (
            .O(N__46400),
            .I(N__46364));
    InMux I__10739 (
            .O(N__46397),
            .I(N__46360));
    Span4Mux_h I__10738 (
            .O(N__46392),
            .I(N__46355));
    LocalMux I__10737 (
            .O(N__46387),
            .I(N__46355));
    Span4Mux_v I__10736 (
            .O(N__46384),
            .I(N__46352));
    InMux I__10735 (
            .O(N__46383),
            .I(N__46349));
    InMux I__10734 (
            .O(N__46382),
            .I(N__46345));
    Span4Mux_h I__10733 (
            .O(N__46379),
            .I(N__46340));
    LocalMux I__10732 (
            .O(N__46376),
            .I(N__46340));
    InMux I__10731 (
            .O(N__46375),
            .I(N__46337));
    Span4Mux_h I__10730 (
            .O(N__46372),
            .I(N__46327));
    Span4Mux_h I__10729 (
            .O(N__46367),
            .I(N__46327));
    Span4Mux_h I__10728 (
            .O(N__46364),
            .I(N__46327));
    InMux I__10727 (
            .O(N__46363),
            .I(N__46324));
    LocalMux I__10726 (
            .O(N__46360),
            .I(N__46321));
    Span4Mux_v I__10725 (
            .O(N__46355),
            .I(N__46318));
    Span4Mux_h I__10724 (
            .O(N__46352),
            .I(N__46312));
    LocalMux I__10723 (
            .O(N__46349),
            .I(N__46309));
    CascadeMux I__10722 (
            .O(N__46348),
            .I(N__46304));
    LocalMux I__10721 (
            .O(N__46345),
            .I(N__46301));
    Span4Mux_v I__10720 (
            .O(N__46340),
            .I(N__46298));
    LocalMux I__10719 (
            .O(N__46337),
            .I(N__46295));
    InMux I__10718 (
            .O(N__46336),
            .I(N__46292));
    InMux I__10717 (
            .O(N__46335),
            .I(N__46287));
    InMux I__10716 (
            .O(N__46334),
            .I(N__46287));
    Span4Mux_v I__10715 (
            .O(N__46327),
            .I(N__46284));
    LocalMux I__10714 (
            .O(N__46324),
            .I(N__46281));
    Span4Mux_s2_v I__10713 (
            .O(N__46321),
            .I(N__46276));
    Span4Mux_h I__10712 (
            .O(N__46318),
            .I(N__46276));
    InMux I__10711 (
            .O(N__46317),
            .I(N__46269));
    InMux I__10710 (
            .O(N__46316),
            .I(N__46269));
    InMux I__10709 (
            .O(N__46315),
            .I(N__46269));
    Span4Mux_v I__10708 (
            .O(N__46312),
            .I(N__46264));
    Span4Mux_s2_v I__10707 (
            .O(N__46309),
            .I(N__46264));
    InMux I__10706 (
            .O(N__46308),
            .I(N__46261));
    InMux I__10705 (
            .O(N__46307),
            .I(N__46256));
    InMux I__10704 (
            .O(N__46304),
            .I(N__46256));
    Span12Mux_v I__10703 (
            .O(N__46301),
            .I(N__46245));
    Sp12to4 I__10702 (
            .O(N__46298),
            .I(N__46245));
    Span12Mux_s2_v I__10701 (
            .O(N__46295),
            .I(N__46245));
    LocalMux I__10700 (
            .O(N__46292),
            .I(N__46245));
    LocalMux I__10699 (
            .O(N__46287),
            .I(N__46245));
    Odrv4 I__10698 (
            .O(N__46284),
            .I(\ALU.b_8 ));
    Odrv4 I__10697 (
            .O(N__46281),
            .I(\ALU.b_8 ));
    Odrv4 I__10696 (
            .O(N__46276),
            .I(\ALU.b_8 ));
    LocalMux I__10695 (
            .O(N__46269),
            .I(\ALU.b_8 ));
    Odrv4 I__10694 (
            .O(N__46264),
            .I(\ALU.b_8 ));
    LocalMux I__10693 (
            .O(N__46261),
            .I(\ALU.b_8 ));
    LocalMux I__10692 (
            .O(N__46256),
            .I(\ALU.b_8 ));
    Odrv12 I__10691 (
            .O(N__46245),
            .I(\ALU.b_8 ));
    CascadeMux I__10690 (
            .O(N__46228),
            .I(N__46224));
    CascadeMux I__10689 (
            .O(N__46227),
            .I(N__46221));
    InMux I__10688 (
            .O(N__46224),
            .I(N__46211));
    InMux I__10687 (
            .O(N__46221),
            .I(N__46211));
    InMux I__10686 (
            .O(N__46220),
            .I(N__46208));
    InMux I__10685 (
            .O(N__46219),
            .I(N__46205));
    InMux I__10684 (
            .O(N__46218),
            .I(N__46201));
    CascadeMux I__10683 (
            .O(N__46217),
            .I(N__46196));
    InMux I__10682 (
            .O(N__46216),
            .I(N__46193));
    LocalMux I__10681 (
            .O(N__46211),
            .I(N__46183));
    LocalMux I__10680 (
            .O(N__46208),
            .I(N__46183));
    LocalMux I__10679 (
            .O(N__46205),
            .I(N__46174));
    InMux I__10678 (
            .O(N__46204),
            .I(N__46169));
    LocalMux I__10677 (
            .O(N__46201),
            .I(N__46166));
    InMux I__10676 (
            .O(N__46200),
            .I(N__46163));
    InMux I__10675 (
            .O(N__46199),
            .I(N__46157));
    InMux I__10674 (
            .O(N__46196),
            .I(N__46154));
    LocalMux I__10673 (
            .O(N__46193),
            .I(N__46148));
    InMux I__10672 (
            .O(N__46192),
            .I(N__46143));
    InMux I__10671 (
            .O(N__46191),
            .I(N__46143));
    InMux I__10670 (
            .O(N__46190),
            .I(N__46140));
    CascadeMux I__10669 (
            .O(N__46189),
            .I(N__46136));
    InMux I__10668 (
            .O(N__46188),
            .I(N__46132));
    Span4Mux_v I__10667 (
            .O(N__46183),
            .I(N__46129));
    InMux I__10666 (
            .O(N__46182),
            .I(N__46126));
    InMux I__10665 (
            .O(N__46181),
            .I(N__46123));
    InMux I__10664 (
            .O(N__46180),
            .I(N__46120));
    InMux I__10663 (
            .O(N__46179),
            .I(N__46115));
    InMux I__10662 (
            .O(N__46178),
            .I(N__46115));
    InMux I__10661 (
            .O(N__46177),
            .I(N__46112));
    Span4Mux_v I__10660 (
            .O(N__46174),
            .I(N__46109));
    InMux I__10659 (
            .O(N__46173),
            .I(N__46104));
    InMux I__10658 (
            .O(N__46172),
            .I(N__46104));
    LocalMux I__10657 (
            .O(N__46169),
            .I(N__46100));
    Span4Mux_v I__10656 (
            .O(N__46166),
            .I(N__46097));
    LocalMux I__10655 (
            .O(N__46163),
            .I(N__46094));
    InMux I__10654 (
            .O(N__46162),
            .I(N__46091));
    InMux I__10653 (
            .O(N__46161),
            .I(N__46086));
    InMux I__10652 (
            .O(N__46160),
            .I(N__46086));
    LocalMux I__10651 (
            .O(N__46157),
            .I(N__46081));
    LocalMux I__10650 (
            .O(N__46154),
            .I(N__46081));
    InMux I__10649 (
            .O(N__46153),
            .I(N__46075));
    InMux I__10648 (
            .O(N__46152),
            .I(N__46075));
    InMux I__10647 (
            .O(N__46151),
            .I(N__46070));
    Span4Mux_h I__10646 (
            .O(N__46148),
            .I(N__46063));
    LocalMux I__10645 (
            .O(N__46143),
            .I(N__46063));
    LocalMux I__10644 (
            .O(N__46140),
            .I(N__46063));
    InMux I__10643 (
            .O(N__46139),
            .I(N__46056));
    InMux I__10642 (
            .O(N__46136),
            .I(N__46056));
    InMux I__10641 (
            .O(N__46135),
            .I(N__46056));
    LocalMux I__10640 (
            .O(N__46132),
            .I(N__46052));
    Span4Mux_h I__10639 (
            .O(N__46129),
            .I(N__46047));
    LocalMux I__10638 (
            .O(N__46126),
            .I(N__46047));
    LocalMux I__10637 (
            .O(N__46123),
            .I(N__46036));
    LocalMux I__10636 (
            .O(N__46120),
            .I(N__46036));
    LocalMux I__10635 (
            .O(N__46115),
            .I(N__46036));
    LocalMux I__10634 (
            .O(N__46112),
            .I(N__46036));
    Sp12to4 I__10633 (
            .O(N__46109),
            .I(N__46036));
    LocalMux I__10632 (
            .O(N__46104),
            .I(N__46033));
    InMux I__10631 (
            .O(N__46103),
            .I(N__46030));
    Span4Mux_s1_v I__10630 (
            .O(N__46100),
            .I(N__46027));
    Span4Mux_h I__10629 (
            .O(N__46097),
            .I(N__46016));
    Span4Mux_v I__10628 (
            .O(N__46094),
            .I(N__46016));
    LocalMux I__10627 (
            .O(N__46091),
            .I(N__46016));
    LocalMux I__10626 (
            .O(N__46086),
            .I(N__46016));
    Span4Mux_v I__10625 (
            .O(N__46081),
            .I(N__46016));
    InMux I__10624 (
            .O(N__46080),
            .I(N__46013));
    LocalMux I__10623 (
            .O(N__46075),
            .I(N__46010));
    CascadeMux I__10622 (
            .O(N__46074),
            .I(N__46005));
    CascadeMux I__10621 (
            .O(N__46073),
            .I(N__46002));
    LocalMux I__10620 (
            .O(N__46070),
            .I(N__45999));
    Span4Mux_h I__10619 (
            .O(N__46063),
            .I(N__45996));
    LocalMux I__10618 (
            .O(N__46056),
            .I(N__45993));
    InMux I__10617 (
            .O(N__46055),
            .I(N__45990));
    Span4Mux_h I__10616 (
            .O(N__46052),
            .I(N__45983));
    Span4Mux_h I__10615 (
            .O(N__46047),
            .I(N__45983));
    Span12Mux_h I__10614 (
            .O(N__46036),
            .I(N__45980));
    Span4Mux_v I__10613 (
            .O(N__46033),
            .I(N__45971));
    LocalMux I__10612 (
            .O(N__46030),
            .I(N__45971));
    Span4Mux_v I__10611 (
            .O(N__46027),
            .I(N__45971));
    Span4Mux_h I__10610 (
            .O(N__46016),
            .I(N__45971));
    LocalMux I__10609 (
            .O(N__46013),
            .I(N__45966));
    Span4Mux_h I__10608 (
            .O(N__46010),
            .I(N__45966));
    InMux I__10607 (
            .O(N__46009),
            .I(N__45957));
    InMux I__10606 (
            .O(N__46008),
            .I(N__45957));
    InMux I__10605 (
            .O(N__46005),
            .I(N__45957));
    InMux I__10604 (
            .O(N__46002),
            .I(N__45957));
    Span12Mux_s5_v I__10603 (
            .O(N__45999),
            .I(N__45954));
    Span4Mux_h I__10602 (
            .O(N__45996),
            .I(N__45947));
    Span4Mux_h I__10601 (
            .O(N__45993),
            .I(N__45947));
    LocalMux I__10600 (
            .O(N__45990),
            .I(N__45947));
    InMux I__10599 (
            .O(N__45989),
            .I(N__45944));
    InMux I__10598 (
            .O(N__45988),
            .I(N__45941));
    Odrv4 I__10597 (
            .O(N__45983),
            .I(\ALU.a_8 ));
    Odrv12 I__10596 (
            .O(N__45980),
            .I(\ALU.a_8 ));
    Odrv4 I__10595 (
            .O(N__45971),
            .I(\ALU.a_8 ));
    Odrv4 I__10594 (
            .O(N__45966),
            .I(\ALU.a_8 ));
    LocalMux I__10593 (
            .O(N__45957),
            .I(\ALU.a_8 ));
    Odrv12 I__10592 (
            .O(N__45954),
            .I(\ALU.a_8 ));
    Odrv4 I__10591 (
            .O(N__45947),
            .I(\ALU.a_8 ));
    LocalMux I__10590 (
            .O(N__45944),
            .I(\ALU.a_8 ));
    LocalMux I__10589 (
            .O(N__45941),
            .I(\ALU.a_8 ));
    CascadeMux I__10588 (
            .O(N__45922),
            .I(N__45919));
    InMux I__10587 (
            .O(N__45919),
            .I(N__45916));
    LocalMux I__10586 (
            .O(N__45916),
            .I(N__45913));
    Odrv4 I__10585 (
            .O(N__45913),
            .I(\ALU.r0_12_prm_7_8_s1_c_RNOZ0 ));
    CascadeMux I__10584 (
            .O(N__45910),
            .I(N__45907));
    InMux I__10583 (
            .O(N__45907),
            .I(N__45904));
    LocalMux I__10582 (
            .O(N__45904),
            .I(N__45901));
    Span4Mux_h I__10581 (
            .O(N__45901),
            .I(N__45898));
    Odrv4 I__10580 (
            .O(N__45898),
            .I(\ALU.r0_12_prm_7_9_s0_c_RNOZ0 ));
    CEMux I__10579 (
            .O(N__45895),
            .I(N__45892));
    LocalMux I__10578 (
            .O(N__45892),
            .I(N__45889));
    Span4Mux_v I__10577 (
            .O(N__45889),
            .I(N__45885));
    CEMux I__10576 (
            .O(N__45888),
            .I(N__45882));
    Span4Mux_h I__10575 (
            .O(N__45885),
            .I(N__45879));
    LocalMux I__10574 (
            .O(N__45882),
            .I(N__45876));
    Span4Mux_h I__10573 (
            .O(N__45879),
            .I(N__45873));
    Span4Mux_v I__10572 (
            .O(N__45876),
            .I(N__45870));
    Span4Mux_h I__10571 (
            .O(N__45873),
            .I(N__45867));
    Span4Mux_h I__10570 (
            .O(N__45870),
            .I(N__45864));
    Span4Mux_h I__10569 (
            .O(N__45867),
            .I(N__45861));
    Span4Mux_h I__10568 (
            .O(N__45864),
            .I(N__45858));
    Odrv4 I__10567 (
            .O(N__45861),
            .I(\ALU.un1_yindexZ0Z_1 ));
    Odrv4 I__10566 (
            .O(N__45858),
            .I(\ALU.un1_yindexZ0Z_1 ));
    CEMux I__10565 (
            .O(N__45853),
            .I(N__45850));
    LocalMux I__10564 (
            .O(N__45850),
            .I(N__45847));
    Span4Mux_h I__10563 (
            .O(N__45847),
            .I(N__45843));
    CEMux I__10562 (
            .O(N__45846),
            .I(N__45839));
    Span4Mux_v I__10561 (
            .O(N__45843),
            .I(N__45836));
    CEMux I__10560 (
            .O(N__45842),
            .I(N__45833));
    LocalMux I__10559 (
            .O(N__45839),
            .I(N__45830));
    Span4Mux_h I__10558 (
            .O(N__45836),
            .I(N__45827));
    LocalMux I__10557 (
            .O(N__45833),
            .I(N__45824));
    Span4Mux_v I__10556 (
            .O(N__45830),
            .I(N__45821));
    Span4Mux_h I__10555 (
            .O(N__45827),
            .I(N__45818));
    Span12Mux_h I__10554 (
            .O(N__45824),
            .I(N__45815));
    Span4Mux_h I__10553 (
            .O(N__45821),
            .I(N__45812));
    Odrv4 I__10552 (
            .O(N__45818),
            .I(\ALU.un1_yindexZ0Z_2 ));
    Odrv12 I__10551 (
            .O(N__45815),
            .I(\ALU.un1_yindexZ0Z_2 ));
    Odrv4 I__10550 (
            .O(N__45812),
            .I(\ALU.un1_yindexZ0Z_2 ));
    CEMux I__10549 (
            .O(N__45805),
            .I(N__45802));
    LocalMux I__10548 (
            .O(N__45802),
            .I(N__45798));
    CEMux I__10547 (
            .O(N__45801),
            .I(N__45795));
    Span4Mux_v I__10546 (
            .O(N__45798),
            .I(N__45792));
    LocalMux I__10545 (
            .O(N__45795),
            .I(N__45789));
    Span4Mux_h I__10544 (
            .O(N__45792),
            .I(N__45786));
    Span4Mux_h I__10543 (
            .O(N__45789),
            .I(N__45783));
    Span4Mux_h I__10542 (
            .O(N__45786),
            .I(N__45780));
    Span4Mux_h I__10541 (
            .O(N__45783),
            .I(N__45777));
    Span4Mux_v I__10540 (
            .O(N__45780),
            .I(N__45774));
    Span4Mux_h I__10539 (
            .O(N__45777),
            .I(N__45771));
    Odrv4 I__10538 (
            .O(N__45774),
            .I(\ALU.un1_yindexZ0Z_3 ));
    Odrv4 I__10537 (
            .O(N__45771),
            .I(\ALU.un1_yindexZ0Z_3 ));
    InMux I__10536 (
            .O(N__45766),
            .I(N__45762));
    InMux I__10535 (
            .O(N__45765),
            .I(N__45759));
    LocalMux I__10534 (
            .O(N__45762),
            .I(N__45756));
    LocalMux I__10533 (
            .O(N__45759),
            .I(N__45753));
    Span4Mux_v I__10532 (
            .O(N__45756),
            .I(N__45748));
    Span4Mux_h I__10531 (
            .O(N__45753),
            .I(N__45748));
    Span4Mux_v I__10530 (
            .O(N__45748),
            .I(N__45745));
    Odrv4 I__10529 (
            .O(N__45745),
            .I(\ALU.r4_RNI8B628_0Z0Z_5 ));
    CascadeMux I__10528 (
            .O(N__45742),
            .I(N__45739));
    InMux I__10527 (
            .O(N__45739),
            .I(N__45736));
    LocalMux I__10526 (
            .O(N__45736),
            .I(\ALU.r0_12_prm_5_5_s1_c_RNOZ0 ));
    InMux I__10525 (
            .O(N__45733),
            .I(N__45730));
    LocalMux I__10524 (
            .O(N__45730),
            .I(N__45727));
    Span4Mux_v I__10523 (
            .O(N__45727),
            .I(N__45724));
    Odrv4 I__10522 (
            .O(N__45724),
            .I(\ALU.r0_12_prm_4_5_s1_c_RNOZ0 ));
    CascadeMux I__10521 (
            .O(N__45721),
            .I(N__45718));
    InMux I__10520 (
            .O(N__45718),
            .I(N__45715));
    LocalMux I__10519 (
            .O(N__45715),
            .I(N__45711));
    InMux I__10518 (
            .O(N__45714),
            .I(N__45708));
    Span4Mux_h I__10517 (
            .O(N__45711),
            .I(N__45705));
    LocalMux I__10516 (
            .O(N__45708),
            .I(\ALU.a_i_5 ));
    Odrv4 I__10515 (
            .O(N__45705),
            .I(\ALU.a_i_5 ));
    InMux I__10514 (
            .O(N__45700),
            .I(N__45697));
    LocalMux I__10513 (
            .O(N__45697),
            .I(N__45694));
    Odrv4 I__10512 (
            .O(N__45694),
            .I(\ALU.r0_12_prm_2_5_s1_c_RNOZ0 ));
    CascadeMux I__10511 (
            .O(N__45691),
            .I(N__45688));
    InMux I__10510 (
            .O(N__45688),
            .I(N__45683));
    InMux I__10509 (
            .O(N__45687),
            .I(N__45680));
    InMux I__10508 (
            .O(N__45686),
            .I(N__45677));
    LocalMux I__10507 (
            .O(N__45683),
            .I(N__45674));
    LocalMux I__10506 (
            .O(N__45680),
            .I(N__45670));
    LocalMux I__10505 (
            .O(N__45677),
            .I(N__45667));
    Span4Mux_v I__10504 (
            .O(N__45674),
            .I(N__45664));
    InMux I__10503 (
            .O(N__45673),
            .I(N__45661));
    Span4Mux_h I__10502 (
            .O(N__45670),
            .I(N__45658));
    Span4Mux_h I__10501 (
            .O(N__45667),
            .I(N__45655));
    Sp12to4 I__10500 (
            .O(N__45664),
            .I(N__45650));
    LocalMux I__10499 (
            .O(N__45661),
            .I(N__45650));
    Odrv4 I__10498 (
            .O(N__45658),
            .I(\ALU.un2_addsub_cry_4_c_RNILPG3DZ0 ));
    Odrv4 I__10497 (
            .O(N__45655),
            .I(\ALU.un2_addsub_cry_4_c_RNILPG3DZ0 ));
    Odrv12 I__10496 (
            .O(N__45650),
            .I(\ALU.un2_addsub_cry_4_c_RNILPG3DZ0 ));
    InMux I__10495 (
            .O(N__45643),
            .I(N__45640));
    LocalMux I__10494 (
            .O(N__45640),
            .I(\ALU.r0_12_prm_1_5_s1_c_RNOZ0 ));
    CascadeMux I__10493 (
            .O(N__45637),
            .I(N__45632));
    InMux I__10492 (
            .O(N__45636),
            .I(N__45629));
    InMux I__10491 (
            .O(N__45635),
            .I(N__45626));
    InMux I__10490 (
            .O(N__45632),
            .I(N__45622));
    LocalMux I__10489 (
            .O(N__45629),
            .I(N__45619));
    LocalMux I__10488 (
            .O(N__45626),
            .I(N__45616));
    InMux I__10487 (
            .O(N__45625),
            .I(N__45613));
    LocalMux I__10486 (
            .O(N__45622),
            .I(N__45610));
    Span4Mux_h I__10485 (
            .O(N__45619),
            .I(N__45607));
    Span4Mux_h I__10484 (
            .O(N__45616),
            .I(N__45604));
    LocalMux I__10483 (
            .O(N__45613),
            .I(\ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88 ));
    Odrv12 I__10482 (
            .O(N__45610),
            .I(\ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88 ));
    Odrv4 I__10481 (
            .O(N__45607),
            .I(\ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88 ));
    Odrv4 I__10480 (
            .O(N__45604),
            .I(\ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88 ));
    InMux I__10479 (
            .O(N__45595),
            .I(\ALU.r0_12_s1_5 ));
    InMux I__10478 (
            .O(N__45592),
            .I(N__45589));
    LocalMux I__10477 (
            .O(N__45589),
            .I(N__45586));
    Span4Mux_h I__10476 (
            .O(N__45586),
            .I(N__45583));
    Odrv4 I__10475 (
            .O(N__45583),
            .I(\ALU.r0_12_s1_5_THRU_CO ));
    CascadeMux I__10474 (
            .O(N__45580),
            .I(N__45577));
    InMux I__10473 (
            .O(N__45577),
            .I(N__45574));
    LocalMux I__10472 (
            .O(N__45574),
            .I(N__45571));
    Span4Mux_h I__10471 (
            .O(N__45571),
            .I(N__45568));
    Odrv4 I__10470 (
            .O(N__45568),
            .I(\ALU.r0_12_prm_5_8_s1_c_RNOZ0 ));
    CascadeMux I__10469 (
            .O(N__45565),
            .I(N__45562));
    InMux I__10468 (
            .O(N__45562),
            .I(N__45559));
    LocalMux I__10467 (
            .O(N__45559),
            .I(N__45556));
    Span4Mux_h I__10466 (
            .O(N__45556),
            .I(N__45553));
    Span4Mux_h I__10465 (
            .O(N__45553),
            .I(N__45550));
    Span4Mux_h I__10464 (
            .O(N__45550),
            .I(N__45547));
    Odrv4 I__10463 (
            .O(N__45547),
            .I(\ALU.r0_12_prm_5_10_s0_c_RNOZ0 ));
    InMux I__10462 (
            .O(N__45544),
            .I(N__45540));
    CascadeMux I__10461 (
            .O(N__45543),
            .I(N__45537));
    LocalMux I__10460 (
            .O(N__45540),
            .I(N__45534));
    InMux I__10459 (
            .O(N__45537),
            .I(N__45531));
    Span4Mux_h I__10458 (
            .O(N__45534),
            .I(N__45528));
    LocalMux I__10457 (
            .O(N__45531),
            .I(N__45525));
    Span4Mux_h I__10456 (
            .O(N__45528),
            .I(N__45520));
    Span4Mux_v I__10455 (
            .O(N__45525),
            .I(N__45520));
    Span4Mux_v I__10454 (
            .O(N__45520),
            .I(N__45517));
    Odrv4 I__10453 (
            .O(N__45517),
            .I(\ALU.un14_log_0_i_9 ));
    CascadeMux I__10452 (
            .O(N__45514),
            .I(N__45507));
    CascadeMux I__10451 (
            .O(N__45513),
            .I(N__45501));
    InMux I__10450 (
            .O(N__45512),
            .I(N__45497));
    InMux I__10449 (
            .O(N__45511),
            .I(N__45491));
    InMux I__10448 (
            .O(N__45510),
            .I(N__45488));
    InMux I__10447 (
            .O(N__45507),
            .I(N__45485));
    InMux I__10446 (
            .O(N__45506),
            .I(N__45480));
    InMux I__10445 (
            .O(N__45505),
            .I(N__45476));
    InMux I__10444 (
            .O(N__45504),
            .I(N__45473));
    InMux I__10443 (
            .O(N__45501),
            .I(N__45470));
    InMux I__10442 (
            .O(N__45500),
            .I(N__45467));
    LocalMux I__10441 (
            .O(N__45497),
            .I(N__45464));
    CascadeMux I__10440 (
            .O(N__45496),
            .I(N__45458));
    CascadeMux I__10439 (
            .O(N__45495),
            .I(N__45455));
    InMux I__10438 (
            .O(N__45494),
            .I(N__45448));
    LocalMux I__10437 (
            .O(N__45491),
            .I(N__45445));
    LocalMux I__10436 (
            .O(N__45488),
            .I(N__45440));
    LocalMux I__10435 (
            .O(N__45485),
            .I(N__45440));
    InMux I__10434 (
            .O(N__45484),
            .I(N__45435));
    InMux I__10433 (
            .O(N__45483),
            .I(N__45435));
    LocalMux I__10432 (
            .O(N__45480),
            .I(N__45432));
    InMux I__10431 (
            .O(N__45479),
            .I(N__45429));
    LocalMux I__10430 (
            .O(N__45476),
            .I(N__45426));
    LocalMux I__10429 (
            .O(N__45473),
            .I(N__45419));
    LocalMux I__10428 (
            .O(N__45470),
            .I(N__45419));
    LocalMux I__10427 (
            .O(N__45467),
            .I(N__45419));
    Span4Mux_h I__10426 (
            .O(N__45464),
            .I(N__45415));
    InMux I__10425 (
            .O(N__45463),
            .I(N__45412));
    InMux I__10424 (
            .O(N__45462),
            .I(N__45409));
    InMux I__10423 (
            .O(N__45461),
            .I(N__45406));
    InMux I__10422 (
            .O(N__45458),
            .I(N__45401));
    InMux I__10421 (
            .O(N__45455),
            .I(N__45398));
    InMux I__10420 (
            .O(N__45454),
            .I(N__45395));
    InMux I__10419 (
            .O(N__45453),
            .I(N__45392));
    InMux I__10418 (
            .O(N__45452),
            .I(N__45388));
    CascadeMux I__10417 (
            .O(N__45451),
            .I(N__45385));
    LocalMux I__10416 (
            .O(N__45448),
            .I(N__45380));
    Span4Mux_h I__10415 (
            .O(N__45445),
            .I(N__45373));
    Span4Mux_v I__10414 (
            .O(N__45440),
            .I(N__45373));
    LocalMux I__10413 (
            .O(N__45435),
            .I(N__45373));
    Span4Mux_v I__10412 (
            .O(N__45432),
            .I(N__45370));
    LocalMux I__10411 (
            .O(N__45429),
            .I(N__45367));
    Span4Mux_v I__10410 (
            .O(N__45426),
            .I(N__45362));
    Span4Mux_s1_v I__10409 (
            .O(N__45419),
            .I(N__45362));
    CascadeMux I__10408 (
            .O(N__45418),
            .I(N__45357));
    Sp12to4 I__10407 (
            .O(N__45415),
            .I(N__45354));
    LocalMux I__10406 (
            .O(N__45412),
            .I(N__45349));
    LocalMux I__10405 (
            .O(N__45409),
            .I(N__45349));
    LocalMux I__10404 (
            .O(N__45406),
            .I(N__45346));
    InMux I__10403 (
            .O(N__45405),
            .I(N__45341));
    InMux I__10402 (
            .O(N__45404),
            .I(N__45341));
    LocalMux I__10401 (
            .O(N__45401),
            .I(N__45334));
    LocalMux I__10400 (
            .O(N__45398),
            .I(N__45334));
    LocalMux I__10399 (
            .O(N__45395),
            .I(N__45334));
    LocalMux I__10398 (
            .O(N__45392),
            .I(N__45331));
    InMux I__10397 (
            .O(N__45391),
            .I(N__45328));
    LocalMux I__10396 (
            .O(N__45388),
            .I(N__45325));
    InMux I__10395 (
            .O(N__45385),
            .I(N__45322));
    InMux I__10394 (
            .O(N__45384),
            .I(N__45317));
    InMux I__10393 (
            .O(N__45383),
            .I(N__45317));
    Span4Mux_s2_v I__10392 (
            .O(N__45380),
            .I(N__45312));
    Span4Mux_v I__10391 (
            .O(N__45373),
            .I(N__45312));
    Span4Mux_h I__10390 (
            .O(N__45370),
            .I(N__45305));
    Span4Mux_v I__10389 (
            .O(N__45367),
            .I(N__45305));
    Span4Mux_h I__10388 (
            .O(N__45362),
            .I(N__45305));
    InMux I__10387 (
            .O(N__45361),
            .I(N__45300));
    InMux I__10386 (
            .O(N__45360),
            .I(N__45300));
    InMux I__10385 (
            .O(N__45357),
            .I(N__45297));
    Span12Mux_v I__10384 (
            .O(N__45354),
            .I(N__45288));
    Span12Mux_v I__10383 (
            .O(N__45349),
            .I(N__45288));
    Span12Mux_s2_h I__10382 (
            .O(N__45346),
            .I(N__45288));
    LocalMux I__10381 (
            .O(N__45341),
            .I(N__45288));
    Span4Mux_h I__10380 (
            .O(N__45334),
            .I(N__45285));
    Odrv12 I__10379 (
            .O(N__45331),
            .I(\ALU.a_5 ));
    LocalMux I__10378 (
            .O(N__45328),
            .I(\ALU.a_5 ));
    Odrv4 I__10377 (
            .O(N__45325),
            .I(\ALU.a_5 ));
    LocalMux I__10376 (
            .O(N__45322),
            .I(\ALU.a_5 ));
    LocalMux I__10375 (
            .O(N__45317),
            .I(\ALU.a_5 ));
    Odrv4 I__10374 (
            .O(N__45312),
            .I(\ALU.a_5 ));
    Odrv4 I__10373 (
            .O(N__45305),
            .I(\ALU.a_5 ));
    LocalMux I__10372 (
            .O(N__45300),
            .I(\ALU.a_5 ));
    LocalMux I__10371 (
            .O(N__45297),
            .I(\ALU.a_5 ));
    Odrv12 I__10370 (
            .O(N__45288),
            .I(\ALU.a_5 ));
    Odrv4 I__10369 (
            .O(N__45285),
            .I(\ALU.a_5 ));
    CascadeMux I__10368 (
            .O(N__45262),
            .I(N__45254));
    InMux I__10367 (
            .O(N__45261),
            .I(N__45251));
    InMux I__10366 (
            .O(N__45260),
            .I(N__45246));
    InMux I__10365 (
            .O(N__45259),
            .I(N__45243));
    CascadeMux I__10364 (
            .O(N__45258),
            .I(N__45240));
    CascadeMux I__10363 (
            .O(N__45257),
            .I(N__45237));
    InMux I__10362 (
            .O(N__45254),
            .I(N__45234));
    LocalMux I__10361 (
            .O(N__45251),
            .I(N__45226));
    InMux I__10360 (
            .O(N__45250),
            .I(N__45223));
    CascadeMux I__10359 (
            .O(N__45249),
            .I(N__45219));
    LocalMux I__10358 (
            .O(N__45246),
            .I(N__45215));
    LocalMux I__10357 (
            .O(N__45243),
            .I(N__45212));
    InMux I__10356 (
            .O(N__45240),
            .I(N__45207));
    InMux I__10355 (
            .O(N__45237),
            .I(N__45207));
    LocalMux I__10354 (
            .O(N__45234),
            .I(N__45202));
    InMux I__10353 (
            .O(N__45233),
            .I(N__45196));
    InMux I__10352 (
            .O(N__45232),
            .I(N__45196));
    InMux I__10351 (
            .O(N__45231),
            .I(N__45191));
    CascadeMux I__10350 (
            .O(N__45230),
            .I(N__45185));
    CascadeMux I__10349 (
            .O(N__45229),
            .I(N__45182));
    Span4Mux_v I__10348 (
            .O(N__45226),
            .I(N__45176));
    LocalMux I__10347 (
            .O(N__45223),
            .I(N__45173));
    InMux I__10346 (
            .O(N__45222),
            .I(N__45170));
    InMux I__10345 (
            .O(N__45219),
            .I(N__45167));
    InMux I__10344 (
            .O(N__45218),
            .I(N__45164));
    Span4Mux_v I__10343 (
            .O(N__45215),
            .I(N__45159));
    Span4Mux_h I__10342 (
            .O(N__45212),
            .I(N__45159));
    LocalMux I__10341 (
            .O(N__45207),
            .I(N__45156));
    InMux I__10340 (
            .O(N__45206),
            .I(N__45151));
    InMux I__10339 (
            .O(N__45205),
            .I(N__45151));
    Span4Mux_v I__10338 (
            .O(N__45202),
            .I(N__45148));
    InMux I__10337 (
            .O(N__45201),
            .I(N__45145));
    LocalMux I__10336 (
            .O(N__45196),
            .I(N__45142));
    InMux I__10335 (
            .O(N__45195),
            .I(N__45137));
    InMux I__10334 (
            .O(N__45194),
            .I(N__45137));
    LocalMux I__10333 (
            .O(N__45191),
            .I(N__45134));
    InMux I__10332 (
            .O(N__45190),
            .I(N__45129));
    InMux I__10331 (
            .O(N__45189),
            .I(N__45129));
    InMux I__10330 (
            .O(N__45188),
            .I(N__45121));
    InMux I__10329 (
            .O(N__45185),
            .I(N__45121));
    InMux I__10328 (
            .O(N__45182),
            .I(N__45121));
    InMux I__10327 (
            .O(N__45181),
            .I(N__45118));
    InMux I__10326 (
            .O(N__45180),
            .I(N__45115));
    InMux I__10325 (
            .O(N__45179),
            .I(N__45112));
    Span4Mux_h I__10324 (
            .O(N__45176),
            .I(N__45107));
    Span4Mux_v I__10323 (
            .O(N__45173),
            .I(N__45107));
    LocalMux I__10322 (
            .O(N__45170),
            .I(N__45103));
    LocalMux I__10321 (
            .O(N__45167),
            .I(N__45100));
    LocalMux I__10320 (
            .O(N__45164),
            .I(N__45097));
    Span4Mux_h I__10319 (
            .O(N__45159),
            .I(N__45094));
    Span4Mux_h I__10318 (
            .O(N__45156),
            .I(N__45089));
    LocalMux I__10317 (
            .O(N__45151),
            .I(N__45089));
    Span4Mux_h I__10316 (
            .O(N__45148),
            .I(N__45086));
    LocalMux I__10315 (
            .O(N__45145),
            .I(N__45081));
    Span4Mux_s0_v I__10314 (
            .O(N__45142),
            .I(N__45081));
    LocalMux I__10313 (
            .O(N__45137),
            .I(N__45078));
    Span4Mux_h I__10312 (
            .O(N__45134),
            .I(N__45073));
    LocalMux I__10311 (
            .O(N__45129),
            .I(N__45073));
    InMux I__10310 (
            .O(N__45128),
            .I(N__45070));
    LocalMux I__10309 (
            .O(N__45121),
            .I(N__45063));
    LocalMux I__10308 (
            .O(N__45118),
            .I(N__45063));
    LocalMux I__10307 (
            .O(N__45115),
            .I(N__45063));
    LocalMux I__10306 (
            .O(N__45112),
            .I(N__45060));
    Span4Mux_h I__10305 (
            .O(N__45107),
            .I(N__45057));
    InMux I__10304 (
            .O(N__45106),
            .I(N__45054));
    Span4Mux_v I__10303 (
            .O(N__45103),
            .I(N__45047));
    Span4Mux_v I__10302 (
            .O(N__45100),
            .I(N__45047));
    Span4Mux_v I__10301 (
            .O(N__45097),
            .I(N__45047));
    Span4Mux_h I__10300 (
            .O(N__45094),
            .I(N__45042));
    Span4Mux_v I__10299 (
            .O(N__45089),
            .I(N__45042));
    Span4Mux_h I__10298 (
            .O(N__45086),
            .I(N__45035));
    Span4Mux_v I__10297 (
            .O(N__45081),
            .I(N__45035));
    Span4Mux_h I__10296 (
            .O(N__45078),
            .I(N__45035));
    Span4Mux_h I__10295 (
            .O(N__45073),
            .I(N__45028));
    LocalMux I__10294 (
            .O(N__45070),
            .I(N__45028));
    Span4Mux_s2_v I__10293 (
            .O(N__45063),
            .I(N__45028));
    Odrv12 I__10292 (
            .O(N__45060),
            .I(\ALU.b_5 ));
    Odrv4 I__10291 (
            .O(N__45057),
            .I(\ALU.b_5 ));
    LocalMux I__10290 (
            .O(N__45054),
            .I(\ALU.b_5 ));
    Odrv4 I__10289 (
            .O(N__45047),
            .I(\ALU.b_5 ));
    Odrv4 I__10288 (
            .O(N__45042),
            .I(\ALU.b_5 ));
    Odrv4 I__10287 (
            .O(N__45035),
            .I(\ALU.b_5 ));
    Odrv4 I__10286 (
            .O(N__45028),
            .I(\ALU.b_5 ));
    InMux I__10285 (
            .O(N__45013),
            .I(N__45009));
    InMux I__10284 (
            .O(N__45012),
            .I(N__45006));
    LocalMux I__10283 (
            .O(N__45009),
            .I(N__45002));
    LocalMux I__10282 (
            .O(N__45006),
            .I(N__44998));
    InMux I__10281 (
            .O(N__45005),
            .I(N__44995));
    Span4Mux_h I__10280 (
            .O(N__45002),
            .I(N__44992));
    InMux I__10279 (
            .O(N__45001),
            .I(N__44989));
    Span4Mux_h I__10278 (
            .O(N__44998),
            .I(N__44986));
    LocalMux I__10277 (
            .O(N__44995),
            .I(\ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8 ));
    Odrv4 I__10276 (
            .O(N__44992),
            .I(\ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8 ));
    LocalMux I__10275 (
            .O(N__44989),
            .I(\ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8 ));
    Odrv4 I__10274 (
            .O(N__44986),
            .I(\ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8 ));
    CascadeMux I__10273 (
            .O(N__44977),
            .I(N__44974));
    InMux I__10272 (
            .O(N__44974),
            .I(N__44971));
    LocalMux I__10271 (
            .O(N__44971),
            .I(N__44968));
    Odrv4 I__10270 (
            .O(N__44968),
            .I(\ALU.r0_12_prm_1_7_s1_c_RNOZ0 ));
    InMux I__10269 (
            .O(N__44965),
            .I(N__44962));
    LocalMux I__10268 (
            .O(N__44962),
            .I(\ALU.r0_12_prm_8_5_s1_c_RNOZ0Z_1 ));
    InMux I__10267 (
            .O(N__44959),
            .I(N__44956));
    LocalMux I__10266 (
            .O(N__44956),
            .I(\ALU.r0_12_prm_8_5_s1_c_RNOZ0 ));
    InMux I__10265 (
            .O(N__44953),
            .I(N__44950));
    LocalMux I__10264 (
            .O(N__44950),
            .I(N__44947));
    Odrv12 I__10263 (
            .O(N__44947),
            .I(\ALU.r0_12_prm_6_5_s1_c_RNOZ0 ));
    InMux I__10262 (
            .O(N__44944),
            .I(N__44941));
    LocalMux I__10261 (
            .O(N__44941),
            .I(N__44937));
    CascadeMux I__10260 (
            .O(N__44940),
            .I(N__44934));
    Span4Mux_v I__10259 (
            .O(N__44937),
            .I(N__44931));
    InMux I__10258 (
            .O(N__44934),
            .I(N__44928));
    Span4Mux_h I__10257 (
            .O(N__44931),
            .I(N__44925));
    LocalMux I__10256 (
            .O(N__44928),
            .I(N__44922));
    Odrv4 I__10255 (
            .O(N__44925),
            .I(\ALU.un14_log_0_i_5 ));
    Odrv4 I__10254 (
            .O(N__44922),
            .I(\ALU.un14_log_0_i_5 ));
    InMux I__10253 (
            .O(N__44917),
            .I(\ALU.r0_12_s1_7 ));
    InMux I__10252 (
            .O(N__44914),
            .I(N__44911));
    LocalMux I__10251 (
            .O(N__44911),
            .I(N__44908));
    Span4Mux_h I__10250 (
            .O(N__44908),
            .I(N__44905));
    Odrv4 I__10249 (
            .O(N__44905),
            .I(\ALU.r0_12_s1_7_THRU_CO ));
    InMux I__10248 (
            .O(N__44902),
            .I(N__44899));
    LocalMux I__10247 (
            .O(N__44899),
            .I(N__44896));
    Span4Mux_h I__10246 (
            .O(N__44896),
            .I(N__44893));
    Span4Mux_h I__10245 (
            .O(N__44893),
            .I(N__44890));
    Span4Mux_v I__10244 (
            .O(N__44890),
            .I(N__44885));
    InMux I__10243 (
            .O(N__44889),
            .I(N__44882));
    InMux I__10242 (
            .O(N__44888),
            .I(N__44879));
    Odrv4 I__10241 (
            .O(N__44885),
            .I(\ALU.r5_RNISMSV4Z0Z_15 ));
    LocalMux I__10240 (
            .O(N__44882),
            .I(\ALU.r5_RNISMSV4Z0Z_15 ));
    LocalMux I__10239 (
            .O(N__44879),
            .I(\ALU.r5_RNISMSV4Z0Z_15 ));
    InMux I__10238 (
            .O(N__44872),
            .I(N__44869));
    LocalMux I__10237 (
            .O(N__44869),
            .I(N__44866));
    Span4Mux_h I__10236 (
            .O(N__44866),
            .I(N__44863));
    Span4Mux_h I__10235 (
            .O(N__44863),
            .I(N__44860));
    Odrv4 I__10234 (
            .O(N__44860),
            .I(\ALU.rshift_15_ns_1_3 ));
    InMux I__10233 (
            .O(N__44857),
            .I(N__44854));
    LocalMux I__10232 (
            .O(N__44854),
            .I(N__44851));
    Span4Mux_h I__10231 (
            .O(N__44851),
            .I(N__44848));
    Span4Mux_v I__10230 (
            .O(N__44848),
            .I(N__44845));
    Span4Mux_v I__10229 (
            .O(N__44845),
            .I(N__44840));
    InMux I__10228 (
            .O(N__44844),
            .I(N__44837));
    InMux I__10227 (
            .O(N__44843),
            .I(N__44834));
    Odrv4 I__10226 (
            .O(N__44840),
            .I(\ALU.r5_RNI465TIZ0Z_13 ));
    LocalMux I__10225 (
            .O(N__44837),
            .I(\ALU.r5_RNI465TIZ0Z_13 ));
    LocalMux I__10224 (
            .O(N__44834),
            .I(\ALU.r5_RNI465TIZ0Z_13 ));
    InMux I__10223 (
            .O(N__44827),
            .I(N__44824));
    LocalMux I__10222 (
            .O(N__44824),
            .I(N__44820));
    InMux I__10221 (
            .O(N__44823),
            .I(N__44817));
    Span4Mux_v I__10220 (
            .O(N__44820),
            .I(N__44814));
    LocalMux I__10219 (
            .O(N__44817),
            .I(N__44811));
    Odrv4 I__10218 (
            .O(N__44814),
            .I(\ALU.r4_RNIF01FKZ0Z_2 ));
    Odrv4 I__10217 (
            .O(N__44811),
            .I(\ALU.r4_RNIF01FKZ0Z_2 ));
    CascadeMux I__10216 (
            .O(N__44806),
            .I(N__44802));
    InMux I__10215 (
            .O(N__44805),
            .I(N__44798));
    InMux I__10214 (
            .O(N__44802),
            .I(N__44794));
    InMux I__10213 (
            .O(N__44801),
            .I(N__44791));
    LocalMux I__10212 (
            .O(N__44798),
            .I(N__44785));
    InMux I__10211 (
            .O(N__44797),
            .I(N__44780));
    LocalMux I__10210 (
            .O(N__44794),
            .I(N__44777));
    LocalMux I__10209 (
            .O(N__44791),
            .I(N__44773));
    InMux I__10208 (
            .O(N__44790),
            .I(N__44770));
    InMux I__10207 (
            .O(N__44789),
            .I(N__44767));
    InMux I__10206 (
            .O(N__44788),
            .I(N__44760));
    Span4Mux_v I__10205 (
            .O(N__44785),
            .I(N__44757));
    InMux I__10204 (
            .O(N__44784),
            .I(N__44754));
    InMux I__10203 (
            .O(N__44783),
            .I(N__44751));
    LocalMux I__10202 (
            .O(N__44780),
            .I(N__44745));
    Span4Mux_v I__10201 (
            .O(N__44777),
            .I(N__44745));
    InMux I__10200 (
            .O(N__44776),
            .I(N__44742));
    Span4Mux_v I__10199 (
            .O(N__44773),
            .I(N__44739));
    LocalMux I__10198 (
            .O(N__44770),
            .I(N__44736));
    LocalMux I__10197 (
            .O(N__44767),
            .I(N__44733));
    InMux I__10196 (
            .O(N__44766),
            .I(N__44730));
    InMux I__10195 (
            .O(N__44765),
            .I(N__44727));
    InMux I__10194 (
            .O(N__44764),
            .I(N__44724));
    CascadeMux I__10193 (
            .O(N__44763),
            .I(N__44720));
    LocalMux I__10192 (
            .O(N__44760),
            .I(N__44712));
    Sp12to4 I__10191 (
            .O(N__44757),
            .I(N__44712));
    LocalMux I__10190 (
            .O(N__44754),
            .I(N__44712));
    LocalMux I__10189 (
            .O(N__44751),
            .I(N__44709));
    InMux I__10188 (
            .O(N__44750),
            .I(N__44706));
    Span4Mux_v I__10187 (
            .O(N__44745),
            .I(N__44701));
    LocalMux I__10186 (
            .O(N__44742),
            .I(N__44698));
    Span4Mux_h I__10185 (
            .O(N__44739),
            .I(N__44691));
    Span4Mux_s2_v I__10184 (
            .O(N__44736),
            .I(N__44691));
    Span4Mux_h I__10183 (
            .O(N__44733),
            .I(N__44691));
    LocalMux I__10182 (
            .O(N__44730),
            .I(N__44688));
    LocalMux I__10181 (
            .O(N__44727),
            .I(N__44685));
    LocalMux I__10180 (
            .O(N__44724),
            .I(N__44682));
    InMux I__10179 (
            .O(N__44723),
            .I(N__44679));
    InMux I__10178 (
            .O(N__44720),
            .I(N__44670));
    InMux I__10177 (
            .O(N__44719),
            .I(N__44670));
    Span12Mux_h I__10176 (
            .O(N__44712),
            .I(N__44667));
    Span4Mux_s3_h I__10175 (
            .O(N__44709),
            .I(N__44664));
    LocalMux I__10174 (
            .O(N__44706),
            .I(N__44661));
    InMux I__10173 (
            .O(N__44705),
            .I(N__44656));
    InMux I__10172 (
            .O(N__44704),
            .I(N__44656));
    Span4Mux_h I__10171 (
            .O(N__44701),
            .I(N__44645));
    Span4Mux_v I__10170 (
            .O(N__44698),
            .I(N__44645));
    Span4Mux_h I__10169 (
            .O(N__44691),
            .I(N__44645));
    Span4Mux_s2_h I__10168 (
            .O(N__44688),
            .I(N__44645));
    Span4Mux_s2_v I__10167 (
            .O(N__44685),
            .I(N__44645));
    Span12Mux_h I__10166 (
            .O(N__44682),
            .I(N__44640));
    LocalMux I__10165 (
            .O(N__44679),
            .I(N__44640));
    InMux I__10164 (
            .O(N__44678),
            .I(N__44631));
    InMux I__10163 (
            .O(N__44677),
            .I(N__44631));
    InMux I__10162 (
            .O(N__44676),
            .I(N__44631));
    InMux I__10161 (
            .O(N__44675),
            .I(N__44631));
    LocalMux I__10160 (
            .O(N__44670),
            .I(N__44628));
    Odrv12 I__10159 (
            .O(N__44667),
            .I(\ALU.b_7 ));
    Odrv4 I__10158 (
            .O(N__44664),
            .I(\ALU.b_7 ));
    Odrv4 I__10157 (
            .O(N__44661),
            .I(\ALU.b_7 ));
    LocalMux I__10156 (
            .O(N__44656),
            .I(\ALU.b_7 ));
    Odrv4 I__10155 (
            .O(N__44645),
            .I(\ALU.b_7 ));
    Odrv12 I__10154 (
            .O(N__44640),
            .I(\ALU.b_7 ));
    LocalMux I__10153 (
            .O(N__44631),
            .I(\ALU.b_7 ));
    Odrv12 I__10152 (
            .O(N__44628),
            .I(\ALU.b_7 ));
    CascadeMux I__10151 (
            .O(N__44611),
            .I(N__44607));
    InMux I__10150 (
            .O(N__44610),
            .I(N__44604));
    InMux I__10149 (
            .O(N__44607),
            .I(N__44597));
    LocalMux I__10148 (
            .O(N__44604),
            .I(N__44590));
    InMux I__10147 (
            .O(N__44603),
            .I(N__44585));
    InMux I__10146 (
            .O(N__44602),
            .I(N__44582));
    InMux I__10145 (
            .O(N__44601),
            .I(N__44579));
    InMux I__10144 (
            .O(N__44600),
            .I(N__44576));
    LocalMux I__10143 (
            .O(N__44597),
            .I(N__44573));
    InMux I__10142 (
            .O(N__44596),
            .I(N__44570));
    InMux I__10141 (
            .O(N__44595),
            .I(N__44567));
    InMux I__10140 (
            .O(N__44594),
            .I(N__44564));
    InMux I__10139 (
            .O(N__44593),
            .I(N__44561));
    Span4Mux_v I__10138 (
            .O(N__44590),
            .I(N__44558));
    InMux I__10137 (
            .O(N__44589),
            .I(N__44553));
    InMux I__10136 (
            .O(N__44588),
            .I(N__44553));
    LocalMux I__10135 (
            .O(N__44585),
            .I(N__44546));
    LocalMux I__10134 (
            .O(N__44582),
            .I(N__44539));
    LocalMux I__10133 (
            .O(N__44579),
            .I(N__44532));
    LocalMux I__10132 (
            .O(N__44576),
            .I(N__44532));
    Span4Mux_v I__10131 (
            .O(N__44573),
            .I(N__44526));
    LocalMux I__10130 (
            .O(N__44570),
            .I(N__44523));
    LocalMux I__10129 (
            .O(N__44567),
            .I(N__44520));
    LocalMux I__10128 (
            .O(N__44564),
            .I(N__44509));
    LocalMux I__10127 (
            .O(N__44561),
            .I(N__44509));
    Span4Mux_h I__10126 (
            .O(N__44558),
            .I(N__44509));
    LocalMux I__10125 (
            .O(N__44553),
            .I(N__44509));
    InMux I__10124 (
            .O(N__44552),
            .I(N__44506));
    InMux I__10123 (
            .O(N__44551),
            .I(N__44501));
    InMux I__10122 (
            .O(N__44550),
            .I(N__44501));
    InMux I__10121 (
            .O(N__44549),
            .I(N__44498));
    Span4Mux_h I__10120 (
            .O(N__44546),
            .I(N__44495));
    InMux I__10119 (
            .O(N__44545),
            .I(N__44490));
    InMux I__10118 (
            .O(N__44544),
            .I(N__44490));
    InMux I__10117 (
            .O(N__44543),
            .I(N__44484));
    InMux I__10116 (
            .O(N__44542),
            .I(N__44481));
    Span4Mux_v I__10115 (
            .O(N__44539),
            .I(N__44478));
    InMux I__10114 (
            .O(N__44538),
            .I(N__44473));
    InMux I__10113 (
            .O(N__44537),
            .I(N__44473));
    Span4Mux_v I__10112 (
            .O(N__44532),
            .I(N__44470));
    InMux I__10111 (
            .O(N__44531),
            .I(N__44465));
    InMux I__10110 (
            .O(N__44530),
            .I(N__44465));
    InMux I__10109 (
            .O(N__44529),
            .I(N__44462));
    Span4Mux_h I__10108 (
            .O(N__44526),
            .I(N__44455));
    Span4Mux_v I__10107 (
            .O(N__44523),
            .I(N__44455));
    Span4Mux_v I__10106 (
            .O(N__44520),
            .I(N__44455));
    InMux I__10105 (
            .O(N__44519),
            .I(N__44450));
    InMux I__10104 (
            .O(N__44518),
            .I(N__44450));
    Span4Mux_v I__10103 (
            .O(N__44509),
            .I(N__44441));
    LocalMux I__10102 (
            .O(N__44506),
            .I(N__44441));
    LocalMux I__10101 (
            .O(N__44501),
            .I(N__44436));
    LocalMux I__10100 (
            .O(N__44498),
            .I(N__44436));
    Span4Mux_h I__10099 (
            .O(N__44495),
            .I(N__44430));
    LocalMux I__10098 (
            .O(N__44490),
            .I(N__44430));
    InMux I__10097 (
            .O(N__44489),
            .I(N__44423));
    InMux I__10096 (
            .O(N__44488),
            .I(N__44423));
    InMux I__10095 (
            .O(N__44487),
            .I(N__44423));
    LocalMux I__10094 (
            .O(N__44484),
            .I(N__44406));
    LocalMux I__10093 (
            .O(N__44481),
            .I(N__44406));
    Sp12to4 I__10092 (
            .O(N__44478),
            .I(N__44406));
    LocalMux I__10091 (
            .O(N__44473),
            .I(N__44406));
    Sp12to4 I__10090 (
            .O(N__44470),
            .I(N__44406));
    LocalMux I__10089 (
            .O(N__44465),
            .I(N__44406));
    LocalMux I__10088 (
            .O(N__44462),
            .I(N__44406));
    Sp12to4 I__10087 (
            .O(N__44455),
            .I(N__44406));
    LocalMux I__10086 (
            .O(N__44450),
            .I(N__44403));
    InMux I__10085 (
            .O(N__44449),
            .I(N__44394));
    InMux I__10084 (
            .O(N__44448),
            .I(N__44394));
    InMux I__10083 (
            .O(N__44447),
            .I(N__44394));
    InMux I__10082 (
            .O(N__44446),
            .I(N__44394));
    Span4Mux_h I__10081 (
            .O(N__44441),
            .I(N__44389));
    Span4Mux_v I__10080 (
            .O(N__44436),
            .I(N__44389));
    InMux I__10079 (
            .O(N__44435),
            .I(N__44386));
    Odrv4 I__10078 (
            .O(N__44430),
            .I(\ALU.a_7 ));
    LocalMux I__10077 (
            .O(N__44423),
            .I(\ALU.a_7 ));
    Odrv12 I__10076 (
            .O(N__44406),
            .I(\ALU.a_7 ));
    Odrv12 I__10075 (
            .O(N__44403),
            .I(\ALU.a_7 ));
    LocalMux I__10074 (
            .O(N__44394),
            .I(\ALU.a_7 ));
    Odrv4 I__10073 (
            .O(N__44389),
            .I(\ALU.a_7 ));
    LocalMux I__10072 (
            .O(N__44386),
            .I(\ALU.a_7 ));
    InMux I__10071 (
            .O(N__44371),
            .I(N__44368));
    LocalMux I__10070 (
            .O(N__44368),
            .I(\ALU.r0_12_prm_6_7_s1_c_RNOZ0 ));
    InMux I__10069 (
            .O(N__44365),
            .I(N__44362));
    LocalMux I__10068 (
            .O(N__44362),
            .I(N__44356));
    InMux I__10067 (
            .O(N__44361),
            .I(N__44353));
    InMux I__10066 (
            .O(N__44360),
            .I(N__44339));
    InMux I__10065 (
            .O(N__44359),
            .I(N__44336));
    Span4Mux_h I__10064 (
            .O(N__44356),
            .I(N__44332));
    LocalMux I__10063 (
            .O(N__44353),
            .I(N__44329));
    InMux I__10062 (
            .O(N__44352),
            .I(N__44322));
    InMux I__10061 (
            .O(N__44351),
            .I(N__44322));
    InMux I__10060 (
            .O(N__44350),
            .I(N__44322));
    InMux I__10059 (
            .O(N__44349),
            .I(N__44319));
    InMux I__10058 (
            .O(N__44348),
            .I(N__44314));
    InMux I__10057 (
            .O(N__44347),
            .I(N__44314));
    InMux I__10056 (
            .O(N__44346),
            .I(N__44310));
    InMux I__10055 (
            .O(N__44345),
            .I(N__44303));
    InMux I__10054 (
            .O(N__44344),
            .I(N__44303));
    InMux I__10053 (
            .O(N__44343),
            .I(N__44300));
    InMux I__10052 (
            .O(N__44342),
            .I(N__44297));
    LocalMux I__10051 (
            .O(N__44339),
            .I(N__44294));
    LocalMux I__10050 (
            .O(N__44336),
            .I(N__44291));
    InMux I__10049 (
            .O(N__44335),
            .I(N__44288));
    Span4Mux_h I__10048 (
            .O(N__44332),
            .I(N__44283));
    Span4Mux_h I__10047 (
            .O(N__44329),
            .I(N__44283));
    LocalMux I__10046 (
            .O(N__44322),
            .I(N__44280));
    LocalMux I__10045 (
            .O(N__44319),
            .I(N__44277));
    LocalMux I__10044 (
            .O(N__44314),
            .I(N__44271));
    InMux I__10043 (
            .O(N__44313),
            .I(N__44268));
    LocalMux I__10042 (
            .O(N__44310),
            .I(N__44265));
    InMux I__10041 (
            .O(N__44309),
            .I(N__44260));
    InMux I__10040 (
            .O(N__44308),
            .I(N__44260));
    LocalMux I__10039 (
            .O(N__44303),
            .I(N__44253));
    LocalMux I__10038 (
            .O(N__44300),
            .I(N__44253));
    LocalMux I__10037 (
            .O(N__44297),
            .I(N__44253));
    Span4Mux_h I__10036 (
            .O(N__44294),
            .I(N__44241));
    Span4Mux_s3_v I__10035 (
            .O(N__44291),
            .I(N__44241));
    LocalMux I__10034 (
            .O(N__44288),
            .I(N__44241));
    Sp12to4 I__10033 (
            .O(N__44283),
            .I(N__44234));
    Span12Mux_h I__10032 (
            .O(N__44280),
            .I(N__44234));
    Span12Mux_s5_h I__10031 (
            .O(N__44277),
            .I(N__44234));
    InMux I__10030 (
            .O(N__44276),
            .I(N__44227));
    InMux I__10029 (
            .O(N__44275),
            .I(N__44227));
    InMux I__10028 (
            .O(N__44274),
            .I(N__44227));
    Span4Mux_h I__10027 (
            .O(N__44271),
            .I(N__44222));
    LocalMux I__10026 (
            .O(N__44268),
            .I(N__44222));
    Span12Mux_h I__10025 (
            .O(N__44265),
            .I(N__44215));
    LocalMux I__10024 (
            .O(N__44260),
            .I(N__44215));
    Span12Mux_s5_h I__10023 (
            .O(N__44253),
            .I(N__44215));
    InMux I__10022 (
            .O(N__44252),
            .I(N__44210));
    InMux I__10021 (
            .O(N__44251),
            .I(N__44210));
    InMux I__10020 (
            .O(N__44250),
            .I(N__44203));
    InMux I__10019 (
            .O(N__44249),
            .I(N__44203));
    InMux I__10018 (
            .O(N__44248),
            .I(N__44203));
    Odrv4 I__10017 (
            .O(N__44241),
            .I(\ALU.b_3 ));
    Odrv12 I__10016 (
            .O(N__44234),
            .I(\ALU.b_3 ));
    LocalMux I__10015 (
            .O(N__44227),
            .I(\ALU.b_3 ));
    Odrv4 I__10014 (
            .O(N__44222),
            .I(\ALU.b_3 ));
    Odrv12 I__10013 (
            .O(N__44215),
            .I(\ALU.b_3 ));
    LocalMux I__10012 (
            .O(N__44210),
            .I(\ALU.b_3 ));
    LocalMux I__10011 (
            .O(N__44203),
            .I(\ALU.b_3 ));
    CascadeMux I__10010 (
            .O(N__44188),
            .I(N__44185));
    InMux I__10009 (
            .O(N__44185),
            .I(N__44182));
    LocalMux I__10008 (
            .O(N__44182),
            .I(N__44179));
    Span4Mux_h I__10007 (
            .O(N__44179),
            .I(N__44176));
    Odrv4 I__10006 (
            .O(N__44176),
            .I(\ALU.r0_12_prm_1_5_s0_c_RNOZ0 ));
    CascadeMux I__10005 (
            .O(N__44173),
            .I(N__44170));
    InMux I__10004 (
            .O(N__44170),
            .I(N__44165));
    InMux I__10003 (
            .O(N__44169),
            .I(N__44162));
    CascadeMux I__10002 (
            .O(N__44168),
            .I(N__44159));
    LocalMux I__10001 (
            .O(N__44165),
            .I(N__44155));
    LocalMux I__10000 (
            .O(N__44162),
            .I(N__44152));
    InMux I__9999 (
            .O(N__44159),
            .I(N__44149));
    InMux I__9998 (
            .O(N__44158),
            .I(N__44146));
    Span4Mux_h I__9997 (
            .O(N__44155),
            .I(N__44141));
    Span4Mux_h I__9996 (
            .O(N__44152),
            .I(N__44141));
    LocalMux I__9995 (
            .O(N__44149),
            .I(N__44136));
    LocalMux I__9994 (
            .O(N__44146),
            .I(N__44136));
    Odrv4 I__9993 (
            .O(N__44141),
            .I(\ALU.rshift_7 ));
    Odrv12 I__9992 (
            .O(N__44136),
            .I(\ALU.rshift_7 ));
    InMux I__9991 (
            .O(N__44131),
            .I(N__44128));
    LocalMux I__9990 (
            .O(N__44128),
            .I(\ALU.r0_12_prm_8_7_s1_c_RNOZ0 ));
    CascadeMux I__9989 (
            .O(N__44125),
            .I(N__44122));
    InMux I__9988 (
            .O(N__44122),
            .I(N__44119));
    LocalMux I__9987 (
            .O(N__44119),
            .I(N__44115));
    CascadeMux I__9986 (
            .O(N__44118),
            .I(N__44112));
    Span4Mux_h I__9985 (
            .O(N__44115),
            .I(N__44108));
    InMux I__9984 (
            .O(N__44112),
            .I(N__44105));
    InMux I__9983 (
            .O(N__44111),
            .I(N__44102));
    Odrv4 I__9982 (
            .O(N__44108),
            .I(\ALU.lshift_7 ));
    LocalMux I__9981 (
            .O(N__44105),
            .I(\ALU.lshift_7 ));
    LocalMux I__9980 (
            .O(N__44102),
            .I(\ALU.lshift_7 ));
    InMux I__9979 (
            .O(N__44095),
            .I(N__44091));
    CascadeMux I__9978 (
            .O(N__44094),
            .I(N__44088));
    LocalMux I__9977 (
            .O(N__44091),
            .I(N__44085));
    InMux I__9976 (
            .O(N__44088),
            .I(N__44082));
    Span4Mux_v I__9975 (
            .O(N__44085),
            .I(N__44079));
    LocalMux I__9974 (
            .O(N__44082),
            .I(N__44076));
    Span4Mux_s1_v I__9973 (
            .O(N__44079),
            .I(N__44071));
    Span4Mux_v I__9972 (
            .O(N__44076),
            .I(N__44071));
    Odrv4 I__9971 (
            .O(N__44071),
            .I(\ALU.un14_log_0_i_7 ));
    InMux I__9970 (
            .O(N__44068),
            .I(N__44065));
    LocalMux I__9969 (
            .O(N__44065),
            .I(\ALU.r0_12_prm_5_7_s1_c_RNOZ0 ));
    CascadeMux I__9968 (
            .O(N__44062),
            .I(N__44059));
    InMux I__9967 (
            .O(N__44059),
            .I(N__44056));
    LocalMux I__9966 (
            .O(N__44056),
            .I(N__44052));
    InMux I__9965 (
            .O(N__44055),
            .I(N__44049));
    Span4Mux_v I__9964 (
            .O(N__44052),
            .I(N__44046));
    LocalMux I__9963 (
            .O(N__44049),
            .I(\ALU.r4_RNIHENK8_0Z0Z_7 ));
    Odrv4 I__9962 (
            .O(N__44046),
            .I(\ALU.r4_RNIHENK8_0Z0Z_7 ));
    InMux I__9961 (
            .O(N__44041),
            .I(N__44038));
    LocalMux I__9960 (
            .O(N__44038),
            .I(\ALU.r0_12_prm_4_7_s1_c_RNOZ0 ));
    CascadeMux I__9959 (
            .O(N__44035),
            .I(N__44032));
    InMux I__9958 (
            .O(N__44032),
            .I(N__44029));
    LocalMux I__9957 (
            .O(N__44029),
            .I(N__44025));
    InMux I__9956 (
            .O(N__44028),
            .I(N__44022));
    Span4Mux_h I__9955 (
            .O(N__44025),
            .I(N__44019));
    LocalMux I__9954 (
            .O(N__44022),
            .I(\ALU.a_i_7 ));
    Odrv4 I__9953 (
            .O(N__44019),
            .I(\ALU.a_i_7 ));
    InMux I__9952 (
            .O(N__44014),
            .I(N__44010));
    InMux I__9951 (
            .O(N__44013),
            .I(N__44005));
    LocalMux I__9950 (
            .O(N__44010),
            .I(N__44002));
    InMux I__9949 (
            .O(N__44009),
            .I(N__43999));
    InMux I__9948 (
            .O(N__44008),
            .I(N__43996));
    LocalMux I__9947 (
            .O(N__44005),
            .I(N__43993));
    Span4Mux_h I__9946 (
            .O(N__44002),
            .I(N__43990));
    LocalMux I__9945 (
            .O(N__43999),
            .I(N__43985));
    LocalMux I__9944 (
            .O(N__43996),
            .I(N__43985));
    Span4Mux_h I__9943 (
            .O(N__43993),
            .I(N__43982));
    Sp12to4 I__9942 (
            .O(N__43990),
            .I(N__43977));
    Span12Mux_h I__9941 (
            .O(N__43985),
            .I(N__43977));
    Odrv4 I__9940 (
            .O(N__43982),
            .I(\ALU.un2_addsub_cry_6_c_RNIPJK8EZ0 ));
    Odrv12 I__9939 (
            .O(N__43977),
            .I(\ALU.un2_addsub_cry_6_c_RNIPJK8EZ0 ));
    CascadeMux I__9938 (
            .O(N__43972),
            .I(N__43969));
    InMux I__9937 (
            .O(N__43969),
            .I(N__43966));
    LocalMux I__9936 (
            .O(N__43966),
            .I(\ALU.r0_12_prm_2_7_s1_c_RNOZ0 ));
    InMux I__9935 (
            .O(N__43963),
            .I(N__43958));
    InMux I__9934 (
            .O(N__43962),
            .I(N__43955));
    InMux I__9933 (
            .O(N__43961),
            .I(N__43951));
    LocalMux I__9932 (
            .O(N__43958),
            .I(N__43944));
    LocalMux I__9931 (
            .O(N__43955),
            .I(N__43941));
    CascadeMux I__9930 (
            .O(N__43954),
            .I(N__43938));
    LocalMux I__9929 (
            .O(N__43951),
            .I(N__43933));
    InMux I__9928 (
            .O(N__43950),
            .I(N__43921));
    InMux I__9927 (
            .O(N__43949),
            .I(N__43921));
    InMux I__9926 (
            .O(N__43948),
            .I(N__43921));
    InMux I__9925 (
            .O(N__43947),
            .I(N__43917));
    Span4Mux_v I__9924 (
            .O(N__43944),
            .I(N__43909));
    Span4Mux_v I__9923 (
            .O(N__43941),
            .I(N__43909));
    InMux I__9922 (
            .O(N__43938),
            .I(N__43904));
    InMux I__9921 (
            .O(N__43937),
            .I(N__43904));
    CascadeMux I__9920 (
            .O(N__43936),
            .I(N__43901));
    Span4Mux_h I__9919 (
            .O(N__43933),
            .I(N__43893));
    InMux I__9918 (
            .O(N__43932),
            .I(N__43888));
    InMux I__9917 (
            .O(N__43931),
            .I(N__43888));
    InMux I__9916 (
            .O(N__43930),
            .I(N__43883));
    InMux I__9915 (
            .O(N__43929),
            .I(N__43880));
    InMux I__9914 (
            .O(N__43928),
            .I(N__43877));
    LocalMux I__9913 (
            .O(N__43921),
            .I(N__43874));
    InMux I__9912 (
            .O(N__43920),
            .I(N__43871));
    LocalMux I__9911 (
            .O(N__43917),
            .I(N__43868));
    InMux I__9910 (
            .O(N__43916),
            .I(N__43863));
    InMux I__9909 (
            .O(N__43915),
            .I(N__43863));
    CascadeMux I__9908 (
            .O(N__43914),
            .I(N__43857));
    Span4Mux_h I__9907 (
            .O(N__43909),
            .I(N__43854));
    LocalMux I__9906 (
            .O(N__43904),
            .I(N__43851));
    InMux I__9905 (
            .O(N__43901),
            .I(N__43844));
    InMux I__9904 (
            .O(N__43900),
            .I(N__43844));
    InMux I__9903 (
            .O(N__43899),
            .I(N__43844));
    InMux I__9902 (
            .O(N__43898),
            .I(N__43841));
    InMux I__9901 (
            .O(N__43897),
            .I(N__43838));
    InMux I__9900 (
            .O(N__43896),
            .I(N__43834));
    Span4Mux_h I__9899 (
            .O(N__43893),
            .I(N__43829));
    LocalMux I__9898 (
            .O(N__43888),
            .I(N__43829));
    InMux I__9897 (
            .O(N__43887),
            .I(N__43824));
    InMux I__9896 (
            .O(N__43886),
            .I(N__43824));
    LocalMux I__9895 (
            .O(N__43883),
            .I(N__43812));
    LocalMux I__9894 (
            .O(N__43880),
            .I(N__43812));
    LocalMux I__9893 (
            .O(N__43877),
            .I(N__43809));
    Span4Mux_v I__9892 (
            .O(N__43874),
            .I(N__43804));
    LocalMux I__9891 (
            .O(N__43871),
            .I(N__43804));
    Span4Mux_v I__9890 (
            .O(N__43868),
            .I(N__43799));
    LocalMux I__9889 (
            .O(N__43863),
            .I(N__43799));
    InMux I__9888 (
            .O(N__43862),
            .I(N__43794));
    InMux I__9887 (
            .O(N__43861),
            .I(N__43794));
    InMux I__9886 (
            .O(N__43860),
            .I(N__43789));
    InMux I__9885 (
            .O(N__43857),
            .I(N__43789));
    Span4Mux_h I__9884 (
            .O(N__43854),
            .I(N__43782));
    Span4Mux_s2_h I__9883 (
            .O(N__43851),
            .I(N__43782));
    LocalMux I__9882 (
            .O(N__43844),
            .I(N__43782));
    LocalMux I__9881 (
            .O(N__43841),
            .I(N__43777));
    LocalMux I__9880 (
            .O(N__43838),
            .I(N__43777));
    InMux I__9879 (
            .O(N__43837),
            .I(N__43774));
    LocalMux I__9878 (
            .O(N__43834),
            .I(N__43767));
    Span4Mux_h I__9877 (
            .O(N__43829),
            .I(N__43767));
    LocalMux I__9876 (
            .O(N__43824),
            .I(N__43767));
    InMux I__9875 (
            .O(N__43823),
            .I(N__43760));
    InMux I__9874 (
            .O(N__43822),
            .I(N__43760));
    InMux I__9873 (
            .O(N__43821),
            .I(N__43760));
    InMux I__9872 (
            .O(N__43820),
            .I(N__43751));
    InMux I__9871 (
            .O(N__43819),
            .I(N__43751));
    InMux I__9870 (
            .O(N__43818),
            .I(N__43751));
    InMux I__9869 (
            .O(N__43817),
            .I(N__43751));
    Span4Mux_s1_v I__9868 (
            .O(N__43812),
            .I(N__43744));
    Span4Mux_h I__9867 (
            .O(N__43809),
            .I(N__43744));
    Span4Mux_h I__9866 (
            .O(N__43804),
            .I(N__43744));
    Odrv4 I__9865 (
            .O(N__43799),
            .I(\ALU.b_2 ));
    LocalMux I__9864 (
            .O(N__43794),
            .I(\ALU.b_2 ));
    LocalMux I__9863 (
            .O(N__43789),
            .I(\ALU.b_2 ));
    Odrv4 I__9862 (
            .O(N__43782),
            .I(\ALU.b_2 ));
    Odrv12 I__9861 (
            .O(N__43777),
            .I(\ALU.b_2 ));
    LocalMux I__9860 (
            .O(N__43774),
            .I(\ALU.b_2 ));
    Odrv4 I__9859 (
            .O(N__43767),
            .I(\ALU.b_2 ));
    LocalMux I__9858 (
            .O(N__43760),
            .I(\ALU.b_2 ));
    LocalMux I__9857 (
            .O(N__43751),
            .I(\ALU.b_2 ));
    Odrv4 I__9856 (
            .O(N__43744),
            .I(\ALU.b_2 ));
    CascadeMux I__9855 (
            .O(N__43723),
            .I(N__43720));
    InMux I__9854 (
            .O(N__43720),
            .I(N__43717));
    LocalMux I__9853 (
            .O(N__43717),
            .I(N__43714));
    Span4Mux_s0_v I__9852 (
            .O(N__43714),
            .I(N__43711));
    Odrv4 I__9851 (
            .O(N__43711),
            .I(\ALU.r0_12_prm_5_2_c_RNOZ0Z_0 ));
    InMux I__9850 (
            .O(N__43708),
            .I(N__43704));
    InMux I__9849 (
            .O(N__43707),
            .I(N__43701));
    LocalMux I__9848 (
            .O(N__43704),
            .I(N__43698));
    LocalMux I__9847 (
            .O(N__43701),
            .I(N__43695));
    Span4Mux_s3_v I__9846 (
            .O(N__43698),
            .I(N__43692));
    Span4Mux_s3_v I__9845 (
            .O(N__43695),
            .I(N__43689));
    Span4Mux_v I__9844 (
            .O(N__43692),
            .I(N__43686));
    Span4Mux_h I__9843 (
            .O(N__43689),
            .I(N__43683));
    Odrv4 I__9842 (
            .O(N__43686),
            .I(\ALU.un9_addsub_cry_1_c_RNIKO6AJZ0 ));
    Odrv4 I__9841 (
            .O(N__43683),
            .I(\ALU.un9_addsub_cry_1_c_RNIKO6AJZ0 ));
    CascadeMux I__9840 (
            .O(N__43678),
            .I(N__43675));
    InMux I__9839 (
            .O(N__43675),
            .I(N__43672));
    LocalMux I__9838 (
            .O(N__43672),
            .I(\ALU.r0_12_prm_1_2_c_RNOZ0 ));
    InMux I__9837 (
            .O(N__43669),
            .I(N__43661));
    InMux I__9836 (
            .O(N__43668),
            .I(N__43658));
    CascadeMux I__9835 (
            .O(N__43667),
            .I(N__43652));
    CascadeMux I__9834 (
            .O(N__43666),
            .I(N__43645));
    CascadeMux I__9833 (
            .O(N__43665),
            .I(N__43640));
    CascadeMux I__9832 (
            .O(N__43664),
            .I(N__43632));
    LocalMux I__9831 (
            .O(N__43661),
            .I(N__43628));
    LocalMux I__9830 (
            .O(N__43658),
            .I(N__43625));
    InMux I__9829 (
            .O(N__43657),
            .I(N__43622));
    InMux I__9828 (
            .O(N__43656),
            .I(N__43619));
    InMux I__9827 (
            .O(N__43655),
            .I(N__43616));
    InMux I__9826 (
            .O(N__43652),
            .I(N__43613));
    InMux I__9825 (
            .O(N__43651),
            .I(N__43608));
    InMux I__9824 (
            .O(N__43650),
            .I(N__43608));
    CascadeMux I__9823 (
            .O(N__43649),
            .I(N__43603));
    InMux I__9822 (
            .O(N__43648),
            .I(N__43600));
    InMux I__9821 (
            .O(N__43645),
            .I(N__43597));
    InMux I__9820 (
            .O(N__43644),
            .I(N__43594));
    CascadeMux I__9819 (
            .O(N__43643),
            .I(N__43591));
    InMux I__9818 (
            .O(N__43640),
            .I(N__43586));
    InMux I__9817 (
            .O(N__43639),
            .I(N__43581));
    InMux I__9816 (
            .O(N__43638),
            .I(N__43581));
    InMux I__9815 (
            .O(N__43637),
            .I(N__43576));
    InMux I__9814 (
            .O(N__43636),
            .I(N__43576));
    InMux I__9813 (
            .O(N__43635),
            .I(N__43571));
    InMux I__9812 (
            .O(N__43632),
            .I(N__43571));
    InMux I__9811 (
            .O(N__43631),
            .I(N__43567));
    Span4Mux_s3_v I__9810 (
            .O(N__43628),
            .I(N__43562));
    Span4Mux_v I__9809 (
            .O(N__43625),
            .I(N__43562));
    LocalMux I__9808 (
            .O(N__43622),
            .I(N__43559));
    LocalMux I__9807 (
            .O(N__43619),
            .I(N__43554));
    LocalMux I__9806 (
            .O(N__43616),
            .I(N__43554));
    LocalMux I__9805 (
            .O(N__43613),
            .I(N__43551));
    LocalMux I__9804 (
            .O(N__43608),
            .I(N__43548));
    InMux I__9803 (
            .O(N__43607),
            .I(N__43545));
    InMux I__9802 (
            .O(N__43606),
            .I(N__43542));
    InMux I__9801 (
            .O(N__43603),
            .I(N__43539));
    LocalMux I__9800 (
            .O(N__43600),
            .I(N__43536));
    LocalMux I__9799 (
            .O(N__43597),
            .I(N__43533));
    LocalMux I__9798 (
            .O(N__43594),
            .I(N__43530));
    InMux I__9797 (
            .O(N__43591),
            .I(N__43527));
    InMux I__9796 (
            .O(N__43590),
            .I(N__43522));
    InMux I__9795 (
            .O(N__43589),
            .I(N__43522));
    LocalMux I__9794 (
            .O(N__43586),
            .I(N__43517));
    LocalMux I__9793 (
            .O(N__43581),
            .I(N__43510));
    LocalMux I__9792 (
            .O(N__43576),
            .I(N__43510));
    LocalMux I__9791 (
            .O(N__43571),
            .I(N__43510));
    InMux I__9790 (
            .O(N__43570),
            .I(N__43507));
    LocalMux I__9789 (
            .O(N__43567),
            .I(N__43504));
    Span4Mux_h I__9788 (
            .O(N__43562),
            .I(N__43495));
    Span4Mux_s3_v I__9787 (
            .O(N__43559),
            .I(N__43495));
    Span4Mux_s3_v I__9786 (
            .O(N__43554),
            .I(N__43495));
    Span4Mux_v I__9785 (
            .O(N__43551),
            .I(N__43495));
    Span4Mux_s2_h I__9784 (
            .O(N__43548),
            .I(N__43492));
    LocalMux I__9783 (
            .O(N__43545),
            .I(N__43487));
    LocalMux I__9782 (
            .O(N__43542),
            .I(N__43487));
    LocalMux I__9781 (
            .O(N__43539),
            .I(N__43484));
    Span4Mux_h I__9780 (
            .O(N__43536),
            .I(N__43473));
    Span4Mux_h I__9779 (
            .O(N__43533),
            .I(N__43473));
    Span4Mux_s0_v I__9778 (
            .O(N__43530),
            .I(N__43473));
    LocalMux I__9777 (
            .O(N__43527),
            .I(N__43473));
    LocalMux I__9776 (
            .O(N__43522),
            .I(N__43473));
    InMux I__9775 (
            .O(N__43521),
            .I(N__43468));
    InMux I__9774 (
            .O(N__43520),
            .I(N__43468));
    Span4Mux_h I__9773 (
            .O(N__43517),
            .I(N__43463));
    Span4Mux_s3_h I__9772 (
            .O(N__43510),
            .I(N__43463));
    LocalMux I__9771 (
            .O(N__43507),
            .I(N__43460));
    Span4Mux_s2_h I__9770 (
            .O(N__43504),
            .I(N__43449));
    Span4Mux_h I__9769 (
            .O(N__43495),
            .I(N__43449));
    Span4Mux_v I__9768 (
            .O(N__43492),
            .I(N__43449));
    Span4Mux_s3_v I__9767 (
            .O(N__43487),
            .I(N__43449));
    Span4Mux_s3_v I__9766 (
            .O(N__43484),
            .I(N__43449));
    Odrv4 I__9765 (
            .O(N__43473),
            .I(\ALU.b_6 ));
    LocalMux I__9764 (
            .O(N__43468),
            .I(\ALU.b_6 ));
    Odrv4 I__9763 (
            .O(N__43463),
            .I(\ALU.b_6 ));
    Odrv4 I__9762 (
            .O(N__43460),
            .I(\ALU.b_6 ));
    Odrv4 I__9761 (
            .O(N__43449),
            .I(\ALU.b_6 ));
    InMux I__9760 (
            .O(N__43438),
            .I(N__43432));
    CascadeMux I__9759 (
            .O(N__43437),
            .I(N__43426));
    InMux I__9758 (
            .O(N__43436),
            .I(N__43421));
    InMux I__9757 (
            .O(N__43435),
            .I(N__43417));
    LocalMux I__9756 (
            .O(N__43432),
            .I(N__43412));
    CascadeMux I__9755 (
            .O(N__43431),
            .I(N__43409));
    InMux I__9754 (
            .O(N__43430),
            .I(N__43405));
    InMux I__9753 (
            .O(N__43429),
            .I(N__43400));
    InMux I__9752 (
            .O(N__43426),
            .I(N__43397));
    CascadeMux I__9751 (
            .O(N__43425),
            .I(N__43390));
    CascadeMux I__9750 (
            .O(N__43424),
            .I(N__43387));
    LocalMux I__9749 (
            .O(N__43421),
            .I(N__43384));
    InMux I__9748 (
            .O(N__43420),
            .I(N__43381));
    LocalMux I__9747 (
            .O(N__43417),
            .I(N__43372));
    InMux I__9746 (
            .O(N__43416),
            .I(N__43369));
    InMux I__9745 (
            .O(N__43415),
            .I(N__43366));
    Span4Mux_v I__9744 (
            .O(N__43412),
            .I(N__43362));
    InMux I__9743 (
            .O(N__43409),
            .I(N__43359));
    InMux I__9742 (
            .O(N__43408),
            .I(N__43356));
    LocalMux I__9741 (
            .O(N__43405),
            .I(N__43352));
    InMux I__9740 (
            .O(N__43404),
            .I(N__43347));
    InMux I__9739 (
            .O(N__43403),
            .I(N__43347));
    LocalMux I__9738 (
            .O(N__43400),
            .I(N__43344));
    LocalMux I__9737 (
            .O(N__43397),
            .I(N__43341));
    InMux I__9736 (
            .O(N__43396),
            .I(N__43338));
    InMux I__9735 (
            .O(N__43395),
            .I(N__43333));
    InMux I__9734 (
            .O(N__43394),
            .I(N__43333));
    InMux I__9733 (
            .O(N__43393),
            .I(N__43330));
    InMux I__9732 (
            .O(N__43390),
            .I(N__43325));
    InMux I__9731 (
            .O(N__43387),
            .I(N__43325));
    Span4Mux_h I__9730 (
            .O(N__43384),
            .I(N__43320));
    LocalMux I__9729 (
            .O(N__43381),
            .I(N__43320));
    InMux I__9728 (
            .O(N__43380),
            .I(N__43315));
    InMux I__9727 (
            .O(N__43379),
            .I(N__43315));
    InMux I__9726 (
            .O(N__43378),
            .I(N__43310));
    InMux I__9725 (
            .O(N__43377),
            .I(N__43310));
    InMux I__9724 (
            .O(N__43376),
            .I(N__43303));
    InMux I__9723 (
            .O(N__43375),
            .I(N__43303));
    Span4Mux_v I__9722 (
            .O(N__43372),
            .I(N__43300));
    LocalMux I__9721 (
            .O(N__43369),
            .I(N__43297));
    LocalMux I__9720 (
            .O(N__43366),
            .I(N__43294));
    InMux I__9719 (
            .O(N__43365),
            .I(N__43291));
    Span4Mux_h I__9718 (
            .O(N__43362),
            .I(N__43284));
    LocalMux I__9717 (
            .O(N__43359),
            .I(N__43284));
    LocalMux I__9716 (
            .O(N__43356),
            .I(N__43284));
    CascadeMux I__9715 (
            .O(N__43355),
            .I(N__43276));
    Span4Mux_h I__9714 (
            .O(N__43352),
            .I(N__43269));
    LocalMux I__9713 (
            .O(N__43347),
            .I(N__43269));
    Span4Mux_s1_v I__9712 (
            .O(N__43344),
            .I(N__43269));
    Span4Mux_h I__9711 (
            .O(N__43341),
            .I(N__43266));
    LocalMux I__9710 (
            .O(N__43338),
            .I(N__43261));
    LocalMux I__9709 (
            .O(N__43333),
            .I(N__43261));
    LocalMux I__9708 (
            .O(N__43330),
            .I(N__43258));
    LocalMux I__9707 (
            .O(N__43325),
            .I(N__43255));
    Span4Mux_h I__9706 (
            .O(N__43320),
            .I(N__43252));
    LocalMux I__9705 (
            .O(N__43315),
            .I(N__43247));
    LocalMux I__9704 (
            .O(N__43310),
            .I(N__43247));
    InMux I__9703 (
            .O(N__43309),
            .I(N__43242));
    InMux I__9702 (
            .O(N__43308),
            .I(N__43242));
    LocalMux I__9701 (
            .O(N__43303),
            .I(N__43239));
    Span4Mux_h I__9700 (
            .O(N__43300),
            .I(N__43228));
    Span4Mux_s1_v I__9699 (
            .O(N__43297),
            .I(N__43228));
    Span4Mux_v I__9698 (
            .O(N__43294),
            .I(N__43228));
    LocalMux I__9697 (
            .O(N__43291),
            .I(N__43228));
    Span4Mux_v I__9696 (
            .O(N__43284),
            .I(N__43228));
    InMux I__9695 (
            .O(N__43283),
            .I(N__43221));
    InMux I__9694 (
            .O(N__43282),
            .I(N__43221));
    InMux I__9693 (
            .O(N__43281),
            .I(N__43221));
    InMux I__9692 (
            .O(N__43280),
            .I(N__43218));
    InMux I__9691 (
            .O(N__43279),
            .I(N__43213));
    InMux I__9690 (
            .O(N__43276),
            .I(N__43213));
    Span4Mux_h I__9689 (
            .O(N__43269),
            .I(N__43202));
    Span4Mux_v I__9688 (
            .O(N__43266),
            .I(N__43202));
    Span4Mux_v I__9687 (
            .O(N__43261),
            .I(N__43202));
    Span4Mux_s3_h I__9686 (
            .O(N__43258),
            .I(N__43202));
    Span4Mux_v I__9685 (
            .O(N__43255),
            .I(N__43202));
    Span4Mux_h I__9684 (
            .O(N__43252),
            .I(N__43199));
    Span12Mux_v I__9683 (
            .O(N__43247),
            .I(N__43194));
    LocalMux I__9682 (
            .O(N__43242),
            .I(N__43194));
    Span4Mux_v I__9681 (
            .O(N__43239),
            .I(N__43189));
    Span4Mux_h I__9680 (
            .O(N__43228),
            .I(N__43189));
    LocalMux I__9679 (
            .O(N__43221),
            .I(\ALU.a_6 ));
    LocalMux I__9678 (
            .O(N__43218),
            .I(\ALU.a_6 ));
    LocalMux I__9677 (
            .O(N__43213),
            .I(\ALU.a_6 ));
    Odrv4 I__9676 (
            .O(N__43202),
            .I(\ALU.a_6 ));
    Odrv4 I__9675 (
            .O(N__43199),
            .I(\ALU.a_6 ));
    Odrv12 I__9674 (
            .O(N__43194),
            .I(\ALU.a_6 ));
    Odrv4 I__9673 (
            .O(N__43189),
            .I(\ALU.a_6 ));
    CascadeMux I__9672 (
            .O(N__43174),
            .I(N__43171));
    InMux I__9671 (
            .O(N__43171),
            .I(N__43168));
    LocalMux I__9670 (
            .O(N__43168),
            .I(N__43165));
    Span4Mux_h I__9669 (
            .O(N__43165),
            .I(N__43162));
    Odrv4 I__9668 (
            .O(N__43162),
            .I(\ALU.r0_12_prm_5_6_s0_c_RNOZ0 ));
    CascadeMux I__9667 (
            .O(N__43159),
            .I(N__43156));
    InMux I__9666 (
            .O(N__43156),
            .I(N__43153));
    LocalMux I__9665 (
            .O(N__43153),
            .I(N__43150));
    Span12Mux_v I__9664 (
            .O(N__43150),
            .I(N__43147));
    Odrv12 I__9663 (
            .O(N__43147),
            .I(\ALU.r0_12_prm_5_7_s0_c_RNOZ0 ));
    InMux I__9662 (
            .O(N__43144),
            .I(N__43141));
    LocalMux I__9661 (
            .O(N__43141),
            .I(N__43135));
    InMux I__9660 (
            .O(N__43140),
            .I(N__43132));
    InMux I__9659 (
            .O(N__43139),
            .I(N__43129));
    InMux I__9658 (
            .O(N__43138),
            .I(N__43124));
    Span4Mux_h I__9657 (
            .O(N__43135),
            .I(N__43118));
    LocalMux I__9656 (
            .O(N__43132),
            .I(N__43118));
    LocalMux I__9655 (
            .O(N__43129),
            .I(N__43115));
    InMux I__9654 (
            .O(N__43128),
            .I(N__43112));
    InMux I__9653 (
            .O(N__43127),
            .I(N__43109));
    LocalMux I__9652 (
            .O(N__43124),
            .I(N__43106));
    InMux I__9651 (
            .O(N__43123),
            .I(N__43103));
    Span4Mux_v I__9650 (
            .O(N__43118),
            .I(N__43100));
    Span4Mux_v I__9649 (
            .O(N__43115),
            .I(N__43097));
    LocalMux I__9648 (
            .O(N__43112),
            .I(N__43092));
    LocalMux I__9647 (
            .O(N__43109),
            .I(N__43092));
    Span12Mux_h I__9646 (
            .O(N__43106),
            .I(N__43089));
    LocalMux I__9645 (
            .O(N__43103),
            .I(N__43086));
    Span4Mux_v I__9644 (
            .O(N__43100),
            .I(N__43079));
    Span4Mux_h I__9643 (
            .O(N__43097),
            .I(N__43079));
    Span4Mux_v I__9642 (
            .O(N__43092),
            .I(N__43079));
    Span12Mux_v I__9641 (
            .O(N__43089),
            .I(N__43076));
    Span12Mux_v I__9640 (
            .O(N__43086),
            .I(N__43071));
    Sp12to4 I__9639 (
            .O(N__43079),
            .I(N__43071));
    Odrv12 I__9638 (
            .O(N__43076),
            .I(\ALU.r5_RNILM5AEZ0Z_15 ));
    Odrv12 I__9637 (
            .O(N__43071),
            .I(\ALU.r5_RNILM5AEZ0Z_15 ));
    InMux I__9636 (
            .O(N__43066),
            .I(N__43062));
    InMux I__9635 (
            .O(N__43065),
            .I(N__43059));
    LocalMux I__9634 (
            .O(N__43062),
            .I(N__43056));
    LocalMux I__9633 (
            .O(N__43059),
            .I(N__43049));
    Span4Mux_v I__9632 (
            .O(N__43056),
            .I(N__43049));
    InMux I__9631 (
            .O(N__43055),
            .I(N__43046));
    InMux I__9630 (
            .O(N__43054),
            .I(N__43043));
    Span4Mux_v I__9629 (
            .O(N__43049),
            .I(N__43038));
    LocalMux I__9628 (
            .O(N__43046),
            .I(N__43038));
    LocalMux I__9627 (
            .O(N__43043),
            .I(\ALU.r5_RNILV3HJZ0Z_12 ));
    Odrv4 I__9626 (
            .O(N__43038),
            .I(\ALU.r5_RNILV3HJZ0Z_12 ));
    InMux I__9625 (
            .O(N__43033),
            .I(N__43030));
    LocalMux I__9624 (
            .O(N__43030),
            .I(N__43027));
    Span4Mux_v I__9623 (
            .O(N__43027),
            .I(N__43024));
    Span4Mux_v I__9622 (
            .O(N__43024),
            .I(N__43021));
    Span4Mux_s2_v I__9621 (
            .O(N__43021),
            .I(N__43018));
    Span4Mux_h I__9620 (
            .O(N__43018),
            .I(N__43015));
    Odrv4 I__9619 (
            .O(N__43015),
            .I(\ALU.rshift_9 ));
    InMux I__9618 (
            .O(N__43012),
            .I(N__43007));
    InMux I__9617 (
            .O(N__43011),
            .I(N__43004));
    InMux I__9616 (
            .O(N__43010),
            .I(N__43001));
    LocalMux I__9615 (
            .O(N__43007),
            .I(N__42998));
    LocalMux I__9614 (
            .O(N__43004),
            .I(N__42993));
    LocalMux I__9613 (
            .O(N__43001),
            .I(N__42993));
    Odrv12 I__9612 (
            .O(N__42998),
            .I(\ALU.r4_RNI9H7SJZ0Z_5 ));
    Odrv12 I__9611 (
            .O(N__42993),
            .I(\ALU.r4_RNI9H7SJZ0Z_5 ));
    CascadeMux I__9610 (
            .O(N__42988),
            .I(\ALU.lshift_7_cascade_ ));
    InMux I__9609 (
            .O(N__42985),
            .I(N__42982));
    LocalMux I__9608 (
            .O(N__42982),
            .I(N__42979));
    Span4Mux_h I__9607 (
            .O(N__42979),
            .I(N__42976));
    Odrv4 I__9606 (
            .O(N__42976),
            .I(\ALU.r0_12_prm_8_7_s0_c_RNOZ0 ));
    InMux I__9605 (
            .O(N__42973),
            .I(\ALU.r0_12_s1_9 ));
    InMux I__9604 (
            .O(N__42970),
            .I(N__42967));
    LocalMux I__9603 (
            .O(N__42967),
            .I(N__42964));
    Span4Mux_h I__9602 (
            .O(N__42964),
            .I(N__42961));
    Span4Mux_h I__9601 (
            .O(N__42961),
            .I(N__42958));
    Odrv4 I__9600 (
            .O(N__42958),
            .I(\ALU.r0_12_s1_9_THRU_CO ));
    CascadeMux I__9599 (
            .O(N__42955),
            .I(N__42952));
    InMux I__9598 (
            .O(N__42952),
            .I(N__42949));
    LocalMux I__9597 (
            .O(N__42949),
            .I(N__42946));
    Span4Mux_v I__9596 (
            .O(N__42946),
            .I(N__42943));
    Span4Mux_h I__9595 (
            .O(N__42943),
            .I(N__42940));
    Odrv4 I__9594 (
            .O(N__42940),
            .I(\ALU.r0_12_prm_7_14_s0_c_RNOZ0 ));
    CascadeMux I__9593 (
            .O(N__42937),
            .I(N__42934));
    InMux I__9592 (
            .O(N__42934),
            .I(N__42931));
    LocalMux I__9591 (
            .O(N__42931),
            .I(N__42928));
    Odrv4 I__9590 (
            .O(N__42928),
            .I(\ALU.un14_log_0_i_2 ));
    CascadeMux I__9589 (
            .O(N__42925),
            .I(N__42922));
    InMux I__9588 (
            .O(N__42922),
            .I(N__42919));
    LocalMux I__9587 (
            .O(N__42919),
            .I(\ALU.mult_2 ));
    InMux I__9586 (
            .O(N__42916),
            .I(N__42910));
    InMux I__9585 (
            .O(N__42915),
            .I(N__42910));
    LocalMux I__9584 (
            .O(N__42910),
            .I(N__42907));
    Span4Mux_h I__9583 (
            .O(N__42907),
            .I(N__42904));
    Span4Mux_h I__9582 (
            .O(N__42904),
            .I(N__42901));
    Odrv4 I__9581 (
            .O(N__42901),
            .I(\ALU.madd_cry_0_THRU_CO ));
    InMux I__9580 (
            .O(N__42898),
            .I(N__42893));
    InMux I__9579 (
            .O(N__42897),
            .I(N__42888));
    InMux I__9578 (
            .O(N__42896),
            .I(N__42888));
    LocalMux I__9577 (
            .O(N__42893),
            .I(N__42885));
    LocalMux I__9576 (
            .O(N__42888),
            .I(N__42882));
    Span4Mux_v I__9575 (
            .O(N__42885),
            .I(N__42879));
    Odrv12 I__9574 (
            .O(N__42882),
            .I(\ALU.madd_axb_1 ));
    Odrv4 I__9573 (
            .O(N__42879),
            .I(\ALU.madd_axb_1 ));
    InMux I__9572 (
            .O(N__42874),
            .I(N__42871));
    LocalMux I__9571 (
            .O(N__42871),
            .I(\ALU.r0_12_prm_3_2_c_RNOZ0 ));
    CascadeMux I__9570 (
            .O(N__42868),
            .I(N__42863));
    InMux I__9569 (
            .O(N__42867),
            .I(N__42858));
    InMux I__9568 (
            .O(N__42866),
            .I(N__42855));
    InMux I__9567 (
            .O(N__42863),
            .I(N__42852));
    CascadeMux I__9566 (
            .O(N__42862),
            .I(N__42845));
    InMux I__9565 (
            .O(N__42861),
            .I(N__42839));
    LocalMux I__9564 (
            .O(N__42858),
            .I(N__42834));
    LocalMux I__9563 (
            .O(N__42855),
            .I(N__42831));
    LocalMux I__9562 (
            .O(N__42852),
            .I(N__42828));
    InMux I__9561 (
            .O(N__42851),
            .I(N__42822));
    InMux I__9560 (
            .O(N__42850),
            .I(N__42819));
    InMux I__9559 (
            .O(N__42849),
            .I(N__42812));
    InMux I__9558 (
            .O(N__42848),
            .I(N__42809));
    InMux I__9557 (
            .O(N__42845),
            .I(N__42804));
    InMux I__9556 (
            .O(N__42844),
            .I(N__42804));
    InMux I__9555 (
            .O(N__42843),
            .I(N__42801));
    InMux I__9554 (
            .O(N__42842),
            .I(N__42798));
    LocalMux I__9553 (
            .O(N__42839),
            .I(N__42795));
    InMux I__9552 (
            .O(N__42838),
            .I(N__42792));
    InMux I__9551 (
            .O(N__42837),
            .I(N__42789));
    Span4Mux_v I__9550 (
            .O(N__42834),
            .I(N__42782));
    Span4Mux_s2_v I__9549 (
            .O(N__42831),
            .I(N__42782));
    Span4Mux_v I__9548 (
            .O(N__42828),
            .I(N__42779));
    InMux I__9547 (
            .O(N__42827),
            .I(N__42774));
    InMux I__9546 (
            .O(N__42826),
            .I(N__42774));
    InMux I__9545 (
            .O(N__42825),
            .I(N__42771));
    LocalMux I__9544 (
            .O(N__42822),
            .I(N__42766));
    LocalMux I__9543 (
            .O(N__42819),
            .I(N__42766));
    InMux I__9542 (
            .O(N__42818),
            .I(N__42759));
    InMux I__9541 (
            .O(N__42817),
            .I(N__42759));
    InMux I__9540 (
            .O(N__42816),
            .I(N__42759));
    InMux I__9539 (
            .O(N__42815),
            .I(N__42756));
    LocalMux I__9538 (
            .O(N__42812),
            .I(N__42747));
    LocalMux I__9537 (
            .O(N__42809),
            .I(N__42747));
    LocalMux I__9536 (
            .O(N__42804),
            .I(N__42744));
    LocalMux I__9535 (
            .O(N__42801),
            .I(N__42739));
    LocalMux I__9534 (
            .O(N__42798),
            .I(N__42739));
    Span4Mux_h I__9533 (
            .O(N__42795),
            .I(N__42734));
    LocalMux I__9532 (
            .O(N__42792),
            .I(N__42734));
    LocalMux I__9531 (
            .O(N__42789),
            .I(N__42731));
    InMux I__9530 (
            .O(N__42788),
            .I(N__42728));
    CascadeMux I__9529 (
            .O(N__42787),
            .I(N__42720));
    Span4Mux_h I__9528 (
            .O(N__42782),
            .I(N__42715));
    Span4Mux_v I__9527 (
            .O(N__42779),
            .I(N__42715));
    LocalMux I__9526 (
            .O(N__42774),
            .I(N__42712));
    LocalMux I__9525 (
            .O(N__42771),
            .I(N__42705));
    Span4Mux_v I__9524 (
            .O(N__42766),
            .I(N__42705));
    LocalMux I__9523 (
            .O(N__42759),
            .I(N__42705));
    LocalMux I__9522 (
            .O(N__42756),
            .I(N__42702));
    CascadeMux I__9521 (
            .O(N__42755),
            .I(N__42699));
    CascadeMux I__9520 (
            .O(N__42754),
            .I(N__42696));
    InMux I__9519 (
            .O(N__42753),
            .I(N__42691));
    InMux I__9518 (
            .O(N__42752),
            .I(N__42691));
    Span4Mux_h I__9517 (
            .O(N__42747),
            .I(N__42686));
    Span4Mux_v I__9516 (
            .O(N__42744),
            .I(N__42686));
    Span4Mux_v I__9515 (
            .O(N__42739),
            .I(N__42683));
    Span4Mux_v I__9514 (
            .O(N__42734),
            .I(N__42678));
    Span4Mux_h I__9513 (
            .O(N__42731),
            .I(N__42678));
    LocalMux I__9512 (
            .O(N__42728),
            .I(N__42675));
    InMux I__9511 (
            .O(N__42727),
            .I(N__42670));
    InMux I__9510 (
            .O(N__42726),
            .I(N__42670));
    InMux I__9509 (
            .O(N__42725),
            .I(N__42663));
    InMux I__9508 (
            .O(N__42724),
            .I(N__42663));
    InMux I__9507 (
            .O(N__42723),
            .I(N__42663));
    InMux I__9506 (
            .O(N__42720),
            .I(N__42660));
    Span4Mux_h I__9505 (
            .O(N__42715),
            .I(N__42655));
    Span4Mux_s2_h I__9504 (
            .O(N__42712),
            .I(N__42655));
    Span4Mux_h I__9503 (
            .O(N__42705),
            .I(N__42650));
    Span4Mux_s2_v I__9502 (
            .O(N__42702),
            .I(N__42650));
    InMux I__9501 (
            .O(N__42699),
            .I(N__42645));
    InMux I__9500 (
            .O(N__42696),
            .I(N__42645));
    LocalMux I__9499 (
            .O(N__42691),
            .I(N__42642));
    Span4Mux_h I__9498 (
            .O(N__42686),
            .I(N__42635));
    Span4Mux_h I__9497 (
            .O(N__42683),
            .I(N__42635));
    Span4Mux_h I__9496 (
            .O(N__42678),
            .I(N__42635));
    Odrv4 I__9495 (
            .O(N__42675),
            .I(\ALU.a_4 ));
    LocalMux I__9494 (
            .O(N__42670),
            .I(\ALU.a_4 ));
    LocalMux I__9493 (
            .O(N__42663),
            .I(\ALU.a_4 ));
    LocalMux I__9492 (
            .O(N__42660),
            .I(\ALU.a_4 ));
    Odrv4 I__9491 (
            .O(N__42655),
            .I(\ALU.a_4 ));
    Odrv4 I__9490 (
            .O(N__42650),
            .I(\ALU.a_4 ));
    LocalMux I__9489 (
            .O(N__42645),
            .I(\ALU.a_4 ));
    Odrv12 I__9488 (
            .O(N__42642),
            .I(\ALU.a_4 ));
    Odrv4 I__9487 (
            .O(N__42635),
            .I(\ALU.a_4 ));
    CascadeMux I__9486 (
            .O(N__42616),
            .I(N__42613));
    InMux I__9485 (
            .O(N__42613),
            .I(N__42610));
    LocalMux I__9484 (
            .O(N__42610),
            .I(N__42607));
    Span4Mux_v I__9483 (
            .O(N__42607),
            .I(N__42604));
    Odrv4 I__9482 (
            .O(N__42604),
            .I(\ALU.r4_RNI87HO5Z0Z_4 ));
    InMux I__9481 (
            .O(N__42601),
            .I(N__42598));
    LocalMux I__9480 (
            .O(N__42598),
            .I(N__42595));
    Span4Mux_h I__9479 (
            .O(N__42595),
            .I(N__42592));
    Span4Mux_v I__9478 (
            .O(N__42592),
            .I(N__42589));
    Odrv4 I__9477 (
            .O(N__42589),
            .I(\ALU.r0_12_prm_8_9_s1_c_RNOZ0 ));
    InMux I__9476 (
            .O(N__42586),
            .I(N__42582));
    CascadeMux I__9475 (
            .O(N__42585),
            .I(N__42579));
    LocalMux I__9474 (
            .O(N__42582),
            .I(N__42576));
    InMux I__9473 (
            .O(N__42579),
            .I(N__42573));
    Span4Mux_v I__9472 (
            .O(N__42576),
            .I(N__42570));
    LocalMux I__9471 (
            .O(N__42573),
            .I(N__42567));
    Span4Mux_h I__9470 (
            .O(N__42570),
            .I(N__42562));
    Span4Mux_h I__9469 (
            .O(N__42567),
            .I(N__42562));
    Span4Mux_v I__9468 (
            .O(N__42562),
            .I(N__42558));
    InMux I__9467 (
            .O(N__42561),
            .I(N__42555));
    Odrv4 I__9466 (
            .O(N__42558),
            .I(\ALU.lshift_9 ));
    LocalMux I__9465 (
            .O(N__42555),
            .I(\ALU.lshift_9 ));
    InMux I__9464 (
            .O(N__42550),
            .I(N__42547));
    LocalMux I__9463 (
            .O(N__42547),
            .I(N__42544));
    Odrv4 I__9462 (
            .O(N__42544),
            .I(\ALU.r0_12_prm_7_9_s1_c_RNOZ0 ));
    InMux I__9461 (
            .O(N__42541),
            .I(N__42537));
    CascadeMux I__9460 (
            .O(N__42540),
            .I(N__42534));
    LocalMux I__9459 (
            .O(N__42537),
            .I(N__42531));
    InMux I__9458 (
            .O(N__42534),
            .I(N__42528));
    Span4Mux_h I__9457 (
            .O(N__42531),
            .I(N__42525));
    LocalMux I__9456 (
            .O(N__42528),
            .I(N__42522));
    Odrv4 I__9455 (
            .O(N__42525),
            .I(\ALU.r4_RNISU5D9_0Z0Z_9 ));
    Odrv4 I__9454 (
            .O(N__42522),
            .I(\ALU.r4_RNISU5D9_0Z0Z_9 ));
    InMux I__9453 (
            .O(N__42517),
            .I(N__42514));
    LocalMux I__9452 (
            .O(N__42514),
            .I(N__42511));
    Odrv4 I__9451 (
            .O(N__42511),
            .I(\ALU.r0_12_prm_6_9_s1_c_RNOZ0 ));
    InMux I__9450 (
            .O(N__42508),
            .I(N__42504));
    InMux I__9449 (
            .O(N__42507),
            .I(N__42501));
    LocalMux I__9448 (
            .O(N__42504),
            .I(N__42498));
    LocalMux I__9447 (
            .O(N__42501),
            .I(N__42495));
    Span4Mux_h I__9446 (
            .O(N__42498),
            .I(N__42492));
    Odrv4 I__9445 (
            .O(N__42495),
            .I(\ALU.r4_RNISU5D9_1Z0Z_9 ));
    Odrv4 I__9444 (
            .O(N__42492),
            .I(\ALU.r4_RNISU5D9_1Z0Z_9 ));
    CascadeMux I__9443 (
            .O(N__42487),
            .I(N__42484));
    InMux I__9442 (
            .O(N__42484),
            .I(N__42481));
    LocalMux I__9441 (
            .O(N__42481),
            .I(\ALU.r0_12_prm_5_9_s1_c_RNOZ0 ));
    CascadeMux I__9440 (
            .O(N__42478),
            .I(N__42475));
    InMux I__9439 (
            .O(N__42475),
            .I(N__42472));
    LocalMux I__9438 (
            .O(N__42472),
            .I(N__42469));
    Span4Mux_v I__9437 (
            .O(N__42469),
            .I(N__42465));
    InMux I__9436 (
            .O(N__42468),
            .I(N__42462));
    Span4Mux_h I__9435 (
            .O(N__42465),
            .I(N__42459));
    LocalMux I__9434 (
            .O(N__42462),
            .I(\ALU.a_i_9 ));
    Odrv4 I__9433 (
            .O(N__42459),
            .I(\ALU.a_i_9 ));
    InMux I__9432 (
            .O(N__42454),
            .I(N__42451));
    LocalMux I__9431 (
            .O(N__42451),
            .I(\ALU.r0_12_prm_2_9_s1_c_RNOZ0 ));
    InMux I__9430 (
            .O(N__42448),
            .I(N__42444));
    CascadeMux I__9429 (
            .O(N__42447),
            .I(N__42441));
    LocalMux I__9428 (
            .O(N__42444),
            .I(N__42437));
    InMux I__9427 (
            .O(N__42441),
            .I(N__42434));
    InMux I__9426 (
            .O(N__42440),
            .I(N__42431));
    Span4Mux_h I__9425 (
            .O(N__42437),
            .I(N__42427));
    LocalMux I__9424 (
            .O(N__42434),
            .I(N__42422));
    LocalMux I__9423 (
            .O(N__42431),
            .I(N__42422));
    InMux I__9422 (
            .O(N__42430),
            .I(N__42419));
    Span4Mux_h I__9421 (
            .O(N__42427),
            .I(N__42416));
    Span4Mux_h I__9420 (
            .O(N__42422),
            .I(N__42413));
    LocalMux I__9419 (
            .O(N__42419),
            .I(\ALU.un2_addsub_cry_8_c_RNINO51FZ0 ));
    Odrv4 I__9418 (
            .O(N__42416),
            .I(\ALU.un2_addsub_cry_8_c_RNINO51FZ0 ));
    Odrv4 I__9417 (
            .O(N__42413),
            .I(\ALU.un2_addsub_cry_8_c_RNINO51FZ0 ));
    InMux I__9416 (
            .O(N__42406),
            .I(N__42403));
    LocalMux I__9415 (
            .O(N__42403),
            .I(\ALU.r0_12_prm_1_9_s1_c_RNOZ0 ));
    CascadeMux I__9414 (
            .O(N__42400),
            .I(N__42396));
    InMux I__9413 (
            .O(N__42399),
            .I(N__42392));
    InMux I__9412 (
            .O(N__42396),
            .I(N__42388));
    InMux I__9411 (
            .O(N__42395),
            .I(N__42385));
    LocalMux I__9410 (
            .O(N__42392),
            .I(N__42382));
    InMux I__9409 (
            .O(N__42391),
            .I(N__42379));
    LocalMux I__9408 (
            .O(N__42388),
            .I(N__42374));
    LocalMux I__9407 (
            .O(N__42385),
            .I(N__42374));
    Span4Mux_h I__9406 (
            .O(N__42382),
            .I(N__42369));
    LocalMux I__9405 (
            .O(N__42379),
            .I(N__42369));
    Span4Mux_v I__9404 (
            .O(N__42374),
            .I(N__42366));
    Odrv4 I__9403 (
            .O(N__42369),
            .I(\ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9 ));
    Odrv4 I__9402 (
            .O(N__42366),
            .I(\ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9 ));
    InMux I__9401 (
            .O(N__42361),
            .I(N__42358));
    LocalMux I__9400 (
            .O(N__42358),
            .I(N__42355));
    Span4Mux_v I__9399 (
            .O(N__42355),
            .I(N__42352));
    Odrv4 I__9398 (
            .O(N__42352),
            .I(\ALU.lshift_3_ns_1_10 ));
    CascadeMux I__9397 (
            .O(N__42349),
            .I(\ALU.r4_RNI67NNKZ0Z_7_cascade_ ));
    CascadeMux I__9396 (
            .O(N__42346),
            .I(N__42343));
    InMux I__9395 (
            .O(N__42343),
            .I(N__42339));
    InMux I__9394 (
            .O(N__42342),
            .I(N__42336));
    LocalMux I__9393 (
            .O(N__42339),
            .I(N__42333));
    LocalMux I__9392 (
            .O(N__42336),
            .I(N__42330));
    Span4Mux_v I__9391 (
            .O(N__42333),
            .I(N__42327));
    Odrv12 I__9390 (
            .O(N__42330),
            .I(\ALU.lshift_10 ));
    Odrv4 I__9389 (
            .O(N__42327),
            .I(\ALU.lshift_10 ));
    InMux I__9388 (
            .O(N__42322),
            .I(N__42318));
    InMux I__9387 (
            .O(N__42321),
            .I(N__42313));
    LocalMux I__9386 (
            .O(N__42318),
            .I(N__42310));
    InMux I__9385 (
            .O(N__42317),
            .I(N__42305));
    InMux I__9384 (
            .O(N__42316),
            .I(N__42305));
    LocalMux I__9383 (
            .O(N__42313),
            .I(\ALU.N_610_1 ));
    Odrv12 I__9382 (
            .O(N__42310),
            .I(\ALU.N_610_1 ));
    LocalMux I__9381 (
            .O(N__42305),
            .I(\ALU.N_610_1 ));
    InMux I__9380 (
            .O(N__42298),
            .I(N__42295));
    LocalMux I__9379 (
            .O(N__42295),
            .I(N__42291));
    InMux I__9378 (
            .O(N__42294),
            .I(N__42288));
    Odrv12 I__9377 (
            .O(N__42291),
            .I(\ALU.r4_RNIAHIIAZ0Z_2 ));
    LocalMux I__9376 (
            .O(N__42288),
            .I(\ALU.r4_RNIAHIIAZ0Z_2 ));
    CascadeMux I__9375 (
            .O(N__42283),
            .I(N__42280));
    InMux I__9374 (
            .O(N__42280),
            .I(N__42274));
    InMux I__9373 (
            .O(N__42279),
            .I(N__42274));
    LocalMux I__9372 (
            .O(N__42274),
            .I(\ALU.r4_RNI38O1GZ0Z_2 ));
    CascadeMux I__9371 (
            .O(N__42271),
            .I(\ALU.r4_RNI38O1GZ0Z_2_cascade_ ));
    InMux I__9370 (
            .O(N__42268),
            .I(N__42259));
    InMux I__9369 (
            .O(N__42267),
            .I(N__42259));
    InMux I__9368 (
            .O(N__42266),
            .I(N__42259));
    LocalMux I__9367 (
            .O(N__42259),
            .I(\ALU.r4_RNICN8R81Z0Z_7 ));
    InMux I__9366 (
            .O(N__42256),
            .I(N__42253));
    LocalMux I__9365 (
            .O(N__42253),
            .I(N__42250));
    Span4Mux_v I__9364 (
            .O(N__42250),
            .I(N__42247));
    Odrv4 I__9363 (
            .O(N__42247),
            .I(\ALU.r0_12_prm_8_10_s1_c_RNOZ0 ));
    InMux I__9362 (
            .O(N__42244),
            .I(N__42241));
    LocalMux I__9361 (
            .O(N__42241),
            .I(\ALU.r4_RNI67NNKZ0Z_7 ));
    InMux I__9360 (
            .O(N__42238),
            .I(N__42235));
    LocalMux I__9359 (
            .O(N__42235),
            .I(\ALU.r5_RNI355TIZ0Z_13 ));
    InMux I__9358 (
            .O(N__42232),
            .I(N__42226));
    InMux I__9357 (
            .O(N__42231),
            .I(N__42226));
    LocalMux I__9356 (
            .O(N__42226),
            .I(N__42223));
    Span4Mux_v I__9355 (
            .O(N__42223),
            .I(N__42219));
    InMux I__9354 (
            .O(N__42222),
            .I(N__42216));
    Span4Mux_v I__9353 (
            .O(N__42219),
            .I(N__42213));
    LocalMux I__9352 (
            .O(N__42216),
            .I(\ALU.r4_RNIO7CSJZ0Z_4 ));
    Odrv4 I__9351 (
            .O(N__42213),
            .I(\ALU.r4_RNIO7CSJZ0Z_4 ));
    CascadeMux I__9350 (
            .O(N__42208),
            .I(\ALU.lshift_15_ns_1_14_cascade_ ));
    InMux I__9349 (
            .O(N__42205),
            .I(N__42200));
    InMux I__9348 (
            .O(N__42204),
            .I(N__42194));
    InMux I__9347 (
            .O(N__42203),
            .I(N__42194));
    LocalMux I__9346 (
            .O(N__42200),
            .I(N__42191));
    InMux I__9345 (
            .O(N__42199),
            .I(N__42188));
    LocalMux I__9344 (
            .O(N__42194),
            .I(N__42185));
    Span4Mux_h I__9343 (
            .O(N__42191),
            .I(N__42182));
    LocalMux I__9342 (
            .O(N__42188),
            .I(N__42179));
    Odrv12 I__9341 (
            .O(N__42185),
            .I(\ALU.r4_RNILVIQFZ0Z_2 ));
    Odrv4 I__9340 (
            .O(N__42182),
            .I(\ALU.r4_RNILVIQFZ0Z_2 ));
    Odrv12 I__9339 (
            .O(N__42179),
            .I(\ALU.r4_RNILVIQFZ0Z_2 ));
    InMux I__9338 (
            .O(N__42172),
            .I(N__42169));
    LocalMux I__9337 (
            .O(N__42169),
            .I(\ALU.r0_12_prm_8_9_s1_c_RNOZ0Z_1 ));
    InMux I__9336 (
            .O(N__42166),
            .I(\ALU.r0_12_1 ));
    InMux I__9335 (
            .O(N__42163),
            .I(N__42160));
    LocalMux I__9334 (
            .O(N__42160),
            .I(N__42157));
    Span4Mux_v I__9333 (
            .O(N__42157),
            .I(N__42151));
    InMux I__9332 (
            .O(N__42156),
            .I(N__42148));
    InMux I__9331 (
            .O(N__42155),
            .I(N__42144));
    InMux I__9330 (
            .O(N__42154),
            .I(N__42140));
    Span4Mux_h I__9329 (
            .O(N__42151),
            .I(N__42136));
    LocalMux I__9328 (
            .O(N__42148),
            .I(N__42133));
    InMux I__9327 (
            .O(N__42147),
            .I(N__42130));
    LocalMux I__9326 (
            .O(N__42144),
            .I(N__42126));
    InMux I__9325 (
            .O(N__42143),
            .I(N__42123));
    LocalMux I__9324 (
            .O(N__42140),
            .I(N__42120));
    InMux I__9323 (
            .O(N__42139),
            .I(N__42117));
    Span4Mux_v I__9322 (
            .O(N__42136),
            .I(N__42112));
    Span4Mux_h I__9321 (
            .O(N__42133),
            .I(N__42112));
    LocalMux I__9320 (
            .O(N__42130),
            .I(N__42109));
    InMux I__9319 (
            .O(N__42129),
            .I(N__42106));
    Span4Mux_h I__9318 (
            .O(N__42126),
            .I(N__42103));
    LocalMux I__9317 (
            .O(N__42123),
            .I(N__42096));
    Span4Mux_v I__9316 (
            .O(N__42120),
            .I(N__42096));
    LocalMux I__9315 (
            .O(N__42117),
            .I(N__42096));
    Span4Mux_h I__9314 (
            .O(N__42112),
            .I(N__42093));
    Span4Mux_h I__9313 (
            .O(N__42109),
            .I(N__42090));
    LocalMux I__9312 (
            .O(N__42106),
            .I(N__42087));
    Span4Mux_h I__9311 (
            .O(N__42103),
            .I(N__42082));
    Span4Mux_v I__9310 (
            .O(N__42096),
            .I(N__42082));
    Span4Mux_v I__9309 (
            .O(N__42093),
            .I(N__42079));
    Span4Mux_h I__9308 (
            .O(N__42090),
            .I(N__42076));
    Span12Mux_h I__9307 (
            .O(N__42087),
            .I(N__42073));
    Span4Mux_h I__9306 (
            .O(N__42082),
            .I(N__42070));
    Odrv4 I__9305 (
            .O(N__42079),
            .I(\ALU.r0_12_1_THRU_CO ));
    Odrv4 I__9304 (
            .O(N__42076),
            .I(\ALU.r0_12_1_THRU_CO ));
    Odrv12 I__9303 (
            .O(N__42073),
            .I(\ALU.r0_12_1_THRU_CO ));
    Odrv4 I__9302 (
            .O(N__42070),
            .I(\ALU.r0_12_1_THRU_CO ));
    CascadeMux I__9301 (
            .O(N__42061),
            .I(N__42058));
    InMux I__9300 (
            .O(N__42058),
            .I(N__42052));
    InMux I__9299 (
            .O(N__42057),
            .I(N__42052));
    LocalMux I__9298 (
            .O(N__42052),
            .I(N__42049));
    Span4Mux_v I__9297 (
            .O(N__42049),
            .I(N__42046));
    Odrv4 I__9296 (
            .O(N__42046),
            .I(\ALU.un9_addsub_cry_0_c_RNIG8GLJZ0 ));
    InMux I__9295 (
            .O(N__42043),
            .I(N__42040));
    LocalMux I__9294 (
            .O(N__42040),
            .I(\ALU.r0_12_prm_1_1_c_RNOZ0 ));
    CascadeMux I__9293 (
            .O(N__42037),
            .I(N__42034));
    InMux I__9292 (
            .O(N__42034),
            .I(N__42031));
    LocalMux I__9291 (
            .O(N__42031),
            .I(N__42028));
    Odrv12 I__9290 (
            .O(N__42028),
            .I(\ALU.r0_12_prm_5_9_s0_c_RNOZ0 ));
    CascadeMux I__9289 (
            .O(N__42025),
            .I(N__42022));
    InMux I__9288 (
            .O(N__42022),
            .I(N__42018));
    InMux I__9287 (
            .O(N__42021),
            .I(N__42015));
    LocalMux I__9286 (
            .O(N__42018),
            .I(N__42012));
    LocalMux I__9285 (
            .O(N__42015),
            .I(\ALU.r4_RNIKUMQ8_0Z0Z_8 ));
    Odrv12 I__9284 (
            .O(N__42012),
            .I(\ALU.r4_RNIKUMQ8_0Z0Z_8 ));
    CascadeMux I__9283 (
            .O(N__42007),
            .I(N__42004));
    InMux I__9282 (
            .O(N__42004),
            .I(N__42001));
    LocalMux I__9281 (
            .O(N__42001),
            .I(\ALU.r0_12_prm_6_8_s1_c_RNOZ0 ));
    CascadeMux I__9280 (
            .O(N__41998),
            .I(N__41995));
    InMux I__9279 (
            .O(N__41995),
            .I(N__41992));
    LocalMux I__9278 (
            .O(N__41992),
            .I(N__41989));
    Span12Mux_s9_h I__9277 (
            .O(N__41989),
            .I(N__41986));
    Odrv12 I__9276 (
            .O(N__41986),
            .I(\ALU.r0_12_prm_8_10_s0_c_RNOZ0 ));
    CascadeMux I__9275 (
            .O(N__41983),
            .I(N__41980));
    InMux I__9274 (
            .O(N__41980),
            .I(N__41976));
    InMux I__9273 (
            .O(N__41979),
            .I(N__41973));
    LocalMux I__9272 (
            .O(N__41976),
            .I(\ALU.rshift_1 ));
    LocalMux I__9271 (
            .O(N__41973),
            .I(\ALU.rshift_1 ));
    CascadeMux I__9270 (
            .O(N__41968),
            .I(N__41965));
    InMux I__9269 (
            .O(N__41965),
            .I(N__41962));
    LocalMux I__9268 (
            .O(N__41962),
            .I(N__41959));
    Odrv4 I__9267 (
            .O(N__41959),
            .I(\ALU.lshift_1 ));
    InMux I__9266 (
            .O(N__41956),
            .I(N__41953));
    LocalMux I__9265 (
            .O(N__41953),
            .I(N__41948));
    InMux I__9264 (
            .O(N__41952),
            .I(N__41943));
    InMux I__9263 (
            .O(N__41951),
            .I(N__41943));
    Span4Mux_v I__9262 (
            .O(N__41948),
            .I(N__41939));
    LocalMux I__9261 (
            .O(N__41943),
            .I(N__41936));
    InMux I__9260 (
            .O(N__41942),
            .I(N__41933));
    Span4Mux_h I__9259 (
            .O(N__41939),
            .I(N__41928));
    Span4Mux_h I__9258 (
            .O(N__41936),
            .I(N__41928));
    LocalMux I__9257 (
            .O(N__41933),
            .I(\ALU.a1_b_1 ));
    Odrv4 I__9256 (
            .O(N__41928),
            .I(\ALU.a1_b_1 ));
    CascadeMux I__9255 (
            .O(N__41923),
            .I(N__41920));
    InMux I__9254 (
            .O(N__41920),
            .I(N__41917));
    LocalMux I__9253 (
            .O(N__41917),
            .I(N__41914));
    Span4Mux_h I__9252 (
            .O(N__41914),
            .I(N__41911));
    Span4Mux_h I__9251 (
            .O(N__41911),
            .I(N__41908));
    Odrv4 I__9250 (
            .O(N__41908),
            .I(\ALU.r0_12_prm_7_1_c_RNOZ0 ));
    InMux I__9249 (
            .O(N__41905),
            .I(N__41902));
    LocalMux I__9248 (
            .O(N__41902),
            .I(N__41899));
    Span4Mux_v I__9247 (
            .O(N__41899),
            .I(N__41896));
    Odrv4 I__9246 (
            .O(N__41896),
            .I(\ALU.r0_12_prm_6_1_c_RNOZ0 ));
    InMux I__9245 (
            .O(N__41893),
            .I(N__41890));
    LocalMux I__9244 (
            .O(N__41890),
            .I(N__41887));
    Span4Mux_h I__9243 (
            .O(N__41887),
            .I(N__41884));
    Odrv4 I__9242 (
            .O(N__41884),
            .I(\ALU.r0_12_prm_5_1_c_RNOZ0 ));
    InMux I__9241 (
            .O(N__41881),
            .I(N__41878));
    LocalMux I__9240 (
            .O(N__41878),
            .I(N__41875));
    Span4Mux_v I__9239 (
            .O(N__41875),
            .I(N__41872));
    Odrv4 I__9238 (
            .O(N__41872),
            .I(\ALU.r4_RNID1636Z0Z_1 ));
    CascadeMux I__9237 (
            .O(N__41869),
            .I(N__41866));
    InMux I__9236 (
            .O(N__41866),
            .I(N__41863));
    LocalMux I__9235 (
            .O(N__41863),
            .I(\ALU.a_i_1 ));
    InMux I__9234 (
            .O(N__41860),
            .I(N__41857));
    LocalMux I__9233 (
            .O(N__41857),
            .I(N__41854));
    Span4Mux_v I__9232 (
            .O(N__41854),
            .I(N__41851));
    Sp12to4 I__9231 (
            .O(N__41851),
            .I(N__41848));
    Span12Mux_h I__9230 (
            .O(N__41848),
            .I(N__41845));
    Odrv12 I__9229 (
            .O(N__41845),
            .I(\ALU.r0_12_prm_3_1_c_RNOZ0 ));
    CascadeMux I__9228 (
            .O(N__41842),
            .I(N__41839));
    InMux I__9227 (
            .O(N__41839),
            .I(N__41836));
    LocalMux I__9226 (
            .O(N__41836),
            .I(N__41833));
    Span4Mux_v I__9225 (
            .O(N__41833),
            .I(N__41830));
    Span4Mux_h I__9224 (
            .O(N__41830),
            .I(N__41827));
    Span4Mux_h I__9223 (
            .O(N__41827),
            .I(N__41824));
    Span4Mux_h I__9222 (
            .O(N__41824),
            .I(N__41820));
    InMux I__9221 (
            .O(N__41823),
            .I(N__41817));
    Span4Mux_s1_h I__9220 (
            .O(N__41820),
            .I(N__41812));
    LocalMux I__9219 (
            .O(N__41817),
            .I(N__41812));
    Odrv4 I__9218 (
            .O(N__41812),
            .I(\ALU.mult_1 ));
    InMux I__9217 (
            .O(N__41809),
            .I(N__41806));
    LocalMux I__9216 (
            .O(N__41806),
            .I(\ALU.r4_RNIVFRGQ_0Z0Z_2 ));
    InMux I__9215 (
            .O(N__41803),
            .I(N__41800));
    LocalMux I__9214 (
            .O(N__41800),
            .I(\ALU.r0_12_prm_8_4_c_RNOZ0 ));
    InMux I__9213 (
            .O(N__41797),
            .I(N__41793));
    InMux I__9212 (
            .O(N__41796),
            .I(N__41790));
    LocalMux I__9211 (
            .O(N__41793),
            .I(N__41787));
    LocalMux I__9210 (
            .O(N__41790),
            .I(N__41784));
    Span4Mux_h I__9209 (
            .O(N__41787),
            .I(N__41781));
    Span4Mux_v I__9208 (
            .O(N__41784),
            .I(N__41778));
    Sp12to4 I__9207 (
            .O(N__41781),
            .I(N__41775));
    Odrv4 I__9206 (
            .O(N__41778),
            .I(\ALU.r4_RNIODO6KZ0Z_7 ));
    Odrv12 I__9205 (
            .O(N__41775),
            .I(\ALU.r4_RNIODO6KZ0Z_7 ));
    InMux I__9204 (
            .O(N__41770),
            .I(N__41767));
    LocalMux I__9203 (
            .O(N__41767),
            .I(N__41764));
    Odrv4 I__9202 (
            .O(N__41764),
            .I(\ALU.r0_12_prm_8_4_c_RNOZ0Z_3 ));
    InMux I__9201 (
            .O(N__41761),
            .I(N__41757));
    InMux I__9200 (
            .O(N__41760),
            .I(N__41754));
    LocalMux I__9199 (
            .O(N__41757),
            .I(N__41751));
    LocalMux I__9198 (
            .O(N__41754),
            .I(N__41748));
    Span4Mux_h I__9197 (
            .O(N__41751),
            .I(N__41745));
    Span4Mux_v I__9196 (
            .O(N__41748),
            .I(N__41742));
    Odrv4 I__9195 (
            .O(N__41745),
            .I(\ALU.un9_addsub_cry_3_c_RNIV8DFIZ0 ));
    Odrv4 I__9194 (
            .O(N__41742),
            .I(\ALU.un9_addsub_cry_3_c_RNIV8DFIZ0 ));
    CascadeMux I__9193 (
            .O(N__41737),
            .I(N__41734));
    InMux I__9192 (
            .O(N__41734),
            .I(N__41731));
    LocalMux I__9191 (
            .O(N__41731),
            .I(\ALU.r0_12_prm_1_4_c_RNOZ0 ));
    InMux I__9190 (
            .O(N__41728),
            .I(N__41723));
    InMux I__9189 (
            .O(N__41727),
            .I(N__41718));
    InMux I__9188 (
            .O(N__41726),
            .I(N__41718));
    LocalMux I__9187 (
            .O(N__41723),
            .I(N__41715));
    LocalMux I__9186 (
            .O(N__41718),
            .I(N__41712));
    Odrv4 I__9185 (
            .O(N__41715),
            .I(\ALU.r5_RNI7NOB9Z0Z_13 ));
    Odrv12 I__9184 (
            .O(N__41712),
            .I(\ALU.r5_RNI7NOB9Z0Z_13 ));
    InMux I__9183 (
            .O(N__41707),
            .I(N__41703));
    InMux I__9182 (
            .O(N__41706),
            .I(N__41700));
    LocalMux I__9181 (
            .O(N__41703),
            .I(N__41697));
    LocalMux I__9180 (
            .O(N__41700),
            .I(N__41694));
    Span4Mux_s2_v I__9179 (
            .O(N__41697),
            .I(N__41691));
    Span4Mux_h I__9178 (
            .O(N__41694),
            .I(N__41688));
    Span4Mux_h I__9177 (
            .O(N__41691),
            .I(N__41682));
    Span4Mux_v I__9176 (
            .O(N__41688),
            .I(N__41679));
    InMux I__9175 (
            .O(N__41687),
            .I(N__41674));
    InMux I__9174 (
            .O(N__41686),
            .I(N__41674));
    InMux I__9173 (
            .O(N__41685),
            .I(N__41671));
    Odrv4 I__9172 (
            .O(N__41682),
            .I(\ALU.r5_RNIUE7TIZ0Z_13 ));
    Odrv4 I__9171 (
            .O(N__41679),
            .I(\ALU.r5_RNIUE7TIZ0Z_13 ));
    LocalMux I__9170 (
            .O(N__41674),
            .I(\ALU.r5_RNIUE7TIZ0Z_13 ));
    LocalMux I__9169 (
            .O(N__41671),
            .I(\ALU.r5_RNIUE7TIZ0Z_13 ));
    InMux I__9168 (
            .O(N__41662),
            .I(N__41658));
    InMux I__9167 (
            .O(N__41661),
            .I(N__41655));
    LocalMux I__9166 (
            .O(N__41658),
            .I(\ALU.r4_RNIRL1V71Z0Z_7 ));
    LocalMux I__9165 (
            .O(N__41655),
            .I(\ALU.r4_RNIRL1V71Z0Z_7 ));
    InMux I__9164 (
            .O(N__41650),
            .I(N__41646));
    InMux I__9163 (
            .O(N__41649),
            .I(N__41643));
    LocalMux I__9162 (
            .O(N__41646),
            .I(N__41639));
    LocalMux I__9161 (
            .O(N__41643),
            .I(N__41636));
    InMux I__9160 (
            .O(N__41642),
            .I(N__41633));
    Span4Mux_v I__9159 (
            .O(N__41639),
            .I(N__41630));
    Span4Mux_h I__9158 (
            .O(N__41636),
            .I(N__41626));
    LocalMux I__9157 (
            .O(N__41633),
            .I(N__41623));
    Span4Mux_h I__9156 (
            .O(N__41630),
            .I(N__41620));
    InMux I__9155 (
            .O(N__41629),
            .I(N__41617));
    Span4Mux_h I__9154 (
            .O(N__41626),
            .I(N__41614));
    Span4Mux_h I__9153 (
            .O(N__41623),
            .I(N__41607));
    Span4Mux_v I__9152 (
            .O(N__41620),
            .I(N__41607));
    LocalMux I__9151 (
            .O(N__41617),
            .I(N__41607));
    Odrv4 I__9150 (
            .O(N__41614),
            .I(\ALU.a6_b_6 ));
    Odrv4 I__9149 (
            .O(N__41607),
            .I(\ALU.a6_b_6 ));
    CascadeMux I__9148 (
            .O(N__41602),
            .I(N__41599));
    InMux I__9147 (
            .O(N__41599),
            .I(N__41596));
    LocalMux I__9146 (
            .O(N__41596),
            .I(N__41593));
    Span4Mux_s2_v I__9145 (
            .O(N__41593),
            .I(N__41590));
    Odrv4 I__9144 (
            .O(N__41590),
            .I(\ALU.r0_12_prm_7_6_s0_c_RNOZ0 ));
    CascadeMux I__9143 (
            .O(N__41587),
            .I(N__41584));
    InMux I__9142 (
            .O(N__41584),
            .I(N__41581));
    LocalMux I__9141 (
            .O(N__41581),
            .I(N__41578));
    Span12Mux_s4_v I__9140 (
            .O(N__41578),
            .I(N__41575));
    Odrv12 I__9139 (
            .O(N__41575),
            .I(\ALU.r0_12_prm_6_6_s0_c_RNOZ0 ));
    InMux I__9138 (
            .O(N__41572),
            .I(N__41567));
    InMux I__9137 (
            .O(N__41571),
            .I(N__41562));
    InMux I__9136 (
            .O(N__41570),
            .I(N__41558));
    LocalMux I__9135 (
            .O(N__41567),
            .I(N__41552));
    InMux I__9134 (
            .O(N__41566),
            .I(N__41549));
    CascadeMux I__9133 (
            .O(N__41565),
            .I(N__41545));
    LocalMux I__9132 (
            .O(N__41562),
            .I(N__41539));
    InMux I__9131 (
            .O(N__41561),
            .I(N__41536));
    LocalMux I__9130 (
            .O(N__41558),
            .I(N__41533));
    InMux I__9129 (
            .O(N__41557),
            .I(N__41530));
    InMux I__9128 (
            .O(N__41556),
            .I(N__41527));
    InMux I__9127 (
            .O(N__41555),
            .I(N__41524));
    Span4Mux_v I__9126 (
            .O(N__41552),
            .I(N__41521));
    LocalMux I__9125 (
            .O(N__41549),
            .I(N__41517));
    InMux I__9124 (
            .O(N__41548),
            .I(N__41512));
    InMux I__9123 (
            .O(N__41545),
            .I(N__41512));
    InMux I__9122 (
            .O(N__41544),
            .I(N__41505));
    InMux I__9121 (
            .O(N__41543),
            .I(N__41505));
    InMux I__9120 (
            .O(N__41542),
            .I(N__41505));
    Span4Mux_h I__9119 (
            .O(N__41539),
            .I(N__41493));
    LocalMux I__9118 (
            .O(N__41536),
            .I(N__41493));
    Span4Mux_v I__9117 (
            .O(N__41533),
            .I(N__41490));
    LocalMux I__9116 (
            .O(N__41530),
            .I(N__41485));
    LocalMux I__9115 (
            .O(N__41527),
            .I(N__41485));
    LocalMux I__9114 (
            .O(N__41524),
            .I(N__41482));
    Span4Mux_v I__9113 (
            .O(N__41521),
            .I(N__41479));
    InMux I__9112 (
            .O(N__41520),
            .I(N__41475));
    Span4Mux_h I__9111 (
            .O(N__41517),
            .I(N__41472));
    LocalMux I__9110 (
            .O(N__41512),
            .I(N__41469));
    LocalMux I__9109 (
            .O(N__41505),
            .I(N__41465));
    InMux I__9108 (
            .O(N__41504),
            .I(N__41449));
    InMux I__9107 (
            .O(N__41503),
            .I(N__41449));
    InMux I__9106 (
            .O(N__41502),
            .I(N__41449));
    InMux I__9105 (
            .O(N__41501),
            .I(N__41449));
    InMux I__9104 (
            .O(N__41500),
            .I(N__41449));
    InMux I__9103 (
            .O(N__41499),
            .I(N__41449));
    InMux I__9102 (
            .O(N__41498),
            .I(N__41449));
    Span4Mux_v I__9101 (
            .O(N__41493),
            .I(N__41446));
    Span4Mux_v I__9100 (
            .O(N__41490),
            .I(N__41442));
    Span4Mux_v I__9099 (
            .O(N__41485),
            .I(N__41437));
    Span4Mux_h I__9098 (
            .O(N__41482),
            .I(N__41437));
    Span4Mux_v I__9097 (
            .O(N__41479),
            .I(N__41434));
    InMux I__9096 (
            .O(N__41478),
            .I(N__41431));
    LocalMux I__9095 (
            .O(N__41475),
            .I(N__41428));
    Span4Mux_v I__9094 (
            .O(N__41472),
            .I(N__41425));
    Span4Mux_v I__9093 (
            .O(N__41469),
            .I(N__41422));
    InMux I__9092 (
            .O(N__41468),
            .I(N__41419));
    Span4Mux_v I__9091 (
            .O(N__41465),
            .I(N__41416));
    InMux I__9090 (
            .O(N__41464),
            .I(N__41413));
    LocalMux I__9089 (
            .O(N__41449),
            .I(N__41408));
    Span4Mux_h I__9088 (
            .O(N__41446),
            .I(N__41408));
    InMux I__9087 (
            .O(N__41445),
            .I(N__41405));
    Span4Mux_h I__9086 (
            .O(N__41442),
            .I(N__41400));
    Span4Mux_h I__9085 (
            .O(N__41437),
            .I(N__41400));
    Sp12to4 I__9084 (
            .O(N__41434),
            .I(N__41395));
    LocalMux I__9083 (
            .O(N__41431),
            .I(N__41395));
    Span4Mux_h I__9082 (
            .O(N__41428),
            .I(N__41390));
    Span4Mux_v I__9081 (
            .O(N__41425),
            .I(N__41390));
    Span4Mux_v I__9080 (
            .O(N__41422),
            .I(N__41387));
    LocalMux I__9079 (
            .O(N__41419),
            .I(\ALU.a_13 ));
    Odrv4 I__9078 (
            .O(N__41416),
            .I(\ALU.a_13 ));
    LocalMux I__9077 (
            .O(N__41413),
            .I(\ALU.a_13 ));
    Odrv4 I__9076 (
            .O(N__41408),
            .I(\ALU.a_13 ));
    LocalMux I__9075 (
            .O(N__41405),
            .I(\ALU.a_13 ));
    Odrv4 I__9074 (
            .O(N__41400),
            .I(\ALU.a_13 ));
    Odrv12 I__9073 (
            .O(N__41395),
            .I(\ALU.a_13 ));
    Odrv4 I__9072 (
            .O(N__41390),
            .I(\ALU.a_13 ));
    Odrv4 I__9071 (
            .O(N__41387),
            .I(\ALU.a_13 ));
    CascadeMux I__9070 (
            .O(N__41368),
            .I(N__41359));
    InMux I__9069 (
            .O(N__41367),
            .I(N__41346));
    InMux I__9068 (
            .O(N__41366),
            .I(N__41343));
    CascadeMux I__9067 (
            .O(N__41365),
            .I(N__41340));
    CascadeMux I__9066 (
            .O(N__41364),
            .I(N__41336));
    CascadeMux I__9065 (
            .O(N__41363),
            .I(N__41333));
    CascadeMux I__9064 (
            .O(N__41362),
            .I(N__41330));
    InMux I__9063 (
            .O(N__41359),
            .I(N__41324));
    InMux I__9062 (
            .O(N__41358),
            .I(N__41324));
    InMux I__9061 (
            .O(N__41357),
            .I(N__41321));
    InMux I__9060 (
            .O(N__41356),
            .I(N__41318));
    InMux I__9059 (
            .O(N__41355),
            .I(N__41311));
    InMux I__9058 (
            .O(N__41354),
            .I(N__41306));
    InMux I__9057 (
            .O(N__41353),
            .I(N__41306));
    InMux I__9056 (
            .O(N__41352),
            .I(N__41303));
    InMux I__9055 (
            .O(N__41351),
            .I(N__41298));
    InMux I__9054 (
            .O(N__41350),
            .I(N__41295));
    InMux I__9053 (
            .O(N__41349),
            .I(N__41290));
    LocalMux I__9052 (
            .O(N__41346),
            .I(N__41285));
    LocalMux I__9051 (
            .O(N__41343),
            .I(N__41285));
    InMux I__9050 (
            .O(N__41340),
            .I(N__41282));
    InMux I__9049 (
            .O(N__41339),
            .I(N__41277));
    InMux I__9048 (
            .O(N__41336),
            .I(N__41277));
    InMux I__9047 (
            .O(N__41333),
            .I(N__41271));
    InMux I__9046 (
            .O(N__41330),
            .I(N__41271));
    InMux I__9045 (
            .O(N__41329),
            .I(N__41268));
    LocalMux I__9044 (
            .O(N__41324),
            .I(N__41265));
    LocalMux I__9043 (
            .O(N__41321),
            .I(N__41262));
    LocalMux I__9042 (
            .O(N__41318),
            .I(N__41259));
    InMux I__9041 (
            .O(N__41317),
            .I(N__41256));
    InMux I__9040 (
            .O(N__41316),
            .I(N__41253));
    InMux I__9039 (
            .O(N__41315),
            .I(N__41248));
    InMux I__9038 (
            .O(N__41314),
            .I(N__41248));
    LocalMux I__9037 (
            .O(N__41311),
            .I(N__41243));
    LocalMux I__9036 (
            .O(N__41306),
            .I(N__41243));
    LocalMux I__9035 (
            .O(N__41303),
            .I(N__41240));
    InMux I__9034 (
            .O(N__41302),
            .I(N__41235));
    InMux I__9033 (
            .O(N__41301),
            .I(N__41235));
    LocalMux I__9032 (
            .O(N__41298),
            .I(N__41232));
    LocalMux I__9031 (
            .O(N__41295),
            .I(N__41229));
    InMux I__9030 (
            .O(N__41294),
            .I(N__41224));
    InMux I__9029 (
            .O(N__41293),
            .I(N__41224));
    LocalMux I__9028 (
            .O(N__41290),
            .I(N__41221));
    Span4Mux_v I__9027 (
            .O(N__41285),
            .I(N__41218));
    LocalMux I__9026 (
            .O(N__41282),
            .I(N__41213));
    LocalMux I__9025 (
            .O(N__41277),
            .I(N__41213));
    InMux I__9024 (
            .O(N__41276),
            .I(N__41210));
    LocalMux I__9023 (
            .O(N__41271),
            .I(N__41207));
    LocalMux I__9022 (
            .O(N__41268),
            .I(N__41204));
    Span4Mux_v I__9021 (
            .O(N__41265),
            .I(N__41199));
    Span4Mux_h I__9020 (
            .O(N__41262),
            .I(N__41199));
    Span4Mux_h I__9019 (
            .O(N__41259),
            .I(N__41196));
    LocalMux I__9018 (
            .O(N__41256),
            .I(N__41193));
    LocalMux I__9017 (
            .O(N__41253),
            .I(N__41190));
    LocalMux I__9016 (
            .O(N__41248),
            .I(N__41187));
    Span4Mux_v I__9015 (
            .O(N__41243),
            .I(N__41180));
    Span4Mux_v I__9014 (
            .O(N__41240),
            .I(N__41180));
    LocalMux I__9013 (
            .O(N__41235),
            .I(N__41180));
    Span4Mux_h I__9012 (
            .O(N__41232),
            .I(N__41173));
    Span4Mux_h I__9011 (
            .O(N__41229),
            .I(N__41173));
    LocalMux I__9010 (
            .O(N__41224),
            .I(N__41173));
    Span4Mux_v I__9009 (
            .O(N__41221),
            .I(N__41170));
    Span4Mux_h I__9008 (
            .O(N__41218),
            .I(N__41167));
    Span4Mux_v I__9007 (
            .O(N__41213),
            .I(N__41162));
    LocalMux I__9006 (
            .O(N__41210),
            .I(N__41162));
    Span4Mux_h I__9005 (
            .O(N__41207),
            .I(N__41155));
    Span4Mux_v I__9004 (
            .O(N__41204),
            .I(N__41155));
    Span4Mux_h I__9003 (
            .O(N__41199),
            .I(N__41155));
    Span4Mux_h I__9002 (
            .O(N__41196),
            .I(N__41150));
    Span4Mux_h I__9001 (
            .O(N__41193),
            .I(N__41150));
    Span4Mux_v I__9000 (
            .O(N__41190),
            .I(N__41145));
    Span4Mux_v I__8999 (
            .O(N__41187),
            .I(N__41145));
    Span4Mux_h I__8998 (
            .O(N__41180),
            .I(N__41140));
    Span4Mux_v I__8997 (
            .O(N__41173),
            .I(N__41140));
    Span4Mux_h I__8996 (
            .O(N__41170),
            .I(N__41135));
    Span4Mux_h I__8995 (
            .O(N__41167),
            .I(N__41135));
    Span4Mux_h I__8994 (
            .O(N__41162),
            .I(N__41132));
    Odrv4 I__8993 (
            .O(N__41155),
            .I(\ALU.a_12 ));
    Odrv4 I__8992 (
            .O(N__41150),
            .I(\ALU.a_12 ));
    Odrv4 I__8991 (
            .O(N__41145),
            .I(\ALU.a_12 ));
    Odrv4 I__8990 (
            .O(N__41140),
            .I(\ALU.a_12 ));
    Odrv4 I__8989 (
            .O(N__41135),
            .I(\ALU.a_12 ));
    Odrv4 I__8988 (
            .O(N__41132),
            .I(\ALU.a_12 ));
    InMux I__8987 (
            .O(N__41119),
            .I(N__41115));
    InMux I__8986 (
            .O(N__41118),
            .I(N__41112));
    LocalMux I__8985 (
            .O(N__41115),
            .I(N__41109));
    LocalMux I__8984 (
            .O(N__41112),
            .I(N__41104));
    Span4Mux_h I__8983 (
            .O(N__41109),
            .I(N__41104));
    Span4Mux_v I__8982 (
            .O(N__41104),
            .I(N__41101));
    Odrv4 I__8981 (
            .O(N__41101),
            .I(\ALU.r4_RNI9H7SJZ0Z_6 ));
    InMux I__8980 (
            .O(N__41098),
            .I(N__41095));
    LocalMux I__8979 (
            .O(N__41095),
            .I(N__41092));
    Span4Mux_h I__8978 (
            .O(N__41092),
            .I(N__41087));
    InMux I__8977 (
            .O(N__41091),
            .I(N__41084));
    InMux I__8976 (
            .O(N__41090),
            .I(N__41081));
    Odrv4 I__8975 (
            .O(N__41087),
            .I(\ALU.r5_RNI0QK3KZ0Z_11 ));
    LocalMux I__8974 (
            .O(N__41084),
            .I(\ALU.r5_RNI0QK3KZ0Z_11 ));
    LocalMux I__8973 (
            .O(N__41081),
            .I(\ALU.r5_RNI0QK3KZ0Z_11 ));
    CascadeMux I__8972 (
            .O(N__41074),
            .I(\ALU.r0_12_prm_8_4_c_RNOZ0Z_2_cascade_ ));
    CascadeMux I__8971 (
            .O(N__41071),
            .I(N__41068));
    InMux I__8970 (
            .O(N__41068),
            .I(N__41064));
    InMux I__8969 (
            .O(N__41067),
            .I(N__41061));
    LocalMux I__8968 (
            .O(N__41064),
            .I(\ALU.rshift_4 ));
    LocalMux I__8967 (
            .O(N__41061),
            .I(\ALU.rshift_4 ));
    InMux I__8966 (
            .O(N__41056),
            .I(N__41053));
    LocalMux I__8965 (
            .O(N__41053),
            .I(\ALU.lshift_15_ns_1_8 ));
    InMux I__8964 (
            .O(N__41050),
            .I(N__41047));
    LocalMux I__8963 (
            .O(N__41047),
            .I(\ALU.lshift_3_ns_1_4 ));
    InMux I__8962 (
            .O(N__41044),
            .I(N__41040));
    InMux I__8961 (
            .O(N__41043),
            .I(N__41037));
    LocalMux I__8960 (
            .O(N__41040),
            .I(\ALU.r4_RNI6PL1LZ0Z_2 ));
    LocalMux I__8959 (
            .O(N__41037),
            .I(\ALU.r4_RNI6PL1LZ0Z_2 ));
    CascadeMux I__8958 (
            .O(N__41032),
            .I(\ALU.r4_RNI6PL1LZ0Z_2_cascade_ ));
    InMux I__8957 (
            .O(N__41029),
            .I(N__41026));
    LocalMux I__8956 (
            .O(N__41026),
            .I(N__41021));
    InMux I__8955 (
            .O(N__41025),
            .I(N__41018));
    InMux I__8954 (
            .O(N__41024),
            .I(N__41015));
    Span4Mux_v I__8953 (
            .O(N__41021),
            .I(N__41008));
    LocalMux I__8952 (
            .O(N__41018),
            .I(N__41008));
    LocalMux I__8951 (
            .O(N__41015),
            .I(N__41008));
    Span4Mux_h I__8950 (
            .O(N__41008),
            .I(N__41005));
    Span4Mux_v I__8949 (
            .O(N__41005),
            .I(N__41002));
    Odrv4 I__8948 (
            .O(N__41002),
            .I(\ALU.r4_RNIVFRGQZ0Z_2 ));
    CascadeMux I__8947 (
            .O(N__40999),
            .I(\ALU.rshift_3_ns_1_9_cascade_ ));
    InMux I__8946 (
            .O(N__40996),
            .I(N__40993));
    LocalMux I__8945 (
            .O(N__40993),
            .I(N__40983));
    InMux I__8944 (
            .O(N__40992),
            .I(N__40974));
    InMux I__8943 (
            .O(N__40991),
            .I(N__40974));
    InMux I__8942 (
            .O(N__40990),
            .I(N__40974));
    CascadeMux I__8941 (
            .O(N__40989),
            .I(N__40971));
    InMux I__8940 (
            .O(N__40988),
            .I(N__40951));
    InMux I__8939 (
            .O(N__40987),
            .I(N__40951));
    InMux I__8938 (
            .O(N__40986),
            .I(N__40948));
    Span4Mux_v I__8937 (
            .O(N__40983),
            .I(N__40945));
    InMux I__8936 (
            .O(N__40982),
            .I(N__40942));
    InMux I__8935 (
            .O(N__40981),
            .I(N__40939));
    LocalMux I__8934 (
            .O(N__40974),
            .I(N__40936));
    InMux I__8933 (
            .O(N__40971),
            .I(N__40933));
    CascadeMux I__8932 (
            .O(N__40970),
            .I(N__40928));
    InMux I__8931 (
            .O(N__40969),
            .I(N__40925));
    InMux I__8930 (
            .O(N__40968),
            .I(N__40912));
    InMux I__8929 (
            .O(N__40967),
            .I(N__40912));
    InMux I__8928 (
            .O(N__40966),
            .I(N__40912));
    InMux I__8927 (
            .O(N__40965),
            .I(N__40912));
    InMux I__8926 (
            .O(N__40964),
            .I(N__40912));
    InMux I__8925 (
            .O(N__40963),
            .I(N__40912));
    InMux I__8924 (
            .O(N__40962),
            .I(N__40908));
    InMux I__8923 (
            .O(N__40961),
            .I(N__40901));
    InMux I__8922 (
            .O(N__40960),
            .I(N__40901));
    InMux I__8921 (
            .O(N__40959),
            .I(N__40901));
    InMux I__8920 (
            .O(N__40958),
            .I(N__40898));
    InMux I__8919 (
            .O(N__40957),
            .I(N__40893));
    InMux I__8918 (
            .O(N__40956),
            .I(N__40893));
    LocalMux I__8917 (
            .O(N__40951),
            .I(N__40889));
    LocalMux I__8916 (
            .O(N__40948),
            .I(N__40886));
    Span4Mux_v I__8915 (
            .O(N__40945),
            .I(N__40883));
    LocalMux I__8914 (
            .O(N__40942),
            .I(N__40878));
    LocalMux I__8913 (
            .O(N__40939),
            .I(N__40878));
    Span4Mux_v I__8912 (
            .O(N__40936),
            .I(N__40871));
    LocalMux I__8911 (
            .O(N__40933),
            .I(N__40871));
    InMux I__8910 (
            .O(N__40932),
            .I(N__40868));
    InMux I__8909 (
            .O(N__40931),
            .I(N__40865));
    InMux I__8908 (
            .O(N__40928),
            .I(N__40862));
    LocalMux I__8907 (
            .O(N__40925),
            .I(N__40857));
    LocalMux I__8906 (
            .O(N__40912),
            .I(N__40857));
    InMux I__8905 (
            .O(N__40911),
            .I(N__40854));
    LocalMux I__8904 (
            .O(N__40908),
            .I(N__40851));
    LocalMux I__8903 (
            .O(N__40901),
            .I(N__40846));
    LocalMux I__8902 (
            .O(N__40898),
            .I(N__40846));
    LocalMux I__8901 (
            .O(N__40893),
            .I(N__40843));
    InMux I__8900 (
            .O(N__40892),
            .I(N__40840));
    Span4Mux_s1_h I__8899 (
            .O(N__40889),
            .I(N__40837));
    Span4Mux_h I__8898 (
            .O(N__40886),
            .I(N__40834));
    Span4Mux_h I__8897 (
            .O(N__40883),
            .I(N__40829));
    Span4Mux_v I__8896 (
            .O(N__40878),
            .I(N__40829));
    InMux I__8895 (
            .O(N__40877),
            .I(N__40824));
    InMux I__8894 (
            .O(N__40876),
            .I(N__40824));
    Span4Mux_h I__8893 (
            .O(N__40871),
            .I(N__40817));
    LocalMux I__8892 (
            .O(N__40868),
            .I(N__40817));
    LocalMux I__8891 (
            .O(N__40865),
            .I(N__40817));
    LocalMux I__8890 (
            .O(N__40862),
            .I(N__40814));
    Span4Mux_v I__8889 (
            .O(N__40857),
            .I(N__40811));
    LocalMux I__8888 (
            .O(N__40854),
            .I(N__40806));
    Span12Mux_v I__8887 (
            .O(N__40851),
            .I(N__40806));
    Span4Mux_v I__8886 (
            .O(N__40846),
            .I(N__40793));
    Span4Mux_v I__8885 (
            .O(N__40843),
            .I(N__40793));
    LocalMux I__8884 (
            .O(N__40840),
            .I(N__40793));
    Span4Mux_v I__8883 (
            .O(N__40837),
            .I(N__40793));
    Span4Mux_v I__8882 (
            .O(N__40834),
            .I(N__40793));
    Span4Mux_h I__8881 (
            .O(N__40829),
            .I(N__40793));
    LocalMux I__8880 (
            .O(N__40824),
            .I(N__40788));
    Span4Mux_h I__8879 (
            .O(N__40817),
            .I(N__40788));
    Span4Mux_v I__8878 (
            .O(N__40814),
            .I(N__40785));
    Odrv4 I__8877 (
            .O(N__40811),
            .I(\ALU.a_11 ));
    Odrv12 I__8876 (
            .O(N__40806),
            .I(\ALU.a_11 ));
    Odrv4 I__8875 (
            .O(N__40793),
            .I(\ALU.a_11 ));
    Odrv4 I__8874 (
            .O(N__40788),
            .I(\ALU.a_11 ));
    Odrv4 I__8873 (
            .O(N__40785),
            .I(\ALU.a_11 ));
    InMux I__8872 (
            .O(N__40774),
            .I(N__40771));
    LocalMux I__8871 (
            .O(N__40771),
            .I(N__40768));
    Span12Mux_v I__8870 (
            .O(N__40768),
            .I(N__40765));
    Odrv12 I__8869 (
            .O(N__40765),
            .I(\ALU.r0_12_prm_5_8_s0_c_RNOZ0 ));
    CascadeMux I__8868 (
            .O(N__40762),
            .I(\ALU.N_610_1_cascade_ ));
    CascadeMux I__8867 (
            .O(N__40759),
            .I(\ALU.r4_RNIVFRGQ_0Z0Z_2_cascade_ ));
    CascadeMux I__8866 (
            .O(N__40756),
            .I(N__40753));
    InMux I__8865 (
            .O(N__40753),
            .I(N__40750));
    LocalMux I__8864 (
            .O(N__40750),
            .I(\ALU.lshift_4 ));
    InMux I__8863 (
            .O(N__40747),
            .I(N__40743));
    InMux I__8862 (
            .O(N__40746),
            .I(N__40740));
    LocalMux I__8861 (
            .O(N__40743),
            .I(N__40737));
    LocalMux I__8860 (
            .O(N__40740),
            .I(N__40732));
    Span4Mux_v I__8859 (
            .O(N__40737),
            .I(N__40732));
    Span4Mux_h I__8858 (
            .O(N__40732),
            .I(N__40727));
    InMux I__8857 (
            .O(N__40731),
            .I(N__40722));
    InMux I__8856 (
            .O(N__40730),
            .I(N__40722));
    Span4Mux_h I__8855 (
            .O(N__40727),
            .I(N__40717));
    LocalMux I__8854 (
            .O(N__40722),
            .I(N__40717));
    Odrv4 I__8853 (
            .O(N__40717),
            .I(\ALU.a2_b_2 ));
    CascadeMux I__8852 (
            .O(N__40714),
            .I(N__40711));
    InMux I__8851 (
            .O(N__40711),
            .I(N__40708));
    LocalMux I__8850 (
            .O(N__40708),
            .I(\ALU.r0_12_prm_7_2_c_RNOZ0 ));
    CascadeMux I__8849 (
            .O(N__40705),
            .I(N__40701));
    InMux I__8848 (
            .O(N__40704),
            .I(N__40698));
    InMux I__8847 (
            .O(N__40701),
            .I(N__40695));
    LocalMux I__8846 (
            .O(N__40698),
            .I(N__40691));
    LocalMux I__8845 (
            .O(N__40695),
            .I(N__40688));
    InMux I__8844 (
            .O(N__40694),
            .I(N__40684));
    Span4Mux_h I__8843 (
            .O(N__40691),
            .I(N__40679));
    Span4Mux_s2_v I__8842 (
            .O(N__40688),
            .I(N__40679));
    InMux I__8841 (
            .O(N__40687),
            .I(N__40676));
    LocalMux I__8840 (
            .O(N__40684),
            .I(N__40673));
    Odrv4 I__8839 (
            .O(N__40679),
            .I(\ALU.lshift_0 ));
    LocalMux I__8838 (
            .O(N__40676),
            .I(\ALU.lshift_0 ));
    Odrv4 I__8837 (
            .O(N__40673),
            .I(\ALU.lshift_0 ));
    CascadeMux I__8836 (
            .O(N__40666),
            .I(N__40663));
    InMux I__8835 (
            .O(N__40663),
            .I(N__40660));
    LocalMux I__8834 (
            .O(N__40660),
            .I(N__40657));
    Span4Mux_h I__8833 (
            .O(N__40657),
            .I(N__40654));
    Span4Mux_v I__8832 (
            .O(N__40654),
            .I(N__40651));
    Odrv4 I__8831 (
            .O(N__40651),
            .I(\ALU.r4_RNIHENK8_1Z0Z_7 ));
    InMux I__8830 (
            .O(N__40648),
            .I(N__40644));
    CascadeMux I__8829 (
            .O(N__40647),
            .I(N__40641));
    LocalMux I__8828 (
            .O(N__40644),
            .I(N__40638));
    InMux I__8827 (
            .O(N__40641),
            .I(N__40635));
    Span4Mux_v I__8826 (
            .O(N__40638),
            .I(N__40632));
    LocalMux I__8825 (
            .O(N__40635),
            .I(N__40629));
    Span4Mux_h I__8824 (
            .O(N__40632),
            .I(N__40624));
    Span4Mux_h I__8823 (
            .O(N__40629),
            .I(N__40624));
    Span4Mux_v I__8822 (
            .O(N__40624),
            .I(N__40621));
    Odrv4 I__8821 (
            .O(N__40621),
            .I(\ALU.b_i_0 ));
    CascadeMux I__8820 (
            .O(N__40618),
            .I(N__40614));
    InMux I__8819 (
            .O(N__40617),
            .I(N__40611));
    InMux I__8818 (
            .O(N__40614),
            .I(N__40608));
    LocalMux I__8817 (
            .O(N__40611),
            .I(N__40603));
    LocalMux I__8816 (
            .O(N__40608),
            .I(N__40600));
    InMux I__8815 (
            .O(N__40607),
            .I(N__40597));
    InMux I__8814 (
            .O(N__40606),
            .I(N__40594));
    Span4Mux_s2_v I__8813 (
            .O(N__40603),
            .I(N__40587));
    Span4Mux_s2_v I__8812 (
            .O(N__40600),
            .I(N__40587));
    LocalMux I__8811 (
            .O(N__40597),
            .I(N__40587));
    LocalMux I__8810 (
            .O(N__40594),
            .I(N__40584));
    Odrv4 I__8809 (
            .O(N__40587),
            .I(\ALU.un2_addsub_axb_0_i ));
    Odrv4 I__8808 (
            .O(N__40584),
            .I(\ALU.un2_addsub_axb_0_i ));
    CascadeMux I__8807 (
            .O(N__40579),
            .I(N__40576));
    InMux I__8806 (
            .O(N__40576),
            .I(N__40573));
    LocalMux I__8805 (
            .O(N__40573),
            .I(N__40569));
    InMux I__8804 (
            .O(N__40572),
            .I(N__40566));
    Span4Mux_s1_v I__8803 (
            .O(N__40569),
            .I(N__40561));
    LocalMux I__8802 (
            .O(N__40566),
            .I(N__40561));
    Span4Mux_v I__8801 (
            .O(N__40561),
            .I(N__40558));
    Span4Mux_h I__8800 (
            .O(N__40558),
            .I(N__40555));
    Odrv4 I__8799 (
            .O(N__40555),
            .I(\ALU.un2_addsub_cry_1_c_RNI1H7SGZ0 ));
    InMux I__8798 (
            .O(N__40552),
            .I(N__40549));
    LocalMux I__8797 (
            .O(N__40549),
            .I(N__40546));
    Odrv4 I__8796 (
            .O(N__40546),
            .I(\ALU.r0_12_prm_2_2_c_RNOZ0 ));
    InMux I__8795 (
            .O(N__40543),
            .I(N__40540));
    LocalMux I__8794 (
            .O(N__40540),
            .I(N__40537));
    Odrv4 I__8793 (
            .O(N__40537),
            .I(\ALU.r0_12_prm_6_2_c_RNOZ0 ));
    InMux I__8792 (
            .O(N__40534),
            .I(N__40527));
    InMux I__8791 (
            .O(N__40533),
            .I(N__40524));
    InMux I__8790 (
            .O(N__40532),
            .I(N__40513));
    InMux I__8789 (
            .O(N__40531),
            .I(N__40513));
    InMux I__8788 (
            .O(N__40530),
            .I(N__40505));
    LocalMux I__8787 (
            .O(N__40527),
            .I(N__40501));
    LocalMux I__8786 (
            .O(N__40524),
            .I(N__40498));
    InMux I__8785 (
            .O(N__40523),
            .I(N__40495));
    InMux I__8784 (
            .O(N__40522),
            .I(N__40492));
    InMux I__8783 (
            .O(N__40521),
            .I(N__40489));
    InMux I__8782 (
            .O(N__40520),
            .I(N__40482));
    InMux I__8781 (
            .O(N__40519),
            .I(N__40477));
    InMux I__8780 (
            .O(N__40518),
            .I(N__40477));
    LocalMux I__8779 (
            .O(N__40513),
            .I(N__40474));
    InMux I__8778 (
            .O(N__40512),
            .I(N__40469));
    InMux I__8777 (
            .O(N__40511),
            .I(N__40469));
    InMux I__8776 (
            .O(N__40510),
            .I(N__40466));
    InMux I__8775 (
            .O(N__40509),
            .I(N__40461));
    InMux I__8774 (
            .O(N__40508),
            .I(N__40461));
    LocalMux I__8773 (
            .O(N__40505),
            .I(N__40458));
    InMux I__8772 (
            .O(N__40504),
            .I(N__40455));
    Span4Mux_h I__8771 (
            .O(N__40501),
            .I(N__40448));
    Span4Mux_s2_v I__8770 (
            .O(N__40498),
            .I(N__40448));
    LocalMux I__8769 (
            .O(N__40495),
            .I(N__40448));
    LocalMux I__8768 (
            .O(N__40492),
            .I(N__40445));
    LocalMux I__8767 (
            .O(N__40489),
            .I(N__40442));
    InMux I__8766 (
            .O(N__40488),
            .I(N__40439));
    InMux I__8765 (
            .O(N__40487),
            .I(N__40434));
    InMux I__8764 (
            .O(N__40486),
            .I(N__40434));
    InMux I__8763 (
            .O(N__40485),
            .I(N__40425));
    LocalMux I__8762 (
            .O(N__40482),
            .I(N__40420));
    LocalMux I__8761 (
            .O(N__40477),
            .I(N__40420));
    Span4Mux_v I__8760 (
            .O(N__40474),
            .I(N__40415));
    LocalMux I__8759 (
            .O(N__40469),
            .I(N__40415));
    LocalMux I__8758 (
            .O(N__40466),
            .I(N__40410));
    LocalMux I__8757 (
            .O(N__40461),
            .I(N__40410));
    Span4Mux_s2_h I__8756 (
            .O(N__40458),
            .I(N__40407));
    LocalMux I__8755 (
            .O(N__40455),
            .I(N__40404));
    Span4Mux_h I__8754 (
            .O(N__40448),
            .I(N__40401));
    Span12Mux_s4_v I__8753 (
            .O(N__40445),
            .I(N__40394));
    Span12Mux_v I__8752 (
            .O(N__40442),
            .I(N__40394));
    LocalMux I__8751 (
            .O(N__40439),
            .I(N__40394));
    LocalMux I__8750 (
            .O(N__40434),
            .I(N__40391));
    InMux I__8749 (
            .O(N__40433),
            .I(N__40386));
    InMux I__8748 (
            .O(N__40432),
            .I(N__40386));
    InMux I__8747 (
            .O(N__40431),
            .I(N__40381));
    InMux I__8746 (
            .O(N__40430),
            .I(N__40381));
    InMux I__8745 (
            .O(N__40429),
            .I(N__40376));
    InMux I__8744 (
            .O(N__40428),
            .I(N__40376));
    LocalMux I__8743 (
            .O(N__40425),
            .I(N__40371));
    Span4Mux_h I__8742 (
            .O(N__40420),
            .I(N__40371));
    Span4Mux_h I__8741 (
            .O(N__40415),
            .I(N__40366));
    Span4Mux_v I__8740 (
            .O(N__40410),
            .I(N__40366));
    Span4Mux_h I__8739 (
            .O(N__40407),
            .I(N__40361));
    Span4Mux_h I__8738 (
            .O(N__40404),
            .I(N__40361));
    Odrv4 I__8737 (
            .O(N__40401),
            .I(\ALU.b_4 ));
    Odrv12 I__8736 (
            .O(N__40394),
            .I(\ALU.b_4 ));
    Odrv12 I__8735 (
            .O(N__40391),
            .I(\ALU.b_4 ));
    LocalMux I__8734 (
            .O(N__40386),
            .I(\ALU.b_4 ));
    LocalMux I__8733 (
            .O(N__40381),
            .I(\ALU.b_4 ));
    LocalMux I__8732 (
            .O(N__40376),
            .I(\ALU.b_4 ));
    Odrv4 I__8731 (
            .O(N__40371),
            .I(\ALU.b_4 ));
    Odrv4 I__8730 (
            .O(N__40366),
            .I(\ALU.b_4 ));
    Odrv4 I__8729 (
            .O(N__40361),
            .I(\ALU.b_4 ));
    InMux I__8728 (
            .O(N__40342),
            .I(N__40339));
    LocalMux I__8727 (
            .O(N__40339),
            .I(\ALU.r0_12_prm_5_4_c_RNOZ0 ));
    InMux I__8726 (
            .O(N__40336),
            .I(N__40333));
    LocalMux I__8725 (
            .O(N__40333),
            .I(N__40330));
    Span4Mux_h I__8724 (
            .O(N__40330),
            .I(N__40327));
    Odrv4 I__8723 (
            .O(N__40327),
            .I(\ALU.r0_12_prm_5_2_c_RNOZ0 ));
    InMux I__8722 (
            .O(N__40324),
            .I(N__40321));
    LocalMux I__8721 (
            .O(N__40321),
            .I(N__40318));
    Span4Mux_h I__8720 (
            .O(N__40318),
            .I(N__40315));
    Odrv4 I__8719 (
            .O(N__40315),
            .I(\ALU.r4_RNIL9636Z0Z_2 ));
    CascadeMux I__8718 (
            .O(N__40312),
            .I(N__40309));
    InMux I__8717 (
            .O(N__40309),
            .I(N__40306));
    LocalMux I__8716 (
            .O(N__40306),
            .I(\ALU.a_i_2 ));
    InMux I__8715 (
            .O(N__40303),
            .I(\ALU.r0_12_2 ));
    InMux I__8714 (
            .O(N__40300),
            .I(N__40297));
    LocalMux I__8713 (
            .O(N__40297),
            .I(N__40293));
    InMux I__8712 (
            .O(N__40296),
            .I(N__40290));
    Span4Mux_v I__8711 (
            .O(N__40293),
            .I(N__40282));
    LocalMux I__8710 (
            .O(N__40290),
            .I(N__40282));
    InMux I__8709 (
            .O(N__40289),
            .I(N__40279));
    InMux I__8708 (
            .O(N__40288),
            .I(N__40276));
    InMux I__8707 (
            .O(N__40287),
            .I(N__40271));
    Span4Mux_v I__8706 (
            .O(N__40282),
            .I(N__40268));
    LocalMux I__8705 (
            .O(N__40279),
            .I(N__40263));
    LocalMux I__8704 (
            .O(N__40276),
            .I(N__40263));
    InMux I__8703 (
            .O(N__40275),
            .I(N__40260));
    InMux I__8702 (
            .O(N__40274),
            .I(N__40257));
    LocalMux I__8701 (
            .O(N__40271),
            .I(N__40254));
    Span4Mux_h I__8700 (
            .O(N__40268),
            .I(N__40251));
    Span4Mux_v I__8699 (
            .O(N__40263),
            .I(N__40244));
    LocalMux I__8698 (
            .O(N__40260),
            .I(N__40244));
    LocalMux I__8697 (
            .O(N__40257),
            .I(N__40244));
    Span4Mux_v I__8696 (
            .O(N__40254),
            .I(N__40240));
    Span4Mux_h I__8695 (
            .O(N__40251),
            .I(N__40235));
    Span4Mux_v I__8694 (
            .O(N__40244),
            .I(N__40235));
    InMux I__8693 (
            .O(N__40243),
            .I(N__40232));
    Span4Mux_v I__8692 (
            .O(N__40240),
            .I(N__40229));
    Span4Mux_h I__8691 (
            .O(N__40235),
            .I(N__40224));
    LocalMux I__8690 (
            .O(N__40232),
            .I(N__40224));
    Span4Mux_h I__8689 (
            .O(N__40229),
            .I(N__40221));
    Span4Mux_v I__8688 (
            .O(N__40224),
            .I(N__40218));
    Odrv4 I__8687 (
            .O(N__40221),
            .I(\ALU.r0_12_2_THRU_CO ));
    Odrv4 I__8686 (
            .O(N__40218),
            .I(\ALU.r0_12_2_THRU_CO ));
    CascadeMux I__8685 (
            .O(N__40213),
            .I(N__40210));
    InMux I__8684 (
            .O(N__40210),
            .I(N__40207));
    LocalMux I__8683 (
            .O(N__40207),
            .I(\ALU.lshift_2 ));
    InMux I__8682 (
            .O(N__40204),
            .I(N__40201));
    LocalMux I__8681 (
            .O(N__40201),
            .I(\ALU.r0_12_prm_8_2_c_RNOZ0 ));
    CascadeMux I__8680 (
            .O(N__40198),
            .I(N__40195));
    InMux I__8679 (
            .O(N__40195),
            .I(N__40192));
    LocalMux I__8678 (
            .O(N__40192),
            .I(N__40189));
    Span4Mux_h I__8677 (
            .O(N__40189),
            .I(N__40186));
    Odrv4 I__8676 (
            .O(N__40186),
            .I(\ALU.r0_12_prm_8_0_s0_c_RNOZ0 ));
    InMux I__8675 (
            .O(N__40183),
            .I(N__40177));
    InMux I__8674 (
            .O(N__40182),
            .I(N__40177));
    LocalMux I__8673 (
            .O(N__40177),
            .I(N__40170));
    InMux I__8672 (
            .O(N__40176),
            .I(N__40167));
    InMux I__8671 (
            .O(N__40175),
            .I(N__40164));
    CascadeMux I__8670 (
            .O(N__40174),
            .I(N__40161));
    InMux I__8669 (
            .O(N__40173),
            .I(N__40151));
    Span4Mux_h I__8668 (
            .O(N__40170),
            .I(N__40146));
    LocalMux I__8667 (
            .O(N__40167),
            .I(N__40146));
    LocalMux I__8666 (
            .O(N__40164),
            .I(N__40143));
    InMux I__8665 (
            .O(N__40161),
            .I(N__40135));
    InMux I__8664 (
            .O(N__40160),
            .I(N__40135));
    InMux I__8663 (
            .O(N__40159),
            .I(N__40135));
    InMux I__8662 (
            .O(N__40158),
            .I(N__40132));
    InMux I__8661 (
            .O(N__40157),
            .I(N__40129));
    InMux I__8660 (
            .O(N__40156),
            .I(N__40126));
    InMux I__8659 (
            .O(N__40155),
            .I(N__40123));
    InMux I__8658 (
            .O(N__40154),
            .I(N__40120));
    LocalMux I__8657 (
            .O(N__40151),
            .I(N__40115));
    Span4Mux_v I__8656 (
            .O(N__40146),
            .I(N__40115));
    Span4Mux_h I__8655 (
            .O(N__40143),
            .I(N__40110));
    InMux I__8654 (
            .O(N__40142),
            .I(N__40107));
    LocalMux I__8653 (
            .O(N__40135),
            .I(N__40103));
    LocalMux I__8652 (
            .O(N__40132),
            .I(N__40098));
    LocalMux I__8651 (
            .O(N__40129),
            .I(N__40098));
    LocalMux I__8650 (
            .O(N__40126),
            .I(N__40092));
    LocalMux I__8649 (
            .O(N__40123),
            .I(N__40092));
    LocalMux I__8648 (
            .O(N__40120),
            .I(N__40087));
    Span4Mux_v I__8647 (
            .O(N__40115),
            .I(N__40087));
    InMux I__8646 (
            .O(N__40114),
            .I(N__40081));
    InMux I__8645 (
            .O(N__40113),
            .I(N__40078));
    Span4Mux_v I__8644 (
            .O(N__40110),
            .I(N__40075));
    LocalMux I__8643 (
            .O(N__40107),
            .I(N__40072));
    InMux I__8642 (
            .O(N__40106),
            .I(N__40069));
    Span4Mux_v I__8641 (
            .O(N__40103),
            .I(N__40066));
    Span4Mux_v I__8640 (
            .O(N__40098),
            .I(N__40063));
    InMux I__8639 (
            .O(N__40097),
            .I(N__40060));
    Span4Mux_v I__8638 (
            .O(N__40092),
            .I(N__40055));
    Span4Mux_v I__8637 (
            .O(N__40087),
            .I(N__40055));
    InMux I__8636 (
            .O(N__40086),
            .I(N__40049));
    InMux I__8635 (
            .O(N__40085),
            .I(N__40049));
    InMux I__8634 (
            .O(N__40084),
            .I(N__40046));
    LocalMux I__8633 (
            .O(N__40081),
            .I(N__40039));
    LocalMux I__8632 (
            .O(N__40078),
            .I(N__40039));
    Span4Mux_h I__8631 (
            .O(N__40075),
            .I(N__40039));
    Span4Mux_h I__8630 (
            .O(N__40072),
            .I(N__40036));
    LocalMux I__8629 (
            .O(N__40069),
            .I(N__40025));
    Sp12to4 I__8628 (
            .O(N__40066),
            .I(N__40025));
    Sp12to4 I__8627 (
            .O(N__40063),
            .I(N__40025));
    LocalMux I__8626 (
            .O(N__40060),
            .I(N__40025));
    Sp12to4 I__8625 (
            .O(N__40055),
            .I(N__40025));
    InMux I__8624 (
            .O(N__40054),
            .I(N__40022));
    LocalMux I__8623 (
            .O(N__40049),
            .I(\ALU.a_15 ));
    LocalMux I__8622 (
            .O(N__40046),
            .I(\ALU.a_15 ));
    Odrv4 I__8621 (
            .O(N__40039),
            .I(\ALU.a_15 ));
    Odrv4 I__8620 (
            .O(N__40036),
            .I(\ALU.a_15 ));
    Odrv12 I__8619 (
            .O(N__40025),
            .I(\ALU.a_15 ));
    LocalMux I__8618 (
            .O(N__40022),
            .I(\ALU.a_15 ));
    InMux I__8617 (
            .O(N__40009),
            .I(N__40004));
    InMux I__8616 (
            .O(N__40008),
            .I(N__40001));
    InMux I__8615 (
            .O(N__40007),
            .I(N__39998));
    LocalMux I__8614 (
            .O(N__40004),
            .I(N__39995));
    LocalMux I__8613 (
            .O(N__40001),
            .I(N__39989));
    LocalMux I__8612 (
            .O(N__39998),
            .I(N__39985));
    Span4Mux_h I__8611 (
            .O(N__39995),
            .I(N__39982));
    InMux I__8610 (
            .O(N__39994),
            .I(N__39974));
    InMux I__8609 (
            .O(N__39993),
            .I(N__39974));
    InMux I__8608 (
            .O(N__39992),
            .I(N__39974));
    Span4Mux_h I__8607 (
            .O(N__39989),
            .I(N__39970));
    InMux I__8606 (
            .O(N__39988),
            .I(N__39967));
    Span4Mux_h I__8605 (
            .O(N__39985),
            .I(N__39964));
    Span4Mux_v I__8604 (
            .O(N__39982),
            .I(N__39961));
    InMux I__8603 (
            .O(N__39981),
            .I(N__39958));
    LocalMux I__8602 (
            .O(N__39974),
            .I(N__39954));
    InMux I__8601 (
            .O(N__39973),
            .I(N__39951));
    Span4Mux_v I__8600 (
            .O(N__39970),
            .I(N__39946));
    LocalMux I__8599 (
            .O(N__39967),
            .I(N__39946));
    Span4Mux_h I__8598 (
            .O(N__39964),
            .I(N__39943));
    Sp12to4 I__8597 (
            .O(N__39961),
            .I(N__39938));
    LocalMux I__8596 (
            .O(N__39958),
            .I(N__39938));
    InMux I__8595 (
            .O(N__39957),
            .I(N__39935));
    Span4Mux_h I__8594 (
            .O(N__39954),
            .I(N__39932));
    LocalMux I__8593 (
            .O(N__39951),
            .I(N__39929));
    Span4Mux_h I__8592 (
            .O(N__39946),
            .I(N__39926));
    Span4Mux_v I__8591 (
            .O(N__39943),
            .I(N__39922));
    Span12Mux_h I__8590 (
            .O(N__39938),
            .I(N__39919));
    LocalMux I__8589 (
            .O(N__39935),
            .I(N__39910));
    Span4Mux_h I__8588 (
            .O(N__39932),
            .I(N__39910));
    Span4Mux_s2_h I__8587 (
            .O(N__39929),
            .I(N__39910));
    Span4Mux_h I__8586 (
            .O(N__39926),
            .I(N__39910));
    InMux I__8585 (
            .O(N__39925),
            .I(N__39907));
    Odrv4 I__8584 (
            .O(N__39922),
            .I(\ALU.b_15 ));
    Odrv12 I__8583 (
            .O(N__39919),
            .I(\ALU.b_15 ));
    Odrv4 I__8582 (
            .O(N__39910),
            .I(\ALU.b_15 ));
    LocalMux I__8581 (
            .O(N__39907),
            .I(\ALU.b_15 ));
    InMux I__8580 (
            .O(N__39898),
            .I(N__39895));
    LocalMux I__8579 (
            .O(N__39895),
            .I(N__39892));
    Odrv4 I__8578 (
            .O(N__39892),
            .I(\ALU.r0_12_prm_7_15_s0_c_RNOZ0 ));
    InMux I__8577 (
            .O(N__39889),
            .I(N__39886));
    LocalMux I__8576 (
            .O(N__39886),
            .I(N__39883));
    Span4Mux_h I__8575 (
            .O(N__39883),
            .I(N__39880));
    Odrv4 I__8574 (
            .O(N__39880),
            .I(\ALU.r0_12_prm_8_13_s1_c_RNOZ0Z_1 ));
    InMux I__8573 (
            .O(N__39877),
            .I(N__39867));
    InMux I__8572 (
            .O(N__39876),
            .I(N__39867));
    CascadeMux I__8571 (
            .O(N__39875),
            .I(N__39864));
    InMux I__8570 (
            .O(N__39874),
            .I(N__39854));
    InMux I__8569 (
            .O(N__39873),
            .I(N__39854));
    InMux I__8568 (
            .O(N__39872),
            .I(N__39851));
    LocalMux I__8567 (
            .O(N__39867),
            .I(N__39846));
    InMux I__8566 (
            .O(N__39864),
            .I(N__39843));
    InMux I__8565 (
            .O(N__39863),
            .I(N__39838));
    InMux I__8564 (
            .O(N__39862),
            .I(N__39838));
    InMux I__8563 (
            .O(N__39861),
            .I(N__39834));
    InMux I__8562 (
            .O(N__39860),
            .I(N__39831));
    InMux I__8561 (
            .O(N__39859),
            .I(N__39827));
    LocalMux I__8560 (
            .O(N__39854),
            .I(N__39823));
    LocalMux I__8559 (
            .O(N__39851),
            .I(N__39820));
    CascadeMux I__8558 (
            .O(N__39850),
            .I(N__39817));
    CascadeMux I__8557 (
            .O(N__39849),
            .I(N__39814));
    Span4Mux_v I__8556 (
            .O(N__39846),
            .I(N__39808));
    LocalMux I__8555 (
            .O(N__39843),
            .I(N__39808));
    LocalMux I__8554 (
            .O(N__39838),
            .I(N__39805));
    InMux I__8553 (
            .O(N__39837),
            .I(N__39802));
    LocalMux I__8552 (
            .O(N__39834),
            .I(N__39797));
    LocalMux I__8551 (
            .O(N__39831),
            .I(N__39797));
    InMux I__8550 (
            .O(N__39830),
            .I(N__39794));
    LocalMux I__8549 (
            .O(N__39827),
            .I(N__39791));
    InMux I__8548 (
            .O(N__39826),
            .I(N__39788));
    Span4Mux_v I__8547 (
            .O(N__39823),
            .I(N__39783));
    Span4Mux_v I__8546 (
            .O(N__39820),
            .I(N__39783));
    InMux I__8545 (
            .O(N__39817),
            .I(N__39780));
    InMux I__8544 (
            .O(N__39814),
            .I(N__39775));
    InMux I__8543 (
            .O(N__39813),
            .I(N__39775));
    Span4Mux_h I__8542 (
            .O(N__39808),
            .I(N__39772));
    Span4Mux_s2_h I__8541 (
            .O(N__39805),
            .I(N__39769));
    LocalMux I__8540 (
            .O(N__39802),
            .I(N__39766));
    Span4Mux_h I__8539 (
            .O(N__39797),
            .I(N__39763));
    LocalMux I__8538 (
            .O(N__39794),
            .I(N__39758));
    Span4Mux_v I__8537 (
            .O(N__39791),
            .I(N__39758));
    LocalMux I__8536 (
            .O(N__39788),
            .I(N__39755));
    Sp12to4 I__8535 (
            .O(N__39783),
            .I(N__39752));
    LocalMux I__8534 (
            .O(N__39780),
            .I(N__39747));
    LocalMux I__8533 (
            .O(N__39775),
            .I(N__39747));
    Span4Mux_h I__8532 (
            .O(N__39772),
            .I(N__39744));
    Span4Mux_v I__8531 (
            .O(N__39769),
            .I(N__39739));
    Span4Mux_s2_h I__8530 (
            .O(N__39766),
            .I(N__39739));
    Span4Mux_h I__8529 (
            .O(N__39763),
            .I(N__39732));
    Span4Mux_h I__8528 (
            .O(N__39758),
            .I(N__39732));
    Span4Mux_v I__8527 (
            .O(N__39755),
            .I(N__39732));
    Span12Mux_h I__8526 (
            .O(N__39752),
            .I(N__39727));
    Sp12to4 I__8525 (
            .O(N__39747),
            .I(N__39727));
    Odrv4 I__8524 (
            .O(N__39744),
            .I(\ALU.b_12 ));
    Odrv4 I__8523 (
            .O(N__39739),
            .I(\ALU.b_12 ));
    Odrv4 I__8522 (
            .O(N__39732),
            .I(\ALU.b_12 ));
    Odrv12 I__8521 (
            .O(N__39727),
            .I(\ALU.b_12 ));
    CascadeMux I__8520 (
            .O(N__39718),
            .I(N__39715));
    InMux I__8519 (
            .O(N__39715),
            .I(N__39712));
    LocalMux I__8518 (
            .O(N__39712),
            .I(\ALU.r0_12_prm_6_12_s1_c_RNOZ0 ));
    InMux I__8517 (
            .O(N__39709),
            .I(N__39706));
    LocalMux I__8516 (
            .O(N__39706),
            .I(N__39703));
    Odrv4 I__8515 (
            .O(N__39703),
            .I(\ALU.r5_RNIPV8A9_0Z0Z_13 ));
    CascadeMux I__8514 (
            .O(N__39700),
            .I(N__39697));
    InMux I__8513 (
            .O(N__39697),
            .I(N__39693));
    InMux I__8512 (
            .O(N__39696),
            .I(N__39690));
    LocalMux I__8511 (
            .O(N__39693),
            .I(\ALU.rshift_2 ));
    LocalMux I__8510 (
            .O(N__39690),
            .I(\ALU.rshift_2 ));
    CascadeMux I__8509 (
            .O(N__39685),
            .I(N__39682));
    InMux I__8508 (
            .O(N__39682),
            .I(N__39679));
    LocalMux I__8507 (
            .O(N__39679),
            .I(N__39676));
    Span4Mux_h I__8506 (
            .O(N__39676),
            .I(N__39673));
    Span4Mux_h I__8505 (
            .O(N__39673),
            .I(N__39670));
    Odrv4 I__8504 (
            .O(N__39670),
            .I(\ALU.r5_RNITG1F5Z0Z_14 ));
    InMux I__8503 (
            .O(N__39667),
            .I(N__39664));
    LocalMux I__8502 (
            .O(N__39664),
            .I(N__39661));
    Odrv12 I__8501 (
            .O(N__39661),
            .I(\ALU.r0_12_prm_5_14_s0_c_RNOZ0 ));
    InMux I__8500 (
            .O(N__39658),
            .I(N__39655));
    LocalMux I__8499 (
            .O(N__39655),
            .I(N__39652));
    Span12Mux_v I__8498 (
            .O(N__39652),
            .I(N__39649));
    Odrv12 I__8497 (
            .O(N__39649),
            .I(\ALU.rshift_13 ));
    CascadeMux I__8496 (
            .O(N__39646),
            .I(N__39643));
    InMux I__8495 (
            .O(N__39643),
            .I(N__39640));
    LocalMux I__8494 (
            .O(N__39640),
            .I(N__39637));
    Odrv12 I__8493 (
            .O(N__39637),
            .I(\ALU.r0_12_prm_6_14_s0_c_RNOZ0 ));
    CascadeMux I__8492 (
            .O(N__39634),
            .I(N__39631));
    InMux I__8491 (
            .O(N__39631),
            .I(N__39628));
    LocalMux I__8490 (
            .O(N__39628),
            .I(N__39625));
    Odrv12 I__8489 (
            .O(N__39625),
            .I(\ALU.r0_12_prm_8_14_s0_c_RNOZ0 ));
    InMux I__8488 (
            .O(N__39622),
            .I(N__39619));
    LocalMux I__8487 (
            .O(N__39619),
            .I(N__39613));
    InMux I__8486 (
            .O(N__39618),
            .I(N__39606));
    InMux I__8485 (
            .O(N__39617),
            .I(N__39606));
    InMux I__8484 (
            .O(N__39616),
            .I(N__39606));
    Span4Mux_v I__8483 (
            .O(N__39613),
            .I(N__39603));
    LocalMux I__8482 (
            .O(N__39606),
            .I(N__39600));
    Sp12to4 I__8481 (
            .O(N__39603),
            .I(N__39597));
    Span4Mux_v I__8480 (
            .O(N__39600),
            .I(N__39594));
    Odrv12 I__8479 (
            .O(N__39597),
            .I(\ALU.un9_addsub_cry_7_c_RNINZ0Z3519 ));
    Odrv4 I__8478 (
            .O(N__39594),
            .I(\ALU.un9_addsub_cry_7_c_RNINZ0Z3519 ));
    CascadeMux I__8477 (
            .O(N__39589),
            .I(N__39586));
    InMux I__8476 (
            .O(N__39586),
            .I(N__39583));
    LocalMux I__8475 (
            .O(N__39583),
            .I(\ALU.r0_12_prm_1_8_s1_c_RNOZ0 ));
    InMux I__8474 (
            .O(N__39580),
            .I(N__39577));
    LocalMux I__8473 (
            .O(N__39577),
            .I(N__39574));
    Span4Mux_h I__8472 (
            .O(N__39574),
            .I(N__39571));
    Span4Mux_h I__8471 (
            .O(N__39571),
            .I(N__39568));
    Span4Mux_v I__8470 (
            .O(N__39568),
            .I(N__39565));
    Odrv4 I__8469 (
            .O(N__39565),
            .I(\ALU.madd_cry_6_THRU_CO ));
    InMux I__8468 (
            .O(N__39562),
            .I(N__39558));
    InMux I__8467 (
            .O(N__39561),
            .I(N__39555));
    LocalMux I__8466 (
            .O(N__39558),
            .I(N__39552));
    LocalMux I__8465 (
            .O(N__39555),
            .I(N__39549));
    Span12Mux_v I__8464 (
            .O(N__39552),
            .I(N__39546));
    Span4Mux_v I__8463 (
            .O(N__39549),
            .I(N__39543));
    Odrv12 I__8462 (
            .O(N__39546),
            .I(\ALU.madd_axb_7 ));
    Odrv4 I__8461 (
            .O(N__39543),
            .I(\ALU.madd_axb_7 ));
    CascadeMux I__8460 (
            .O(N__39538),
            .I(N__39535));
    InMux I__8459 (
            .O(N__39535),
            .I(N__39532));
    LocalMux I__8458 (
            .O(N__39532),
            .I(\ALU.r0_12_s0_8_THRU_CO ));
    InMux I__8457 (
            .O(N__39529),
            .I(\ALU.r0_12_s1_8 ));
    InMux I__8456 (
            .O(N__39526),
            .I(N__39520));
    InMux I__8455 (
            .O(N__39525),
            .I(N__39517));
    InMux I__8454 (
            .O(N__39524),
            .I(N__39514));
    InMux I__8453 (
            .O(N__39523),
            .I(N__39510));
    LocalMux I__8452 (
            .O(N__39520),
            .I(N__39507));
    LocalMux I__8451 (
            .O(N__39517),
            .I(N__39504));
    LocalMux I__8450 (
            .O(N__39514),
            .I(N__39501));
    InMux I__8449 (
            .O(N__39513),
            .I(N__39498));
    LocalMux I__8448 (
            .O(N__39510),
            .I(N__39495));
    Span4Mux_h I__8447 (
            .O(N__39507),
            .I(N__39490));
    Span4Mux_h I__8446 (
            .O(N__39504),
            .I(N__39485));
    Span4Mux_v I__8445 (
            .O(N__39501),
            .I(N__39485));
    LocalMux I__8444 (
            .O(N__39498),
            .I(N__39482));
    Span4Mux_h I__8443 (
            .O(N__39495),
            .I(N__39479));
    InMux I__8442 (
            .O(N__39494),
            .I(N__39476));
    InMux I__8441 (
            .O(N__39493),
            .I(N__39473));
    Span4Mux_h I__8440 (
            .O(N__39490),
            .I(N__39469));
    Span4Mux_h I__8439 (
            .O(N__39485),
            .I(N__39466));
    Span4Mux_h I__8438 (
            .O(N__39482),
            .I(N__39463));
    Span4Mux_h I__8437 (
            .O(N__39479),
            .I(N__39458));
    LocalMux I__8436 (
            .O(N__39476),
            .I(N__39458));
    LocalMux I__8435 (
            .O(N__39473),
            .I(N__39455));
    InMux I__8434 (
            .O(N__39472),
            .I(N__39452));
    Odrv4 I__8433 (
            .O(N__39469),
            .I(\ALU.r0_12_8 ));
    Odrv4 I__8432 (
            .O(N__39466),
            .I(\ALU.r0_12_8 ));
    Odrv4 I__8431 (
            .O(N__39463),
            .I(\ALU.r0_12_8 ));
    Odrv4 I__8430 (
            .O(N__39458),
            .I(\ALU.r0_12_8 ));
    Odrv12 I__8429 (
            .O(N__39455),
            .I(\ALU.r0_12_8 ));
    LocalMux I__8428 (
            .O(N__39452),
            .I(\ALU.r0_12_8 ));
    InMux I__8427 (
            .O(N__39439),
            .I(N__39435));
    InMux I__8426 (
            .O(N__39438),
            .I(N__39432));
    LocalMux I__8425 (
            .O(N__39435),
            .I(N__39428));
    LocalMux I__8424 (
            .O(N__39432),
            .I(N__39425));
    InMux I__8423 (
            .O(N__39431),
            .I(N__39422));
    Span4Mux_h I__8422 (
            .O(N__39428),
            .I(N__39419));
    Span4Mux_h I__8421 (
            .O(N__39425),
            .I(N__39414));
    LocalMux I__8420 (
            .O(N__39422),
            .I(N__39414));
    Span4Mux_h I__8419 (
            .O(N__39419),
            .I(N__39411));
    Span4Mux_h I__8418 (
            .O(N__39414),
            .I(N__39408));
    Odrv4 I__8417 (
            .O(N__39411),
            .I(r0_8));
    Odrv4 I__8416 (
            .O(N__39408),
            .I(r0_8));
    InMux I__8415 (
            .O(N__39403),
            .I(N__39398));
    InMux I__8414 (
            .O(N__39402),
            .I(N__39395));
    InMux I__8413 (
            .O(N__39401),
            .I(N__39392));
    LocalMux I__8412 (
            .O(N__39398),
            .I(N__39388));
    LocalMux I__8411 (
            .O(N__39395),
            .I(N__39383));
    LocalMux I__8410 (
            .O(N__39392),
            .I(N__39383));
    InMux I__8409 (
            .O(N__39391),
            .I(N__39380));
    Span4Mux_h I__8408 (
            .O(N__39388),
            .I(N__39377));
    Odrv4 I__8407 (
            .O(N__39383),
            .I(\ALU.un2_addsub_cry_7_c_RNI5ELEEZ0 ));
    LocalMux I__8406 (
            .O(N__39380),
            .I(\ALU.un2_addsub_cry_7_c_RNI5ELEEZ0 ));
    Odrv4 I__8405 (
            .O(N__39377),
            .I(\ALU.un2_addsub_cry_7_c_RNI5ELEEZ0 ));
    CascadeMux I__8404 (
            .O(N__39370),
            .I(N__39367));
    InMux I__8403 (
            .O(N__39367),
            .I(N__39364));
    LocalMux I__8402 (
            .O(N__39364),
            .I(N__39361));
    Odrv4 I__8401 (
            .O(N__39361),
            .I(\ALU.r0_12_prm_2_8_s0_c_RNOZ0 ));
    InMux I__8400 (
            .O(N__39358),
            .I(N__39355));
    LocalMux I__8399 (
            .O(N__39355),
            .I(N__39352));
    Odrv4 I__8398 (
            .O(N__39352),
            .I(\ALU.r5_RNITTMB9Z0Z_12 ));
    CascadeMux I__8397 (
            .O(N__39349),
            .I(\ALU.r5_RNITTMB9Z0Z_12_cascade_ ));
    CascadeMux I__8396 (
            .O(N__39346),
            .I(\ALU.rshift_15_ns_1_1_cascade_ ));
    CascadeMux I__8395 (
            .O(N__39343),
            .I(N__39340));
    InMux I__8394 (
            .O(N__39340),
            .I(N__39337));
    LocalMux I__8393 (
            .O(N__39337),
            .I(N__39334));
    Odrv12 I__8392 (
            .O(N__39334),
            .I(\ALU.r0_12_prm_8_8_s1_c_RNOZ0Z_1 ));
    CascadeMux I__8391 (
            .O(N__39331),
            .I(N__39328));
    InMux I__8390 (
            .O(N__39328),
            .I(N__39324));
    InMux I__8389 (
            .O(N__39327),
            .I(N__39321));
    LocalMux I__8388 (
            .O(N__39324),
            .I(N__39318));
    LocalMux I__8387 (
            .O(N__39321),
            .I(N__39312));
    Span4Mux_h I__8386 (
            .O(N__39318),
            .I(N__39312));
    InMux I__8385 (
            .O(N__39317),
            .I(N__39309));
    Odrv4 I__8384 (
            .O(N__39312),
            .I(\ALU.lshift_8 ));
    LocalMux I__8383 (
            .O(N__39309),
            .I(\ALU.lshift_8 ));
    CascadeMux I__8382 (
            .O(N__39304),
            .I(N__39301));
    InMux I__8381 (
            .O(N__39301),
            .I(N__39298));
    LocalMux I__8380 (
            .O(N__39298),
            .I(N__39295));
    Odrv12 I__8379 (
            .O(N__39295),
            .I(\ALU.r0_12_prm_8_8_s1_c_RNOZ0 ));
    CascadeMux I__8378 (
            .O(N__39292),
            .I(N__39288));
    InMux I__8377 (
            .O(N__39291),
            .I(N__39285));
    InMux I__8376 (
            .O(N__39288),
            .I(N__39282));
    LocalMux I__8375 (
            .O(N__39285),
            .I(N__39277));
    LocalMux I__8374 (
            .O(N__39282),
            .I(N__39277));
    Span4Mux_v I__8373 (
            .O(N__39277),
            .I(N__39274));
    Span4Mux_v I__8372 (
            .O(N__39274),
            .I(N__39271));
    Sp12to4 I__8371 (
            .O(N__39271),
            .I(N__39268));
    Odrv12 I__8370 (
            .O(N__39268),
            .I(\ALU.a8_b_8 ));
    InMux I__8369 (
            .O(N__39265),
            .I(N__39261));
    CascadeMux I__8368 (
            .O(N__39264),
            .I(N__39258));
    LocalMux I__8367 (
            .O(N__39261),
            .I(N__39255));
    InMux I__8366 (
            .O(N__39258),
            .I(N__39252));
    Span4Mux_h I__8365 (
            .O(N__39255),
            .I(N__39247));
    LocalMux I__8364 (
            .O(N__39252),
            .I(N__39247));
    Span4Mux_v I__8363 (
            .O(N__39247),
            .I(N__39244));
    Odrv4 I__8362 (
            .O(N__39244),
            .I(\ALU.un14_log_0_i_8 ));
    InMux I__8361 (
            .O(N__39241),
            .I(N__39238));
    LocalMux I__8360 (
            .O(N__39238),
            .I(\ALU.r0_12_prm_4_8_s1_c_RNOZ0 ));
    CascadeMux I__8359 (
            .O(N__39235),
            .I(N__39231));
    CascadeMux I__8358 (
            .O(N__39234),
            .I(N__39228));
    InMux I__8357 (
            .O(N__39231),
            .I(N__39225));
    InMux I__8356 (
            .O(N__39228),
            .I(N__39222));
    LocalMux I__8355 (
            .O(N__39225),
            .I(\ALU.a_i_8 ));
    LocalMux I__8354 (
            .O(N__39222),
            .I(\ALU.a_i_8 ));
    CascadeMux I__8353 (
            .O(N__39217),
            .I(N__39214));
    InMux I__8352 (
            .O(N__39214),
            .I(N__39211));
    LocalMux I__8351 (
            .O(N__39211),
            .I(N__39208));
    Odrv4 I__8350 (
            .O(N__39208),
            .I(\ALU.r0_12_prm_2_8_s1_c_RNOZ0 ));
    InMux I__8349 (
            .O(N__39205),
            .I(N__39202));
    LocalMux I__8348 (
            .O(N__39202),
            .I(N__39197));
    InMux I__8347 (
            .O(N__39201),
            .I(N__39192));
    InMux I__8346 (
            .O(N__39200),
            .I(N__39192));
    Span4Mux_h I__8345 (
            .O(N__39197),
            .I(N__39189));
    LocalMux I__8344 (
            .O(N__39192),
            .I(N__39186));
    Sp12to4 I__8343 (
            .O(N__39189),
            .I(N__39183));
    Span4Mux_h I__8342 (
            .O(N__39186),
            .I(N__39180));
    Span12Mux_v I__8341 (
            .O(N__39183),
            .I(N__39177));
    Span4Mux_h I__8340 (
            .O(N__39180),
            .I(N__39174));
    Odrv12 I__8339 (
            .O(N__39177),
            .I(r6_8));
    Odrv4 I__8338 (
            .O(N__39174),
            .I(r6_8));
    InMux I__8337 (
            .O(N__39169),
            .I(N__39164));
    InMux I__8336 (
            .O(N__39168),
            .I(N__39159));
    InMux I__8335 (
            .O(N__39167),
            .I(N__39159));
    LocalMux I__8334 (
            .O(N__39164),
            .I(N__39156));
    LocalMux I__8333 (
            .O(N__39159),
            .I(N__39153));
    Span4Mux_h I__8332 (
            .O(N__39156),
            .I(N__39150));
    Span12Mux_s5_h I__8331 (
            .O(N__39153),
            .I(N__39147));
    Span4Mux_h I__8330 (
            .O(N__39150),
            .I(N__39144));
    Odrv12 I__8329 (
            .O(N__39147),
            .I(r6_2));
    Odrv4 I__8328 (
            .O(N__39144),
            .I(r6_2));
    InMux I__8327 (
            .O(N__39139),
            .I(N__39136));
    LocalMux I__8326 (
            .O(N__39136),
            .I(N__39133));
    Span4Mux_v I__8325 (
            .O(N__39133),
            .I(N__39129));
    InMux I__8324 (
            .O(N__39132),
            .I(N__39125));
    Span4Mux_h I__8323 (
            .O(N__39129),
            .I(N__39122));
    InMux I__8322 (
            .O(N__39128),
            .I(N__39119));
    LocalMux I__8321 (
            .O(N__39125),
            .I(N__39116));
    Span4Mux_h I__8320 (
            .O(N__39122),
            .I(N__39113));
    LocalMux I__8319 (
            .O(N__39119),
            .I(N__39110));
    Span4Mux_h I__8318 (
            .O(N__39116),
            .I(N__39107));
    Span4Mux_h I__8317 (
            .O(N__39113),
            .I(N__39104));
    Span12Mux_v I__8316 (
            .O(N__39110),
            .I(N__39101));
    Span4Mux_h I__8315 (
            .O(N__39107),
            .I(N__39098));
    Odrv4 I__8314 (
            .O(N__39104),
            .I(r6_3));
    Odrv12 I__8313 (
            .O(N__39101),
            .I(r6_3));
    Odrv4 I__8312 (
            .O(N__39098),
            .I(r6_3));
    InMux I__8311 (
            .O(N__39091),
            .I(N__39087));
    InMux I__8310 (
            .O(N__39090),
            .I(N__39084));
    LocalMux I__8309 (
            .O(N__39087),
            .I(N__39079));
    LocalMux I__8308 (
            .O(N__39084),
            .I(N__39075));
    InMux I__8307 (
            .O(N__39083),
            .I(N__39072));
    InMux I__8306 (
            .O(N__39082),
            .I(N__39069));
    Span4Mux_h I__8305 (
            .O(N__39079),
            .I(N__39066));
    InMux I__8304 (
            .O(N__39078),
            .I(N__39063));
    Span4Mux_v I__8303 (
            .O(N__39075),
            .I(N__39059));
    LocalMux I__8302 (
            .O(N__39072),
            .I(N__39056));
    LocalMux I__8301 (
            .O(N__39069),
            .I(N__39053));
    Span4Mux_v I__8300 (
            .O(N__39066),
            .I(N__39047));
    LocalMux I__8299 (
            .O(N__39063),
            .I(N__39047));
    InMux I__8298 (
            .O(N__39062),
            .I(N__39044));
    Span4Mux_h I__8297 (
            .O(N__39059),
            .I(N__39038));
    Span4Mux_h I__8296 (
            .O(N__39056),
            .I(N__39038));
    Span4Mux_h I__8295 (
            .O(N__39053),
            .I(N__39035));
    InMux I__8294 (
            .O(N__39052),
            .I(N__39032));
    Span4Mux_v I__8293 (
            .O(N__39047),
            .I(N__39027));
    LocalMux I__8292 (
            .O(N__39044),
            .I(N__39027));
    InMux I__8291 (
            .O(N__39043),
            .I(N__39024));
    Span4Mux_v I__8290 (
            .O(N__39038),
            .I(N__39021));
    Span4Mux_v I__8289 (
            .O(N__39035),
            .I(N__39018));
    LocalMux I__8288 (
            .O(N__39032),
            .I(N__39015));
    Span4Mux_h I__8287 (
            .O(N__39027),
            .I(N__39010));
    LocalMux I__8286 (
            .O(N__39024),
            .I(N__39010));
    Odrv4 I__8285 (
            .O(N__39021),
            .I(\ALU.r0_12_4_THRU_CO ));
    Odrv4 I__8284 (
            .O(N__39018),
            .I(\ALU.r0_12_4_THRU_CO ));
    Odrv12 I__8283 (
            .O(N__39015),
            .I(\ALU.r0_12_4_THRU_CO ));
    Odrv4 I__8282 (
            .O(N__39010),
            .I(\ALU.r0_12_4_THRU_CO ));
    InMux I__8281 (
            .O(N__39001),
            .I(N__38992));
    InMux I__8280 (
            .O(N__39000),
            .I(N__38992));
    InMux I__8279 (
            .O(N__38999),
            .I(N__38992));
    LocalMux I__8278 (
            .O(N__38992),
            .I(N__38989));
    Span4Mux_h I__8277 (
            .O(N__38989),
            .I(N__38986));
    Span4Mux_h I__8276 (
            .O(N__38986),
            .I(N__38983));
    Odrv4 I__8275 (
            .O(N__38983),
            .I(r6_4));
    InMux I__8274 (
            .O(N__38980),
            .I(N__38977));
    LocalMux I__8273 (
            .O(N__38977),
            .I(\ALU.r4_RNIN3236Z0Z_8 ));
    InMux I__8272 (
            .O(N__38974),
            .I(N__38971));
    LocalMux I__8271 (
            .O(N__38971),
            .I(N__38968));
    Span4Mux_v I__8270 (
            .O(N__38968),
            .I(N__38965));
    Span4Mux_h I__8269 (
            .O(N__38965),
            .I(N__38962));
    Span4Mux_h I__8268 (
            .O(N__38962),
            .I(N__38959));
    Odrv4 I__8267 (
            .O(N__38959),
            .I(\ALU.rshift_3_ns_1_1 ));
    CascadeMux I__8266 (
            .O(N__38956),
            .I(\ALU.r0_12_prm_8_1_c_RNOZ0Z_3_cascade_ ));
    CascadeMux I__8265 (
            .O(N__38953),
            .I(N__38950));
    InMux I__8264 (
            .O(N__38950),
            .I(N__38947));
    LocalMux I__8263 (
            .O(N__38947),
            .I(\ALU.r0_12_prm_2_7_s0_c_RNOZ0 ));
    InMux I__8262 (
            .O(N__38944),
            .I(N__38940));
    InMux I__8261 (
            .O(N__38943),
            .I(N__38937));
    LocalMux I__8260 (
            .O(N__38940),
            .I(N__38934));
    LocalMux I__8259 (
            .O(N__38937),
            .I(N__38931));
    Span4Mux_h I__8258 (
            .O(N__38934),
            .I(N__38928));
    Span12Mux_v I__8257 (
            .O(N__38931),
            .I(N__38925));
    Odrv4 I__8256 (
            .O(N__38928),
            .I(\ALU.r4_RNIODO6KZ0Z_5 ));
    Odrv12 I__8255 (
            .O(N__38925),
            .I(\ALU.r4_RNIODO6KZ0Z_5 ));
    CascadeMux I__8254 (
            .O(N__38920),
            .I(\ALU.lshift_8_cascade_ ));
    InMux I__8253 (
            .O(N__38917),
            .I(N__38914));
    LocalMux I__8252 (
            .O(N__38914),
            .I(N__38911));
    Span4Mux_h I__8251 (
            .O(N__38911),
            .I(N__38908));
    Odrv4 I__8250 (
            .O(N__38908),
            .I(\ALU.r0_12_prm_8_8_s0_c_RNOZ0 ));
    InMux I__8249 (
            .O(N__38905),
            .I(N__38902));
    LocalMux I__8248 (
            .O(N__38902),
            .I(N__38899));
    Span4Mux_v I__8247 (
            .O(N__38899),
            .I(N__38896));
    Odrv4 I__8246 (
            .O(N__38896),
            .I(\ALU.r0_12_prm_8_12_s1_c_RNOZ0Z_1 ));
    InMux I__8245 (
            .O(N__38893),
            .I(N__38890));
    LocalMux I__8244 (
            .O(N__38890),
            .I(N__38887));
    Odrv4 I__8243 (
            .O(N__38887),
            .I(\ALU.r0_12_prm_7_8_s0_c_RNOZ0 ));
    InMux I__8242 (
            .O(N__38884),
            .I(N__38881));
    LocalMux I__8241 (
            .O(N__38881),
            .I(\ALU.rshift_5 ));
    InMux I__8240 (
            .O(N__38878),
            .I(N__38875));
    LocalMux I__8239 (
            .O(N__38875),
            .I(N__38868));
    InMux I__8238 (
            .O(N__38874),
            .I(N__38865));
    InMux I__8237 (
            .O(N__38873),
            .I(N__38862));
    InMux I__8236 (
            .O(N__38872),
            .I(N__38859));
    InMux I__8235 (
            .O(N__38871),
            .I(N__38856));
    Span4Mux_v I__8234 (
            .O(N__38868),
            .I(N__38850));
    LocalMux I__8233 (
            .O(N__38865),
            .I(N__38850));
    LocalMux I__8232 (
            .O(N__38862),
            .I(N__38845));
    LocalMux I__8231 (
            .O(N__38859),
            .I(N__38845));
    LocalMux I__8230 (
            .O(N__38856),
            .I(N__38842));
    InMux I__8229 (
            .O(N__38855),
            .I(N__38839));
    Span4Mux_h I__8228 (
            .O(N__38850),
            .I(N__38836));
    Span4Mux_h I__8227 (
            .O(N__38845),
            .I(N__38833));
    Span4Mux_h I__8226 (
            .O(N__38842),
            .I(N__38828));
    LocalMux I__8225 (
            .O(N__38839),
            .I(N__38828));
    Span4Mux_h I__8224 (
            .O(N__38836),
            .I(N__38824));
    Span4Mux_h I__8223 (
            .O(N__38833),
            .I(N__38819));
    Span4Mux_h I__8222 (
            .O(N__38828),
            .I(N__38819));
    InMux I__8221 (
            .O(N__38827),
            .I(N__38816));
    Sp12to4 I__8220 (
            .O(N__38824),
            .I(N__38808));
    Sp12to4 I__8219 (
            .O(N__38819),
            .I(N__38808));
    LocalMux I__8218 (
            .O(N__38816),
            .I(N__38808));
    InMux I__8217 (
            .O(N__38815),
            .I(N__38805));
    Odrv12 I__8216 (
            .O(N__38808),
            .I(\ALU.r0_12_6 ));
    LocalMux I__8215 (
            .O(N__38805),
            .I(\ALU.r0_12_6 ));
    CascadeMux I__8214 (
            .O(N__38800),
            .I(N__38797));
    InMux I__8213 (
            .O(N__38797),
            .I(N__38794));
    LocalMux I__8212 (
            .O(N__38794),
            .I(N__38790));
    InMux I__8211 (
            .O(N__38793),
            .I(N__38787));
    Span4Mux_v I__8210 (
            .O(N__38790),
            .I(N__38783));
    LocalMux I__8209 (
            .O(N__38787),
            .I(N__38780));
    InMux I__8208 (
            .O(N__38786),
            .I(N__38777));
    Span4Mux_h I__8207 (
            .O(N__38783),
            .I(N__38774));
    Span4Mux_h I__8206 (
            .O(N__38780),
            .I(N__38771));
    LocalMux I__8205 (
            .O(N__38777),
            .I(N__38768));
    Span4Mux_v I__8204 (
            .O(N__38774),
            .I(N__38761));
    Span4Mux_v I__8203 (
            .O(N__38771),
            .I(N__38761));
    Span4Mux_h I__8202 (
            .O(N__38768),
            .I(N__38761));
    Span4Mux_h I__8201 (
            .O(N__38761),
            .I(N__38758));
    Odrv4 I__8200 (
            .O(N__38758),
            .I(r6_6));
    InMux I__8199 (
            .O(N__38755),
            .I(N__38751));
    InMux I__8198 (
            .O(N__38754),
            .I(N__38748));
    LocalMux I__8197 (
            .O(N__38751),
            .I(N__38742));
    LocalMux I__8196 (
            .O(N__38748),
            .I(N__38742));
    InMux I__8195 (
            .O(N__38747),
            .I(N__38737));
    Span4Mux_v I__8194 (
            .O(N__38742),
            .I(N__38734));
    InMux I__8193 (
            .O(N__38741),
            .I(N__38731));
    InMux I__8192 (
            .O(N__38740),
            .I(N__38728));
    LocalMux I__8191 (
            .O(N__38737),
            .I(N__38724));
    Span4Mux_h I__8190 (
            .O(N__38734),
            .I(N__38719));
    LocalMux I__8189 (
            .O(N__38731),
            .I(N__38719));
    LocalMux I__8188 (
            .O(N__38728),
            .I(N__38716));
    InMux I__8187 (
            .O(N__38727),
            .I(N__38713));
    Span4Mux_v I__8186 (
            .O(N__38724),
            .I(N__38708));
    Span4Mux_h I__8185 (
            .O(N__38719),
            .I(N__38705));
    Span12Mux_v I__8184 (
            .O(N__38716),
            .I(N__38700));
    LocalMux I__8183 (
            .O(N__38713),
            .I(N__38700));
    InMux I__8182 (
            .O(N__38712),
            .I(N__38697));
    InMux I__8181 (
            .O(N__38711),
            .I(N__38694));
    Odrv4 I__8180 (
            .O(N__38708),
            .I(\ALU.r0_12_7 ));
    Odrv4 I__8179 (
            .O(N__38705),
            .I(\ALU.r0_12_7 ));
    Odrv12 I__8178 (
            .O(N__38700),
            .I(\ALU.r0_12_7 ));
    LocalMux I__8177 (
            .O(N__38697),
            .I(\ALU.r0_12_7 ));
    LocalMux I__8176 (
            .O(N__38694),
            .I(\ALU.r0_12_7 ));
    InMux I__8175 (
            .O(N__38683),
            .I(N__38674));
    InMux I__8174 (
            .O(N__38682),
            .I(N__38674));
    InMux I__8173 (
            .O(N__38681),
            .I(N__38674));
    LocalMux I__8172 (
            .O(N__38674),
            .I(N__38671));
    Span4Mux_h I__8171 (
            .O(N__38671),
            .I(N__38668));
    Span4Mux_h I__8170 (
            .O(N__38668),
            .I(N__38665));
    Span4Mux_h I__8169 (
            .O(N__38665),
            .I(N__38662));
    Odrv4 I__8168 (
            .O(N__38662),
            .I(r6_7));
    InMux I__8167 (
            .O(N__38659),
            .I(\ALU.r0_12_4 ));
    InMux I__8166 (
            .O(N__38656),
            .I(N__38653));
    LocalMux I__8165 (
            .O(N__38653),
            .I(N__38650));
    Span4Mux_v I__8164 (
            .O(N__38650),
            .I(N__38646));
    InMux I__8163 (
            .O(N__38649),
            .I(N__38643));
    Sp12to4 I__8162 (
            .O(N__38646),
            .I(N__38640));
    LocalMux I__8161 (
            .O(N__38643),
            .I(N__38637));
    Odrv12 I__8160 (
            .O(N__38640),
            .I(\ALU.r5_RNIKS4A9Z0Z_11 ));
    Odrv4 I__8159 (
            .O(N__38637),
            .I(\ALU.r5_RNIKS4A9Z0Z_11 ));
    InMux I__8158 (
            .O(N__38632),
            .I(N__38628));
    InMux I__8157 (
            .O(N__38631),
            .I(N__38625));
    LocalMux I__8156 (
            .O(N__38628),
            .I(N__38622));
    LocalMux I__8155 (
            .O(N__38625),
            .I(\ALU.r4_RNIVLAIAZ0Z_9 ));
    Odrv4 I__8154 (
            .O(N__38622),
            .I(\ALU.r4_RNIVLAIAZ0Z_9 ));
    CascadeMux I__8153 (
            .O(N__38617),
            .I(\ALU.r5_RNI0QK3KZ0Z_11_cascade_ ));
    InMux I__8152 (
            .O(N__38614),
            .I(N__38611));
    LocalMux I__8151 (
            .O(N__38611),
            .I(N__38608));
    Span4Mux_v I__8150 (
            .O(N__38608),
            .I(N__38605));
    Odrv4 I__8149 (
            .O(N__38605),
            .I(\ALU.rshift_8 ));
    InMux I__8148 (
            .O(N__38602),
            .I(N__38599));
    LocalMux I__8147 (
            .O(N__38599),
            .I(N__38595));
    InMux I__8146 (
            .O(N__38598),
            .I(N__38592));
    Span4Mux_h I__8145 (
            .O(N__38595),
            .I(N__38589));
    LocalMux I__8144 (
            .O(N__38592),
            .I(N__38586));
    Span4Mux_v I__8143 (
            .O(N__38589),
            .I(N__38581));
    Span4Mux_v I__8142 (
            .O(N__38586),
            .I(N__38581));
    Odrv4 I__8141 (
            .O(N__38581),
            .I(\ALU.un2_addsub_cry_3_c_RNI8MVBGZ0 ));
    CascadeMux I__8140 (
            .O(N__38578),
            .I(N__38575));
    InMux I__8139 (
            .O(N__38575),
            .I(N__38572));
    LocalMux I__8138 (
            .O(N__38572),
            .I(\ALU.r0_12_prm_2_4_c_RNOZ0 ));
    InMux I__8137 (
            .O(N__38569),
            .I(N__38566));
    LocalMux I__8136 (
            .O(N__38566),
            .I(N__38563));
    Span4Mux_v I__8135 (
            .O(N__38563),
            .I(N__38560));
    Span4Mux_h I__8134 (
            .O(N__38560),
            .I(N__38556));
    InMux I__8133 (
            .O(N__38559),
            .I(N__38553));
    Odrv4 I__8132 (
            .O(N__38556),
            .I(\ALU.madd_axb_3 ));
    LocalMux I__8131 (
            .O(N__38553),
            .I(\ALU.madd_axb_3 ));
    InMux I__8130 (
            .O(N__38548),
            .I(N__38545));
    LocalMux I__8129 (
            .O(N__38545),
            .I(N__38541));
    InMux I__8128 (
            .O(N__38544),
            .I(N__38538));
    Span4Mux_h I__8127 (
            .O(N__38541),
            .I(N__38535));
    LocalMux I__8126 (
            .O(N__38538),
            .I(\ALU.madd_cry_2_THRU_CO ));
    Odrv4 I__8125 (
            .O(N__38535),
            .I(\ALU.madd_cry_2_THRU_CO ));
    InMux I__8124 (
            .O(N__38530),
            .I(N__38527));
    LocalMux I__8123 (
            .O(N__38527),
            .I(\ALU.r0_12_prm_3_4_c_RNOZ0 ));
    InMux I__8122 (
            .O(N__38524),
            .I(N__38521));
    LocalMux I__8121 (
            .O(N__38521),
            .I(N__38516));
    CascadeMux I__8120 (
            .O(N__38520),
            .I(N__38513));
    InMux I__8119 (
            .O(N__38519),
            .I(N__38510));
    Span4Mux_v I__8118 (
            .O(N__38516),
            .I(N__38507));
    InMux I__8117 (
            .O(N__38513),
            .I(N__38504));
    LocalMux I__8116 (
            .O(N__38510),
            .I(N__38501));
    Span4Mux_h I__8115 (
            .O(N__38507),
            .I(N__38498));
    LocalMux I__8114 (
            .O(N__38504),
            .I(N__38495));
    Span4Mux_v I__8113 (
            .O(N__38501),
            .I(N__38492));
    Span4Mux_h I__8112 (
            .O(N__38498),
            .I(N__38489));
    Span4Mux_h I__8111 (
            .O(N__38495),
            .I(N__38486));
    Span4Mux_h I__8110 (
            .O(N__38492),
            .I(N__38483));
    Sp12to4 I__8109 (
            .O(N__38489),
            .I(N__38480));
    Span4Mux_h I__8108 (
            .O(N__38486),
            .I(N__38477));
    Span4Mux_h I__8107 (
            .O(N__38483),
            .I(N__38474));
    Odrv12 I__8106 (
            .O(N__38480),
            .I(r1_6));
    Odrv4 I__8105 (
            .O(N__38477),
            .I(r1_6));
    Odrv4 I__8104 (
            .O(N__38474),
            .I(r1_6));
    InMux I__8103 (
            .O(N__38467),
            .I(N__38464));
    LocalMux I__8102 (
            .O(N__38464),
            .I(N__38460));
    InMux I__8101 (
            .O(N__38463),
            .I(N__38457));
    Span4Mux_h I__8100 (
            .O(N__38460),
            .I(N__38452));
    LocalMux I__8099 (
            .O(N__38457),
            .I(N__38452));
    Span4Mux_v I__8098 (
            .O(N__38452),
            .I(N__38448));
    CascadeMux I__8097 (
            .O(N__38451),
            .I(N__38445));
    Span4Mux_h I__8096 (
            .O(N__38448),
            .I(N__38442));
    InMux I__8095 (
            .O(N__38445),
            .I(N__38439));
    Odrv4 I__8094 (
            .O(N__38442),
            .I(\ALU.a4_b_4 ));
    LocalMux I__8093 (
            .O(N__38439),
            .I(\ALU.a4_b_4 ));
    CascadeMux I__8092 (
            .O(N__38434),
            .I(N__38431));
    InMux I__8091 (
            .O(N__38431),
            .I(N__38428));
    LocalMux I__8090 (
            .O(N__38428),
            .I(\ALU.r0_12_prm_7_4_c_RNOZ0 ));
    InMux I__8089 (
            .O(N__38425),
            .I(N__38422));
    LocalMux I__8088 (
            .O(N__38422),
            .I(N__38419));
    Span4Mux_v I__8087 (
            .O(N__38419),
            .I(N__38416));
    Span4Mux_h I__8086 (
            .O(N__38416),
            .I(N__38413));
    Odrv4 I__8085 (
            .O(N__38413),
            .I(\ALU.r0_12_prm_6_4_c_RNOZ0 ));
    CascadeMux I__8084 (
            .O(N__38410),
            .I(N__38407));
    InMux I__8083 (
            .O(N__38407),
            .I(N__38404));
    LocalMux I__8082 (
            .O(N__38404),
            .I(N__38401));
    Span4Mux_h I__8081 (
            .O(N__38401),
            .I(N__38398));
    Odrv4 I__8080 (
            .O(N__38398),
            .I(\ALU.un14_log_0_i_4 ));
    CascadeMux I__8079 (
            .O(N__38395),
            .I(N__38392));
    InMux I__8078 (
            .O(N__38392),
            .I(N__38389));
    LocalMux I__8077 (
            .O(N__38389),
            .I(N__38386));
    Odrv4 I__8076 (
            .O(N__38386),
            .I(\ALU.r0_12_prm_5_4_c_RNOZ0Z_0 ));
    InMux I__8075 (
            .O(N__38383),
            .I(N__38380));
    LocalMux I__8074 (
            .O(N__38380),
            .I(\ALU.a_i_4 ));
    CascadeMux I__8073 (
            .O(N__38377),
            .I(N__38374));
    InMux I__8072 (
            .O(N__38374),
            .I(N__38371));
    LocalMux I__8071 (
            .O(N__38371),
            .I(N__38368));
    Odrv12 I__8070 (
            .O(N__38368),
            .I(\ALU.mult_4 ));
    InMux I__8069 (
            .O(N__38365),
            .I(N__38362));
    LocalMux I__8068 (
            .O(N__38362),
            .I(N__38358));
    CascadeMux I__8067 (
            .O(N__38361),
            .I(N__38355));
    Span4Mux_v I__8066 (
            .O(N__38358),
            .I(N__38352));
    InMux I__8065 (
            .O(N__38355),
            .I(N__38349));
    Sp12to4 I__8064 (
            .O(N__38352),
            .I(N__38344));
    LocalMux I__8063 (
            .O(N__38349),
            .I(N__38344));
    Odrv12 I__8062 (
            .O(N__38344),
            .I(\ALU.un14_log_0_i_6 ));
    InMux I__8061 (
            .O(N__38341),
            .I(N__38337));
    CascadeMux I__8060 (
            .O(N__38340),
            .I(N__38334));
    LocalMux I__8059 (
            .O(N__38337),
            .I(N__38331));
    InMux I__8058 (
            .O(N__38334),
            .I(N__38328));
    Span4Mux_v I__8057 (
            .O(N__38331),
            .I(N__38325));
    LocalMux I__8056 (
            .O(N__38328),
            .I(N__38322));
    Odrv4 I__8055 (
            .O(N__38325),
            .I(\ALU.r4_RNI2BKQ8_0Z0Z_6 ));
    Odrv4 I__8054 (
            .O(N__38322),
            .I(\ALU.r4_RNI2BKQ8_0Z0Z_6 ));
    CascadeMux I__8053 (
            .O(N__38317),
            .I(N__38314));
    InMux I__8052 (
            .O(N__38314),
            .I(N__38311));
    LocalMux I__8051 (
            .O(N__38311),
            .I(N__38308));
    Span4Mux_h I__8050 (
            .O(N__38308),
            .I(N__38305));
    IoSpan4Mux I__8049 (
            .O(N__38305),
            .I(N__38302));
    Span4Mux_s0_v I__8048 (
            .O(N__38302),
            .I(N__38299));
    Odrv4 I__8047 (
            .O(N__38299),
            .I(\ALU.r4_RNIUGHG5Z0Z_6 ));
    CascadeMux I__8046 (
            .O(N__38296),
            .I(N__38293));
    InMux I__8045 (
            .O(N__38293),
            .I(N__38290));
    LocalMux I__8044 (
            .O(N__38290),
            .I(N__38286));
    InMux I__8043 (
            .O(N__38289),
            .I(N__38283));
    Span4Mux_s2_v I__8042 (
            .O(N__38286),
            .I(N__38280));
    LocalMux I__8041 (
            .O(N__38283),
            .I(\ALU.a_i_6 ));
    Odrv4 I__8040 (
            .O(N__38280),
            .I(\ALU.a_i_6 ));
    CascadeMux I__8039 (
            .O(N__38275),
            .I(N__38272));
    InMux I__8038 (
            .O(N__38272),
            .I(N__38269));
    LocalMux I__8037 (
            .O(N__38269),
            .I(\ALU.r0_12_prm_3_6_s0_sf ));
    InMux I__8036 (
            .O(N__38266),
            .I(N__38262));
    InMux I__8035 (
            .O(N__38265),
            .I(N__38259));
    LocalMux I__8034 (
            .O(N__38262),
            .I(N__38254));
    LocalMux I__8033 (
            .O(N__38259),
            .I(N__38251));
    InMux I__8032 (
            .O(N__38258),
            .I(N__38248));
    InMux I__8031 (
            .O(N__38257),
            .I(N__38245));
    Span4Mux_s1_v I__8030 (
            .O(N__38254),
            .I(N__38242));
    Span4Mux_h I__8029 (
            .O(N__38251),
            .I(N__38239));
    LocalMux I__8028 (
            .O(N__38248),
            .I(N__38236));
    LocalMux I__8027 (
            .O(N__38245),
            .I(N__38233));
    Span4Mux_v I__8026 (
            .O(N__38242),
            .I(N__38230));
    Span4Mux_v I__8025 (
            .O(N__38239),
            .I(N__38227));
    Span12Mux_h I__8024 (
            .O(N__38236),
            .I(N__38222));
    Span12Mux_s2_v I__8023 (
            .O(N__38233),
            .I(N__38222));
    Odrv4 I__8022 (
            .O(N__38230),
            .I(\ALU.un2_addsub_cry_5_c_RNIO30SDZ0 ));
    Odrv4 I__8021 (
            .O(N__38227),
            .I(\ALU.un2_addsub_cry_5_c_RNIO30SDZ0 ));
    Odrv12 I__8020 (
            .O(N__38222),
            .I(\ALU.un2_addsub_cry_5_c_RNIO30SDZ0 ));
    CascadeMux I__8019 (
            .O(N__38215),
            .I(N__38212));
    InMux I__8018 (
            .O(N__38212),
            .I(N__38209));
    LocalMux I__8017 (
            .O(N__38209),
            .I(\ALU.r0_12_prm_2_6_s0_c_RNOZ0 ));
    InMux I__8016 (
            .O(N__38206),
            .I(N__38201));
    InMux I__8015 (
            .O(N__38205),
            .I(N__38198));
    InMux I__8014 (
            .O(N__38204),
            .I(N__38195));
    LocalMux I__8013 (
            .O(N__38201),
            .I(N__38192));
    LocalMux I__8012 (
            .O(N__38198),
            .I(N__38189));
    LocalMux I__8011 (
            .O(N__38195),
            .I(N__38186));
    Span4Mux_s0_v I__8010 (
            .O(N__38192),
            .I(N__38182));
    Span12Mux_s7_v I__8009 (
            .O(N__38189),
            .I(N__38179));
    Span4Mux_v I__8008 (
            .O(N__38186),
            .I(N__38176));
    InMux I__8007 (
            .O(N__38185),
            .I(N__38173));
    Span4Mux_v I__8006 (
            .O(N__38182),
            .I(N__38170));
    Odrv12 I__8005 (
            .O(N__38179),
            .I(\ALU.un9_addsub_cry_5_c_RNI3CZ0Z019 ));
    Odrv4 I__8004 (
            .O(N__38176),
            .I(\ALU.un9_addsub_cry_5_c_RNI3CZ0Z019 ));
    LocalMux I__8003 (
            .O(N__38173),
            .I(\ALU.un9_addsub_cry_5_c_RNI3CZ0Z019 ));
    Odrv4 I__8002 (
            .O(N__38170),
            .I(\ALU.un9_addsub_cry_5_c_RNI3CZ0Z019 ));
    CascadeMux I__8001 (
            .O(N__38161),
            .I(N__38158));
    InMux I__8000 (
            .O(N__38158),
            .I(N__38155));
    LocalMux I__7999 (
            .O(N__38155),
            .I(N__38152));
    Span4Mux_v I__7998 (
            .O(N__38152),
            .I(N__38149));
    Odrv4 I__7997 (
            .O(N__38149),
            .I(\ALU.r0_12_prm_1_6_s0_c_RNOZ0 ));
    InMux I__7996 (
            .O(N__38146),
            .I(N__38143));
    LocalMux I__7995 (
            .O(N__38143),
            .I(N__38140));
    Span4Mux_h I__7994 (
            .O(N__38140),
            .I(N__38137));
    Odrv4 I__7993 (
            .O(N__38137),
            .I(\ALU.r0_12_s1_6_THRU_CO ));
    InMux I__7992 (
            .O(N__38134),
            .I(N__38131));
    LocalMux I__7991 (
            .O(N__38131),
            .I(N__38128));
    Span4Mux_h I__7990 (
            .O(N__38128),
            .I(N__38125));
    Span4Mux_h I__7989 (
            .O(N__38125),
            .I(N__38122));
    Odrv4 I__7988 (
            .O(N__38122),
            .I(\ALU.mult_6 ));
    InMux I__7987 (
            .O(N__38119),
            .I(\ALU.r0_12_s0_6 ));
    InMux I__7986 (
            .O(N__38116),
            .I(N__38113));
    LocalMux I__7985 (
            .O(N__38113),
            .I(\ALU.r0_12_prm_2_0_s1_c_RNOZ0 ));
    InMux I__7984 (
            .O(N__38110),
            .I(N__38107));
    LocalMux I__7983 (
            .O(N__38107),
            .I(N__38104));
    Span4Mux_h I__7982 (
            .O(N__38104),
            .I(N__38101));
    Odrv4 I__7981 (
            .O(N__38101),
            .I(\ALU.r0_12_prm_8_2_c_RNOZ0Z_3 ));
    InMux I__7980 (
            .O(N__38098),
            .I(N__38095));
    LocalMux I__7979 (
            .O(N__38095),
            .I(N__38092));
    Span4Mux_h I__7978 (
            .O(N__38092),
            .I(N__38089));
    Span4Mux_s1_v I__7977 (
            .O(N__38089),
            .I(N__38086));
    Odrv4 I__7976 (
            .O(N__38086),
            .I(\ALU.r4_RNI1G9PKZ0Z_6 ));
    InMux I__7975 (
            .O(N__38083),
            .I(N__38080));
    LocalMux I__7974 (
            .O(N__38080),
            .I(N__38077));
    Span4Mux_s3_v I__7973 (
            .O(N__38077),
            .I(N__38072));
    InMux I__7972 (
            .O(N__38076),
            .I(N__38067));
    InMux I__7971 (
            .O(N__38075),
            .I(N__38067));
    Odrv4 I__7970 (
            .O(N__38072),
            .I(\ALU.N_845_1 ));
    LocalMux I__7969 (
            .O(N__38067),
            .I(\ALU.N_845_1 ));
    CascadeMux I__7968 (
            .O(N__38062),
            .I(\ALU.rshift_15_ns_1_2_cascade_ ));
    InMux I__7967 (
            .O(N__38059),
            .I(N__38056));
    LocalMux I__7966 (
            .O(N__38056),
            .I(N__38053));
    Span4Mux_h I__7965 (
            .O(N__38053),
            .I(N__38047));
    InMux I__7964 (
            .O(N__38052),
            .I(N__38044));
    InMux I__7963 (
            .O(N__38051),
            .I(N__38039));
    InMux I__7962 (
            .O(N__38050),
            .I(N__38039));
    Odrv4 I__7961 (
            .O(N__38047),
            .I(\ALU.r5_RNI8R2TIZ0Z_11 ));
    LocalMux I__7960 (
            .O(N__38044),
            .I(\ALU.r5_RNI8R2TIZ0Z_11 ));
    LocalMux I__7959 (
            .O(N__38039),
            .I(\ALU.r5_RNI8R2TIZ0Z_11 ));
    InMux I__7958 (
            .O(N__38032),
            .I(N__38022));
    InMux I__7957 (
            .O(N__38031),
            .I(N__38012));
    InMux I__7956 (
            .O(N__38030),
            .I(N__38009));
    InMux I__7955 (
            .O(N__38029),
            .I(N__38002));
    InMux I__7954 (
            .O(N__38028),
            .I(N__38002));
    InMux I__7953 (
            .O(N__38027),
            .I(N__37995));
    InMux I__7952 (
            .O(N__38026),
            .I(N__37995));
    InMux I__7951 (
            .O(N__38025),
            .I(N__37995));
    LocalMux I__7950 (
            .O(N__38022),
            .I(N__37989));
    InMux I__7949 (
            .O(N__38021),
            .I(N__37985));
    InMux I__7948 (
            .O(N__38020),
            .I(N__37982));
    InMux I__7947 (
            .O(N__38019),
            .I(N__37977));
    InMux I__7946 (
            .O(N__38018),
            .I(N__37977));
    InMux I__7945 (
            .O(N__38017),
            .I(N__37974));
    InMux I__7944 (
            .O(N__38016),
            .I(N__37970));
    InMux I__7943 (
            .O(N__38015),
            .I(N__37961));
    LocalMux I__7942 (
            .O(N__38012),
            .I(N__37955));
    LocalMux I__7941 (
            .O(N__38009),
            .I(N__37955));
    InMux I__7940 (
            .O(N__38008),
            .I(N__37950));
    InMux I__7939 (
            .O(N__38007),
            .I(N__37950));
    LocalMux I__7938 (
            .O(N__38002),
            .I(N__37945));
    LocalMux I__7937 (
            .O(N__37995),
            .I(N__37945));
    InMux I__7936 (
            .O(N__37994),
            .I(N__37938));
    InMux I__7935 (
            .O(N__37993),
            .I(N__37938));
    InMux I__7934 (
            .O(N__37992),
            .I(N__37938));
    Span4Mux_s3_v I__7933 (
            .O(N__37989),
            .I(N__37935));
    InMux I__7932 (
            .O(N__37988),
            .I(N__37932));
    LocalMux I__7931 (
            .O(N__37985),
            .I(N__37929));
    LocalMux I__7930 (
            .O(N__37982),
            .I(N__37924));
    LocalMux I__7929 (
            .O(N__37977),
            .I(N__37924));
    LocalMux I__7928 (
            .O(N__37974),
            .I(N__37921));
    InMux I__7927 (
            .O(N__37973),
            .I(N__37918));
    LocalMux I__7926 (
            .O(N__37970),
            .I(N__37915));
    InMux I__7925 (
            .O(N__37969),
            .I(N__37908));
    InMux I__7924 (
            .O(N__37968),
            .I(N__37908));
    InMux I__7923 (
            .O(N__37967),
            .I(N__37908));
    InMux I__7922 (
            .O(N__37966),
            .I(N__37903));
    InMux I__7921 (
            .O(N__37965),
            .I(N__37903));
    InMux I__7920 (
            .O(N__37964),
            .I(N__37900));
    LocalMux I__7919 (
            .O(N__37961),
            .I(N__37892));
    InMux I__7918 (
            .O(N__37960),
            .I(N__37889));
    Span4Mux_h I__7917 (
            .O(N__37955),
            .I(N__37875));
    LocalMux I__7916 (
            .O(N__37950),
            .I(N__37875));
    Span4Mux_v I__7915 (
            .O(N__37945),
            .I(N__37875));
    LocalMux I__7914 (
            .O(N__37938),
            .I(N__37875));
    Span4Mux_h I__7913 (
            .O(N__37935),
            .I(N__37870));
    LocalMux I__7912 (
            .O(N__37932),
            .I(N__37870));
    Span4Mux_v I__7911 (
            .O(N__37929),
            .I(N__37867));
    Span4Mux_s3_v I__7910 (
            .O(N__37924),
            .I(N__37860));
    Span4Mux_s1_h I__7909 (
            .O(N__37921),
            .I(N__37860));
    LocalMux I__7908 (
            .O(N__37918),
            .I(N__37860));
    Span4Mux_h I__7907 (
            .O(N__37915),
            .I(N__37855));
    LocalMux I__7906 (
            .O(N__37908),
            .I(N__37855));
    LocalMux I__7905 (
            .O(N__37903),
            .I(N__37852));
    LocalMux I__7904 (
            .O(N__37900),
            .I(N__37849));
    InMux I__7903 (
            .O(N__37899),
            .I(N__37842));
    InMux I__7902 (
            .O(N__37898),
            .I(N__37842));
    InMux I__7901 (
            .O(N__37897),
            .I(N__37842));
    InMux I__7900 (
            .O(N__37896),
            .I(N__37837));
    InMux I__7899 (
            .O(N__37895),
            .I(N__37837));
    Sp12to4 I__7898 (
            .O(N__37892),
            .I(N__37832));
    LocalMux I__7897 (
            .O(N__37889),
            .I(N__37832));
    InMux I__7896 (
            .O(N__37888),
            .I(N__37823));
    InMux I__7895 (
            .O(N__37887),
            .I(N__37814));
    InMux I__7894 (
            .O(N__37886),
            .I(N__37814));
    InMux I__7893 (
            .O(N__37885),
            .I(N__37814));
    InMux I__7892 (
            .O(N__37884),
            .I(N__37814));
    Span4Mux_h I__7891 (
            .O(N__37875),
            .I(N__37811));
    Span4Mux_h I__7890 (
            .O(N__37870),
            .I(N__37804));
    Span4Mux_h I__7889 (
            .O(N__37867),
            .I(N__37804));
    Span4Mux_h I__7888 (
            .O(N__37860),
            .I(N__37804));
    Span4Mux_h I__7887 (
            .O(N__37855),
            .I(N__37799));
    Span4Mux_h I__7886 (
            .O(N__37852),
            .I(N__37799));
    Span4Mux_h I__7885 (
            .O(N__37849),
            .I(N__37794));
    LocalMux I__7884 (
            .O(N__37842),
            .I(N__37794));
    LocalMux I__7883 (
            .O(N__37837),
            .I(N__37789));
    Span12Mux_v I__7882 (
            .O(N__37832),
            .I(N__37789));
    InMux I__7881 (
            .O(N__37831),
            .I(N__37784));
    InMux I__7880 (
            .O(N__37830),
            .I(N__37784));
    InMux I__7879 (
            .O(N__37829),
            .I(N__37775));
    InMux I__7878 (
            .O(N__37828),
            .I(N__37775));
    InMux I__7877 (
            .O(N__37827),
            .I(N__37775));
    InMux I__7876 (
            .O(N__37826),
            .I(N__37775));
    LocalMux I__7875 (
            .O(N__37823),
            .I(\ALU.bZ0Z_0 ));
    LocalMux I__7874 (
            .O(N__37814),
            .I(\ALU.bZ0Z_0 ));
    Odrv4 I__7873 (
            .O(N__37811),
            .I(\ALU.bZ0Z_0 ));
    Odrv4 I__7872 (
            .O(N__37804),
            .I(\ALU.bZ0Z_0 ));
    Odrv4 I__7871 (
            .O(N__37799),
            .I(\ALU.bZ0Z_0 ));
    Odrv4 I__7870 (
            .O(N__37794),
            .I(\ALU.bZ0Z_0 ));
    Odrv12 I__7869 (
            .O(N__37789),
            .I(\ALU.bZ0Z_0 ));
    LocalMux I__7868 (
            .O(N__37784),
            .I(\ALU.bZ0Z_0 ));
    LocalMux I__7867 (
            .O(N__37775),
            .I(\ALU.bZ0Z_0 ));
    InMux I__7866 (
            .O(N__37756),
            .I(N__37753));
    LocalMux I__7865 (
            .O(N__37753),
            .I(N__37749));
    CascadeMux I__7864 (
            .O(N__37752),
            .I(N__37746));
    Span4Mux_h I__7863 (
            .O(N__37749),
            .I(N__37743));
    InMux I__7862 (
            .O(N__37746),
            .I(N__37740));
    Odrv4 I__7861 (
            .O(N__37743),
            .I(\ALU.r4_RNID26E8_0Z0Z_0 ));
    LocalMux I__7860 (
            .O(N__37740),
            .I(\ALU.r4_RNID26E8_0Z0Z_0 ));
    CascadeMux I__7859 (
            .O(N__37735),
            .I(N__37731));
    CascadeMux I__7858 (
            .O(N__37734),
            .I(N__37727));
    InMux I__7857 (
            .O(N__37731),
            .I(N__37723));
    InMux I__7856 (
            .O(N__37730),
            .I(N__37720));
    InMux I__7855 (
            .O(N__37727),
            .I(N__37717));
    InMux I__7854 (
            .O(N__37726),
            .I(N__37714));
    LocalMux I__7853 (
            .O(N__37723),
            .I(N__37709));
    LocalMux I__7852 (
            .O(N__37720),
            .I(N__37709));
    LocalMux I__7851 (
            .O(N__37717),
            .I(N__37704));
    LocalMux I__7850 (
            .O(N__37714),
            .I(N__37704));
    Span4Mux_h I__7849 (
            .O(N__37709),
            .I(N__37701));
    Span4Mux_s0_v I__7848 (
            .O(N__37704),
            .I(N__37698));
    Odrv4 I__7847 (
            .O(N__37701),
            .I(\ALU.rshift_6 ));
    Odrv4 I__7846 (
            .O(N__37698),
            .I(\ALU.rshift_6 ));
    InMux I__7845 (
            .O(N__37693),
            .I(N__37690));
    LocalMux I__7844 (
            .O(N__37690),
            .I(N__37685));
    CascadeMux I__7843 (
            .O(N__37689),
            .I(N__37682));
    InMux I__7842 (
            .O(N__37688),
            .I(N__37679));
    Span4Mux_h I__7841 (
            .O(N__37685),
            .I(N__37676));
    InMux I__7840 (
            .O(N__37682),
            .I(N__37673));
    LocalMux I__7839 (
            .O(N__37679),
            .I(N__37670));
    Odrv4 I__7838 (
            .O(N__37676),
            .I(\ALU.lshift_6 ));
    LocalMux I__7837 (
            .O(N__37673),
            .I(\ALU.lshift_6 ));
    Odrv4 I__7836 (
            .O(N__37670),
            .I(\ALU.lshift_6 ));
    CascadeMux I__7835 (
            .O(N__37663),
            .I(N__37660));
    InMux I__7834 (
            .O(N__37660),
            .I(N__37657));
    LocalMux I__7833 (
            .O(N__37657),
            .I(\ALU.r0_12_prm_8_6_s0_c_RNOZ0 ));
    InMux I__7832 (
            .O(N__37654),
            .I(N__37651));
    LocalMux I__7831 (
            .O(N__37651),
            .I(N__37647));
    InMux I__7830 (
            .O(N__37650),
            .I(N__37644));
    Span4Mux_v I__7829 (
            .O(N__37647),
            .I(N__37641));
    LocalMux I__7828 (
            .O(N__37644),
            .I(N__37638));
    Span4Mux_h I__7827 (
            .O(N__37641),
            .I(N__37633));
    Span4Mux_h I__7826 (
            .O(N__37638),
            .I(N__37630));
    InMux I__7825 (
            .O(N__37637),
            .I(N__37627));
    InMux I__7824 (
            .O(N__37636),
            .I(N__37624));
    Odrv4 I__7823 (
            .O(N__37633),
            .I(\ALU.un2_addsub_cry_11_c_RNICP8AEZ0 ));
    Odrv4 I__7822 (
            .O(N__37630),
            .I(\ALU.un2_addsub_cry_11_c_RNICP8AEZ0 ));
    LocalMux I__7821 (
            .O(N__37627),
            .I(\ALU.un2_addsub_cry_11_c_RNICP8AEZ0 ));
    LocalMux I__7820 (
            .O(N__37624),
            .I(\ALU.un2_addsub_cry_11_c_RNICP8AEZ0 ));
    CascadeMux I__7819 (
            .O(N__37615),
            .I(N__37612));
    InMux I__7818 (
            .O(N__37612),
            .I(N__37609));
    LocalMux I__7817 (
            .O(N__37609),
            .I(N__37606));
    Odrv4 I__7816 (
            .O(N__37606),
            .I(\ALU.r0_12_prm_2_12_s1_c_RNOZ0 ));
    InMux I__7815 (
            .O(N__37603),
            .I(N__37600));
    LocalMux I__7814 (
            .O(N__37600),
            .I(N__37597));
    Odrv4 I__7813 (
            .O(N__37597),
            .I(\ALU.r0_12_prm_1_12_s1_c_RNOZ0 ));
    InMux I__7812 (
            .O(N__37594),
            .I(N__37590));
    CascadeMux I__7811 (
            .O(N__37593),
            .I(N__37587));
    LocalMux I__7810 (
            .O(N__37590),
            .I(N__37583));
    InMux I__7809 (
            .O(N__37587),
            .I(N__37580));
    InMux I__7808 (
            .O(N__37586),
            .I(N__37577));
    Span4Mux_v I__7807 (
            .O(N__37583),
            .I(N__37573));
    LocalMux I__7806 (
            .O(N__37580),
            .I(N__37568));
    LocalMux I__7805 (
            .O(N__37577),
            .I(N__37568));
    InMux I__7804 (
            .O(N__37576),
            .I(N__37565));
    Span4Mux_h I__7803 (
            .O(N__37573),
            .I(N__37558));
    Span4Mux_v I__7802 (
            .O(N__37568),
            .I(N__37558));
    LocalMux I__7801 (
            .O(N__37565),
            .I(N__37558));
    Odrv4 I__7800 (
            .O(N__37558),
            .I(\ALU.un9_addsub_cry_11_c_RNIAHI1AZ0 ));
    InMux I__7799 (
            .O(N__37555),
            .I(\ALU.r0_12_s1_12 ));
    InMux I__7798 (
            .O(N__37552),
            .I(N__37549));
    LocalMux I__7797 (
            .O(N__37549),
            .I(N__37546));
    Span12Mux_v I__7796 (
            .O(N__37546),
            .I(N__37543));
    Odrv12 I__7795 (
            .O(N__37543),
            .I(\ALU.r0_12_s1_12_THRU_CO ));
    CascadeMux I__7794 (
            .O(N__37540),
            .I(N__37537));
    InMux I__7793 (
            .O(N__37537),
            .I(N__37534));
    LocalMux I__7792 (
            .O(N__37534),
            .I(N__37531));
    Span4Mux_v I__7791 (
            .O(N__37531),
            .I(N__37528));
    Span4Mux_h I__7790 (
            .O(N__37528),
            .I(N__37525));
    Span4Mux_h I__7789 (
            .O(N__37525),
            .I(N__37522));
    Odrv4 I__7788 (
            .O(N__37522),
            .I(\ALU.r0_12_prm_5_15_s1_c_RNOZ0 ));
    InMux I__7787 (
            .O(N__37519),
            .I(N__37516));
    LocalMux I__7786 (
            .O(N__37516),
            .I(N__37513));
    Span12Mux_s7_h I__7785 (
            .O(N__37513),
            .I(N__37510));
    Span12Mux_v I__7784 (
            .O(N__37510),
            .I(N__37507));
    Odrv12 I__7783 (
            .O(N__37507),
            .I(\ALU.r0_12_prm_8_15_s1_c_RNOZ0Z_1 ));
    InMux I__7782 (
            .O(N__37504),
            .I(N__37501));
    LocalMux I__7781 (
            .O(N__37501),
            .I(\ALU.r0_12_prm_8_0_s1_c_RNOZ0 ));
    InMux I__7780 (
            .O(N__37498),
            .I(N__37495));
    LocalMux I__7779 (
            .O(N__37495),
            .I(N__37492));
    Span4Mux_h I__7778 (
            .O(N__37492),
            .I(N__37489));
    Odrv4 I__7777 (
            .O(N__37489),
            .I(\ALU.r5_RNIAV175Z0Z_15 ));
    InMux I__7776 (
            .O(N__37486),
            .I(N__37482));
    InMux I__7775 (
            .O(N__37485),
            .I(N__37479));
    LocalMux I__7774 (
            .O(N__37482),
            .I(\ALU.r4_RNIQK1V71Z0Z_5 ));
    LocalMux I__7773 (
            .O(N__37479),
            .I(\ALU.r4_RNIQK1V71Z0Z_5 ));
    InMux I__7772 (
            .O(N__37474),
            .I(N__37471));
    LocalMux I__7771 (
            .O(N__37471),
            .I(\ALU.r0_12_prm_8_12_s1_c_RNOZ0 ));
    InMux I__7770 (
            .O(N__37468),
            .I(N__37465));
    LocalMux I__7769 (
            .O(N__37465),
            .I(N__37461));
    CascadeMux I__7768 (
            .O(N__37464),
            .I(N__37458));
    Span4Mux_h I__7767 (
            .O(N__37461),
            .I(N__37455));
    InMux I__7766 (
            .O(N__37458),
            .I(N__37452));
    Odrv4 I__7765 (
            .O(N__37455),
            .I(\ALU.lshift_12 ));
    LocalMux I__7764 (
            .O(N__37452),
            .I(\ALU.lshift_12 ));
    InMux I__7763 (
            .O(N__37447),
            .I(N__37444));
    LocalMux I__7762 (
            .O(N__37444),
            .I(\ALU.r0_12_prm_7_12_s1_c_RNOZ0 ));
    CascadeMux I__7761 (
            .O(N__37441),
            .I(N__37438));
    InMux I__7760 (
            .O(N__37438),
            .I(N__37434));
    InMux I__7759 (
            .O(N__37437),
            .I(N__37431));
    LocalMux I__7758 (
            .O(N__37434),
            .I(N__37428));
    LocalMux I__7757 (
            .O(N__37431),
            .I(N__37425));
    Span4Mux_v I__7756 (
            .O(N__37428),
            .I(N__37422));
    Span4Mux_v I__7755 (
            .O(N__37425),
            .I(N__37417));
    Span4Mux_h I__7754 (
            .O(N__37422),
            .I(N__37417));
    Odrv4 I__7753 (
            .O(N__37417),
            .I(\ALU.r5_RNISP2L9_0Z0Z_12 ));
    InMux I__7752 (
            .O(N__37414),
            .I(N__37411));
    LocalMux I__7751 (
            .O(N__37411),
            .I(N__37407));
    InMux I__7750 (
            .O(N__37410),
            .I(N__37404));
    Span4Mux_h I__7749 (
            .O(N__37407),
            .I(N__37401));
    LocalMux I__7748 (
            .O(N__37404),
            .I(N__37398));
    Sp12to4 I__7747 (
            .O(N__37401),
            .I(N__37395));
    Span4Mux_h I__7746 (
            .O(N__37398),
            .I(N__37392));
    Span12Mux_v I__7745 (
            .O(N__37395),
            .I(N__37389));
    Odrv4 I__7744 (
            .O(N__37392),
            .I(\ALU.un14_log_0_i_12 ));
    Odrv12 I__7743 (
            .O(N__37389),
            .I(\ALU.un14_log_0_i_12 ));
    InMux I__7742 (
            .O(N__37384),
            .I(N__37381));
    LocalMux I__7741 (
            .O(N__37381),
            .I(N__37378));
    Span4Mux_h I__7740 (
            .O(N__37378),
            .I(N__37375));
    Span4Mux_v I__7739 (
            .O(N__37375),
            .I(N__37372));
    Odrv4 I__7738 (
            .O(N__37372),
            .I(\ALU.r0_12_prm_5_12_s1_c_RNOZ0 ));
    InMux I__7737 (
            .O(N__37369),
            .I(N__37366));
    LocalMux I__7736 (
            .O(N__37366),
            .I(N__37363));
    Span4Mux_h I__7735 (
            .O(N__37363),
            .I(N__37359));
    CascadeMux I__7734 (
            .O(N__37362),
            .I(N__37356));
    Span4Mux_h I__7733 (
            .O(N__37359),
            .I(N__37353));
    InMux I__7732 (
            .O(N__37356),
            .I(N__37350));
    Odrv4 I__7731 (
            .O(N__37353),
            .I(\ALU.r5_RNISP2L9_1Z0Z_12 ));
    LocalMux I__7730 (
            .O(N__37350),
            .I(\ALU.r5_RNISP2L9_1Z0Z_12 ));
    InMux I__7729 (
            .O(N__37345),
            .I(N__37342));
    LocalMux I__7728 (
            .O(N__37342),
            .I(N__37339));
    Span4Mux_v I__7727 (
            .O(N__37339),
            .I(N__37336));
    Odrv4 I__7726 (
            .O(N__37336),
            .I(\ALU.r0_12_prm_4_12_s1_c_RNOZ0 ));
    CascadeMux I__7725 (
            .O(N__37333),
            .I(N__37330));
    InMux I__7724 (
            .O(N__37330),
            .I(N__37327));
    LocalMux I__7723 (
            .O(N__37327),
            .I(N__37324));
    Span4Mux_h I__7722 (
            .O(N__37324),
            .I(N__37320));
    InMux I__7721 (
            .O(N__37323),
            .I(N__37317));
    Span4Mux_h I__7720 (
            .O(N__37320),
            .I(N__37314));
    LocalMux I__7719 (
            .O(N__37317),
            .I(\ALU.a_i_12 ));
    Odrv4 I__7718 (
            .O(N__37314),
            .I(\ALU.a_i_12 ));
    InMux I__7717 (
            .O(N__37309),
            .I(\ALU.r0_12_s0_8 ));
    CascadeMux I__7716 (
            .O(N__37306),
            .I(N__37303));
    InMux I__7715 (
            .O(N__37303),
            .I(N__37300));
    LocalMux I__7714 (
            .O(N__37300),
            .I(\ALU.r0_12_prm_1_8_s0_c_RNOZ0 ));
    InMux I__7713 (
            .O(N__37297),
            .I(N__37294));
    LocalMux I__7712 (
            .O(N__37294),
            .I(N__37291));
    Span4Mux_h I__7711 (
            .O(N__37291),
            .I(N__37287));
    CascadeMux I__7710 (
            .O(N__37290),
            .I(N__37284));
    Span4Mux_h I__7709 (
            .O(N__37287),
            .I(N__37280));
    InMux I__7708 (
            .O(N__37284),
            .I(N__37277));
    InMux I__7707 (
            .O(N__37283),
            .I(N__37274));
    Span4Mux_v I__7706 (
            .O(N__37280),
            .I(N__37270));
    LocalMux I__7705 (
            .O(N__37277),
            .I(N__37267));
    LocalMux I__7704 (
            .O(N__37274),
            .I(N__37264));
    InMux I__7703 (
            .O(N__37273),
            .I(N__37261));
    Odrv4 I__7702 (
            .O(N__37270),
            .I(\ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9 ));
    Odrv12 I__7701 (
            .O(N__37267),
            .I(\ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9 ));
    Odrv4 I__7700 (
            .O(N__37264),
            .I(\ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9 ));
    LocalMux I__7699 (
            .O(N__37261),
            .I(\ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9 ));
    CascadeMux I__7698 (
            .O(N__37252),
            .I(N__37249));
    InMux I__7697 (
            .O(N__37249),
            .I(N__37246));
    LocalMux I__7696 (
            .O(N__37246),
            .I(N__37243));
    Span4Mux_h I__7695 (
            .O(N__37243),
            .I(N__37240));
    Span4Mux_h I__7694 (
            .O(N__37240),
            .I(N__37237));
    Odrv4 I__7693 (
            .O(N__37237),
            .I(\ALU.r0_12_prm_1_15_s1_c_RNOZ0 ));
    InMux I__7692 (
            .O(N__37234),
            .I(N__37231));
    LocalMux I__7691 (
            .O(N__37231),
            .I(N__37228));
    Span4Mux_h I__7690 (
            .O(N__37228),
            .I(N__37225));
    Span4Mux_h I__7689 (
            .O(N__37225),
            .I(N__37222));
    Odrv4 I__7688 (
            .O(N__37222),
            .I(\ALU.mult_5 ));
    InMux I__7687 (
            .O(N__37219),
            .I(\ALU.r0_12_s0_5 ));
    InMux I__7686 (
            .O(N__37216),
            .I(N__37213));
    LocalMux I__7685 (
            .O(N__37213),
            .I(N__37205));
    InMux I__7684 (
            .O(N__37212),
            .I(N__37202));
    InMux I__7683 (
            .O(N__37211),
            .I(N__37199));
    InMux I__7682 (
            .O(N__37210),
            .I(N__37196));
    InMux I__7681 (
            .O(N__37209),
            .I(N__37193));
    InMux I__7680 (
            .O(N__37208),
            .I(N__37190));
    Span4Mux_v I__7679 (
            .O(N__37205),
            .I(N__37180));
    LocalMux I__7678 (
            .O(N__37202),
            .I(N__37180));
    LocalMux I__7677 (
            .O(N__37199),
            .I(N__37180));
    LocalMux I__7676 (
            .O(N__37196),
            .I(N__37180));
    LocalMux I__7675 (
            .O(N__37193),
            .I(N__37177));
    LocalMux I__7674 (
            .O(N__37190),
            .I(N__37174));
    InMux I__7673 (
            .O(N__37189),
            .I(N__37171));
    Span4Mux_v I__7672 (
            .O(N__37180),
            .I(N__37168));
    Span4Mux_h I__7671 (
            .O(N__37177),
            .I(N__37165));
    Span4Mux_v I__7670 (
            .O(N__37174),
            .I(N__37160));
    LocalMux I__7669 (
            .O(N__37171),
            .I(N__37160));
    Span4Mux_h I__7668 (
            .O(N__37168),
            .I(N__37157));
    Span4Mux_h I__7667 (
            .O(N__37165),
            .I(N__37154));
    Span4Mux_v I__7666 (
            .O(N__37160),
            .I(N__37151));
    Span4Mux_h I__7665 (
            .O(N__37157),
            .I(N__37147));
    Span4Mux_h I__7664 (
            .O(N__37154),
            .I(N__37144));
    Span4Mux_h I__7663 (
            .O(N__37151),
            .I(N__37141));
    InMux I__7662 (
            .O(N__37150),
            .I(N__37138));
    Odrv4 I__7661 (
            .O(N__37147),
            .I(\ALU.r0_12_5 ));
    Odrv4 I__7660 (
            .O(N__37144),
            .I(\ALU.r0_12_5 ));
    Odrv4 I__7659 (
            .O(N__37141),
            .I(\ALU.r0_12_5 ));
    LocalMux I__7658 (
            .O(N__37138),
            .I(\ALU.r0_12_5 ));
    CascadeMux I__7657 (
            .O(N__37129),
            .I(N__37126));
    InMux I__7656 (
            .O(N__37126),
            .I(N__37121));
    InMux I__7655 (
            .O(N__37125),
            .I(N__37118));
    CascadeMux I__7654 (
            .O(N__37124),
            .I(N__37115));
    LocalMux I__7653 (
            .O(N__37121),
            .I(N__37112));
    LocalMux I__7652 (
            .O(N__37118),
            .I(N__37109));
    InMux I__7651 (
            .O(N__37115),
            .I(N__37106));
    Span4Mux_v I__7650 (
            .O(N__37112),
            .I(N__37103));
    Sp12to4 I__7649 (
            .O(N__37109),
            .I(N__37100));
    LocalMux I__7648 (
            .O(N__37106),
            .I(N__37097));
    Span4Mux_h I__7647 (
            .O(N__37103),
            .I(N__37094));
    Span12Mux_v I__7646 (
            .O(N__37100),
            .I(N__37089));
    Span12Mux_s5_h I__7645 (
            .O(N__37097),
            .I(N__37089));
    Odrv4 I__7644 (
            .O(N__37094),
            .I(r1_5));
    Odrv12 I__7643 (
            .O(N__37089),
            .I(r1_5));
    InMux I__7642 (
            .O(N__37084),
            .I(N__37081));
    LocalMux I__7641 (
            .O(N__37081),
            .I(N__37078));
    Span4Mux_v I__7640 (
            .O(N__37078),
            .I(N__37075));
    Span4Mux_v I__7639 (
            .O(N__37075),
            .I(N__37072));
    Span4Mux_h I__7638 (
            .O(N__37072),
            .I(N__37069));
    Odrv4 I__7637 (
            .O(N__37069),
            .I(\ALU.r0_12_prm_6_8_s0_c_RNOZ0 ));
    InMux I__7636 (
            .O(N__37066),
            .I(N__37063));
    LocalMux I__7635 (
            .O(N__37063),
            .I(\ALU.r0_12_prm_3_8_s0_sf ));
    CascadeMux I__7634 (
            .O(N__37060),
            .I(N__37057));
    InMux I__7633 (
            .O(N__37057),
            .I(N__37054));
    LocalMux I__7632 (
            .O(N__37054),
            .I(N__37051));
    Span4Mux_v I__7631 (
            .O(N__37051),
            .I(N__37048));
    Sp12to4 I__7630 (
            .O(N__37048),
            .I(N__37045));
    Odrv12 I__7629 (
            .O(N__37045),
            .I(\ALU.r0_12_prm_7_5_s0_c_RNOZ0 ));
    CascadeMux I__7628 (
            .O(N__37042),
            .I(N__37039));
    InMux I__7627 (
            .O(N__37039),
            .I(N__37036));
    LocalMux I__7626 (
            .O(N__37036),
            .I(N__37033));
    Span4Mux_v I__7625 (
            .O(N__37033),
            .I(N__37030));
    Span4Mux_h I__7624 (
            .O(N__37030),
            .I(N__37027));
    Odrv4 I__7623 (
            .O(N__37027),
            .I(\ALU.r0_12_prm_6_5_s0_c_RNOZ0 ));
    CascadeMux I__7622 (
            .O(N__37024),
            .I(N__37021));
    InMux I__7621 (
            .O(N__37021),
            .I(N__37018));
    LocalMux I__7620 (
            .O(N__37018),
            .I(N__37015));
    Odrv12 I__7619 (
            .O(N__37015),
            .I(\ALU.r0_12_prm_5_5_s0_c_RNOZ0 ));
    CascadeMux I__7618 (
            .O(N__37012),
            .I(N__37009));
    InMux I__7617 (
            .O(N__37009),
            .I(N__37006));
    LocalMux I__7616 (
            .O(N__37006),
            .I(N__37003));
    Span4Mux_h I__7615 (
            .O(N__37003),
            .I(N__37000));
    Span4Mux_v I__7614 (
            .O(N__37000),
            .I(N__36997));
    Odrv4 I__7613 (
            .O(N__36997),
            .I(\ALU.r4_RNIM8HG5Z0Z_5 ));
    InMux I__7612 (
            .O(N__36994),
            .I(N__36991));
    LocalMux I__7611 (
            .O(N__36991),
            .I(\ALU.r0_12_prm_3_5_s0_sf ));
    CascadeMux I__7610 (
            .O(N__36988),
            .I(N__36985));
    InMux I__7609 (
            .O(N__36985),
            .I(N__36982));
    LocalMux I__7608 (
            .O(N__36982),
            .I(N__36979));
    Odrv4 I__7607 (
            .O(N__36979),
            .I(\ALU.r0_12_prm_2_5_s0_c_RNOZ0 ));
    CascadeMux I__7606 (
            .O(N__36976),
            .I(N__36973));
    InMux I__7605 (
            .O(N__36973),
            .I(N__36970));
    LocalMux I__7604 (
            .O(N__36970),
            .I(N__36967));
    Odrv4 I__7603 (
            .O(N__36967),
            .I(\ALU.r0_12_prm_6_7_s0_c_RNOZ0 ));
    CascadeMux I__7602 (
            .O(N__36964),
            .I(N__36961));
    InMux I__7601 (
            .O(N__36961),
            .I(N__36958));
    LocalMux I__7600 (
            .O(N__36958),
            .I(\ALU.r4_RNIFR136Z0Z_7 ));
    InMux I__7599 (
            .O(N__36955),
            .I(N__36952));
    LocalMux I__7598 (
            .O(N__36952),
            .I(\ALU.r0_12_prm_3_7_s0_sf ));
    CascadeMux I__7597 (
            .O(N__36949),
            .I(N__36946));
    InMux I__7596 (
            .O(N__36946),
            .I(N__36943));
    LocalMux I__7595 (
            .O(N__36943),
            .I(\ALU.r0_12_prm_1_7_s0_c_RNOZ0 ));
    InMux I__7594 (
            .O(N__36940),
            .I(N__36937));
    LocalMux I__7593 (
            .O(N__36937),
            .I(N__36934));
    Span4Mux_v I__7592 (
            .O(N__36934),
            .I(N__36931));
    Span4Mux_h I__7591 (
            .O(N__36931),
            .I(N__36928));
    Odrv4 I__7590 (
            .O(N__36928),
            .I(\ALU.mult_7 ));
    InMux I__7589 (
            .O(N__36925),
            .I(\ALU.r0_12_s0_7 ));
    CascadeMux I__7588 (
            .O(N__36922),
            .I(N__36919));
    InMux I__7587 (
            .O(N__36919),
            .I(N__36914));
    InMux I__7586 (
            .O(N__36918),
            .I(N__36909));
    InMux I__7585 (
            .O(N__36917),
            .I(N__36909));
    LocalMux I__7584 (
            .O(N__36914),
            .I(N__36906));
    LocalMux I__7583 (
            .O(N__36909),
            .I(N__36903));
    Span4Mux_h I__7582 (
            .O(N__36906),
            .I(N__36900));
    Odrv4 I__7581 (
            .O(N__36903),
            .I(r1_7));
    Odrv4 I__7580 (
            .O(N__36900),
            .I(r1_7));
    CascadeMux I__7579 (
            .O(N__36895),
            .I(N__36892));
    InMux I__7578 (
            .O(N__36892),
            .I(N__36889));
    LocalMux I__7577 (
            .O(N__36889),
            .I(\ALU.lshift_3_ns_1_5 ));
    InMux I__7576 (
            .O(N__36886),
            .I(N__36883));
    LocalMux I__7575 (
            .O(N__36883),
            .I(N__36880));
    Odrv4 I__7574 (
            .O(N__36880),
            .I(\ALU.lshift_15_ns_1_9 ));
    CascadeMux I__7573 (
            .O(N__36877),
            .I(\ALU.r4_RNIF01FKZ0Z_2_cascade_ ));
    InMux I__7572 (
            .O(N__36874),
            .I(N__36871));
    LocalMux I__7571 (
            .O(N__36871),
            .I(N__36868));
    Span4Mux_h I__7570 (
            .O(N__36868),
            .I(N__36864));
    InMux I__7569 (
            .O(N__36867),
            .I(N__36861));
    Odrv4 I__7568 (
            .O(N__36864),
            .I(\ALU.r4_RNI2H9PKZ0Z_6 ));
    LocalMux I__7567 (
            .O(N__36861),
            .I(\ALU.r4_RNI2H9PKZ0Z_6 ));
    CascadeMux I__7566 (
            .O(N__36856),
            .I(\ALU.lshift_9_cascade_ ));
    CascadeMux I__7565 (
            .O(N__36853),
            .I(N__36850));
    InMux I__7564 (
            .O(N__36850),
            .I(N__36847));
    LocalMux I__7563 (
            .O(N__36847),
            .I(N__36844));
    Span4Mux_v I__7562 (
            .O(N__36844),
            .I(N__36841));
    Span4Mux_h I__7561 (
            .O(N__36841),
            .I(N__36838));
    Odrv4 I__7560 (
            .O(N__36838),
            .I(\ALU.r0_12_prm_8_9_s0_c_RNOZ0 ));
    InMux I__7559 (
            .O(N__36835),
            .I(N__36832));
    LocalMux I__7558 (
            .O(N__36832),
            .I(N__36829));
    Odrv4 I__7557 (
            .O(N__36829),
            .I(\ALU.rshift_15_ns_1_6 ));
    InMux I__7556 (
            .O(N__36826),
            .I(N__36823));
    LocalMux I__7555 (
            .O(N__36823),
            .I(\ALU.rshift_3_ns_1_5 ));
    CascadeMux I__7554 (
            .O(N__36820),
            .I(\ALU.r4_RNI9OH6AZ0Z_1_cascade_ ));
    InMux I__7553 (
            .O(N__36817),
            .I(N__36814));
    LocalMux I__7552 (
            .O(N__36814),
            .I(N__36811));
    Span12Mux_s9_v I__7551 (
            .O(N__36811),
            .I(N__36808));
    Odrv12 I__7550 (
            .O(N__36808),
            .I(\ALU.r5_RNIVQN52Z0Z_10 ));
    InMux I__7549 (
            .O(N__36805),
            .I(N__36802));
    LocalMux I__7548 (
            .O(N__36802),
            .I(N__36799));
    Span4Mux_h I__7547 (
            .O(N__36799),
            .I(N__36796));
    Span4Mux_h I__7546 (
            .O(N__36796),
            .I(N__36792));
    InMux I__7545 (
            .O(N__36795),
            .I(N__36789));
    Odrv4 I__7544 (
            .O(N__36792),
            .I(\ALU.r6_RNIP3372Z0Z_10 ));
    LocalMux I__7543 (
            .O(N__36789),
            .I(\ALU.r6_RNIP3372Z0Z_10 ));
    CascadeMux I__7542 (
            .O(N__36784),
            .I(N__36779));
    CascadeMux I__7541 (
            .O(N__36783),
            .I(N__36775));
    CascadeMux I__7540 (
            .O(N__36782),
            .I(N__36772));
    InMux I__7539 (
            .O(N__36779),
            .I(N__36760));
    CascadeMux I__7538 (
            .O(N__36778),
            .I(N__36756));
    InMux I__7537 (
            .O(N__36775),
            .I(N__36750));
    InMux I__7536 (
            .O(N__36772),
            .I(N__36747));
    CascadeMux I__7535 (
            .O(N__36771),
            .I(N__36744));
    CascadeMux I__7534 (
            .O(N__36770),
            .I(N__36741));
    CascadeMux I__7533 (
            .O(N__36769),
            .I(N__36738));
    CascadeMux I__7532 (
            .O(N__36768),
            .I(N__36735));
    CascadeMux I__7531 (
            .O(N__36767),
            .I(N__36731));
    CascadeMux I__7530 (
            .O(N__36766),
            .I(N__36728));
    CascadeMux I__7529 (
            .O(N__36765),
            .I(N__36725));
    InMux I__7528 (
            .O(N__36764),
            .I(N__36722));
    CascadeMux I__7527 (
            .O(N__36763),
            .I(N__36719));
    LocalMux I__7526 (
            .O(N__36760),
            .I(N__36716));
    InMux I__7525 (
            .O(N__36759),
            .I(N__36711));
    InMux I__7524 (
            .O(N__36756),
            .I(N__36711));
    CascadeMux I__7523 (
            .O(N__36755),
            .I(N__36708));
    CascadeMux I__7522 (
            .O(N__36754),
            .I(N__36705));
    CascadeMux I__7521 (
            .O(N__36753),
            .I(N__36702));
    LocalMux I__7520 (
            .O(N__36750),
            .I(N__36699));
    LocalMux I__7519 (
            .O(N__36747),
            .I(N__36694));
    InMux I__7518 (
            .O(N__36744),
            .I(N__36689));
    InMux I__7517 (
            .O(N__36741),
            .I(N__36689));
    InMux I__7516 (
            .O(N__36738),
            .I(N__36686));
    InMux I__7515 (
            .O(N__36735),
            .I(N__36682));
    InMux I__7514 (
            .O(N__36734),
            .I(N__36677));
    InMux I__7513 (
            .O(N__36731),
            .I(N__36674));
    InMux I__7512 (
            .O(N__36728),
            .I(N__36671));
    InMux I__7511 (
            .O(N__36725),
            .I(N__36668));
    LocalMux I__7510 (
            .O(N__36722),
            .I(N__36665));
    InMux I__7509 (
            .O(N__36719),
            .I(N__36661));
    Span4Mux_h I__7508 (
            .O(N__36716),
            .I(N__36656));
    LocalMux I__7507 (
            .O(N__36711),
            .I(N__36656));
    InMux I__7506 (
            .O(N__36708),
            .I(N__36651));
    InMux I__7505 (
            .O(N__36705),
            .I(N__36651));
    InMux I__7504 (
            .O(N__36702),
            .I(N__36648));
    Span4Mux_h I__7503 (
            .O(N__36699),
            .I(N__36645));
    InMux I__7502 (
            .O(N__36698),
            .I(N__36640));
    InMux I__7501 (
            .O(N__36697),
            .I(N__36640));
    Span4Mux_s1_v I__7500 (
            .O(N__36694),
            .I(N__36635));
    LocalMux I__7499 (
            .O(N__36689),
            .I(N__36635));
    LocalMux I__7498 (
            .O(N__36686),
            .I(N__36632));
    CascadeMux I__7497 (
            .O(N__36685),
            .I(N__36629));
    LocalMux I__7496 (
            .O(N__36682),
            .I(N__36626));
    CascadeMux I__7495 (
            .O(N__36681),
            .I(N__36622));
    CascadeMux I__7494 (
            .O(N__36680),
            .I(N__36618));
    LocalMux I__7493 (
            .O(N__36677),
            .I(N__36615));
    LocalMux I__7492 (
            .O(N__36674),
            .I(N__36610));
    LocalMux I__7491 (
            .O(N__36671),
            .I(N__36610));
    LocalMux I__7490 (
            .O(N__36668),
            .I(N__36607));
    Span4Mux_s2_h I__7489 (
            .O(N__36665),
            .I(N__36604));
    InMux I__7488 (
            .O(N__36664),
            .I(N__36601));
    LocalMux I__7487 (
            .O(N__36661),
            .I(N__36596));
    Span4Mux_v I__7486 (
            .O(N__36656),
            .I(N__36596));
    LocalMux I__7485 (
            .O(N__36651),
            .I(N__36593));
    LocalMux I__7484 (
            .O(N__36648),
            .I(N__36590));
    Span4Mux_s1_h I__7483 (
            .O(N__36645),
            .I(N__36585));
    LocalMux I__7482 (
            .O(N__36640),
            .I(N__36585));
    Span4Mux_h I__7481 (
            .O(N__36635),
            .I(N__36580));
    Span4Mux_v I__7480 (
            .O(N__36632),
            .I(N__36580));
    InMux I__7479 (
            .O(N__36629),
            .I(N__36577));
    Span4Mux_h I__7478 (
            .O(N__36626),
            .I(N__36574));
    InMux I__7477 (
            .O(N__36625),
            .I(N__36571));
    InMux I__7476 (
            .O(N__36622),
            .I(N__36564));
    InMux I__7475 (
            .O(N__36621),
            .I(N__36564));
    InMux I__7474 (
            .O(N__36618),
            .I(N__36564));
    Span4Mux_v I__7473 (
            .O(N__36615),
            .I(N__36560));
    Span4Mux_v I__7472 (
            .O(N__36610),
            .I(N__36557));
    Sp12to4 I__7471 (
            .O(N__36607),
            .I(N__36554));
    Span4Mux_h I__7470 (
            .O(N__36604),
            .I(N__36549));
    LocalMux I__7469 (
            .O(N__36601),
            .I(N__36549));
    Span4Mux_s2_h I__7468 (
            .O(N__36596),
            .I(N__36546));
    Span4Mux_v I__7467 (
            .O(N__36593),
            .I(N__36543));
    Span4Mux_s1_v I__7466 (
            .O(N__36590),
            .I(N__36534));
    Span4Mux_h I__7465 (
            .O(N__36585),
            .I(N__36534));
    Span4Mux_h I__7464 (
            .O(N__36580),
            .I(N__36534));
    LocalMux I__7463 (
            .O(N__36577),
            .I(N__36534));
    Span4Mux_v I__7462 (
            .O(N__36574),
            .I(N__36531));
    LocalMux I__7461 (
            .O(N__36571),
            .I(N__36526));
    LocalMux I__7460 (
            .O(N__36564),
            .I(N__36526));
    InMux I__7459 (
            .O(N__36563),
            .I(N__36523));
    Span4Mux_h I__7458 (
            .O(N__36560),
            .I(N__36520));
    Sp12to4 I__7457 (
            .O(N__36557),
            .I(N__36515));
    Span12Mux_s8_v I__7456 (
            .O(N__36554),
            .I(N__36515));
    Span4Mux_v I__7455 (
            .O(N__36549),
            .I(N__36508));
    Span4Mux_v I__7454 (
            .O(N__36546),
            .I(N__36508));
    Span4Mux_s2_h I__7453 (
            .O(N__36543),
            .I(N__36508));
    Span4Mux_v I__7452 (
            .O(N__36534),
            .I(N__36505));
    Sp12to4 I__7451 (
            .O(N__36531),
            .I(N__36500));
    Span12Mux_s8_v I__7450 (
            .O(N__36526),
            .I(N__36500));
    LocalMux I__7449 (
            .O(N__36523),
            .I(a_1_repZ0Z2));
    Odrv4 I__7448 (
            .O(N__36520),
            .I(a_1_repZ0Z2));
    Odrv12 I__7447 (
            .O(N__36515),
            .I(a_1_repZ0Z2));
    Odrv4 I__7446 (
            .O(N__36508),
            .I(a_1_repZ0Z2));
    Odrv4 I__7445 (
            .O(N__36505),
            .I(a_1_repZ0Z2));
    Odrv12 I__7444 (
            .O(N__36500),
            .I(a_1_repZ0Z2));
    InMux I__7443 (
            .O(N__36487),
            .I(N__36481));
    InMux I__7442 (
            .O(N__36486),
            .I(N__36481));
    LocalMux I__7441 (
            .O(N__36481),
            .I(N__36478));
    Span4Mux_s3_h I__7440 (
            .O(N__36478),
            .I(N__36475));
    Span4Mux_h I__7439 (
            .O(N__36475),
            .I(N__36472));
    Span4Mux_h I__7438 (
            .O(N__36472),
            .I(N__36469));
    Sp12to4 I__7437 (
            .O(N__36469),
            .I(N__36466));
    Odrv12 I__7436 (
            .O(N__36466),
            .I(\ALU.a10_b_4 ));
    InMux I__7435 (
            .O(N__36463),
            .I(N__36460));
    LocalMux I__7434 (
            .O(N__36460),
            .I(N__36457));
    Span4Mux_s2_v I__7433 (
            .O(N__36457),
            .I(N__36454));
    Span4Mux_h I__7432 (
            .O(N__36454),
            .I(N__36451));
    Odrv4 I__7431 (
            .O(N__36451),
            .I(\ALU.r0_12_prm_3_0_s1_c_RNOZ0 ));
    CascadeMux I__7430 (
            .O(N__36448),
            .I(N__36444));
    CascadeMux I__7429 (
            .O(N__36447),
            .I(N__36441));
    InMux I__7428 (
            .O(N__36444),
            .I(N__36434));
    InMux I__7427 (
            .O(N__36441),
            .I(N__36434));
    InMux I__7426 (
            .O(N__36440),
            .I(N__36429));
    InMux I__7425 (
            .O(N__36439),
            .I(N__36429));
    LocalMux I__7424 (
            .O(N__36434),
            .I(N__36426));
    LocalMux I__7423 (
            .O(N__36429),
            .I(N__36421));
    Span4Mux_h I__7422 (
            .O(N__36426),
            .I(N__36421));
    Span4Mux_v I__7421 (
            .O(N__36421),
            .I(N__36418));
    Odrv4 I__7420 (
            .O(N__36418),
            .I(\ALU.mult_0 ));
    InMux I__7419 (
            .O(N__36415),
            .I(N__36412));
    LocalMux I__7418 (
            .O(N__36412),
            .I(N__36409));
    Span4Mux_v I__7417 (
            .O(N__36409),
            .I(N__36406));
    Sp12to4 I__7416 (
            .O(N__36406),
            .I(N__36403));
    Odrv12 I__7415 (
            .O(N__36403),
            .I(\ALU.r0_12_prm_1_0_s1_c_RNOZ0 ));
    CascadeMux I__7414 (
            .O(N__36400),
            .I(N__36396));
    InMux I__7413 (
            .O(N__36399),
            .I(N__36393));
    InMux I__7412 (
            .O(N__36396),
            .I(N__36390));
    LocalMux I__7411 (
            .O(N__36393),
            .I(\ALU.un9_addsub_axb_0 ));
    LocalMux I__7410 (
            .O(N__36390),
            .I(\ALU.un9_addsub_axb_0 ));
    InMux I__7409 (
            .O(N__36385),
            .I(bfn_12_3_0_));
    InMux I__7408 (
            .O(N__36382),
            .I(N__36379));
    LocalMux I__7407 (
            .O(N__36379),
            .I(\ALU.r0_12_s1_0_THRU_CO ));
    InMux I__7406 (
            .O(N__36376),
            .I(N__36373));
    LocalMux I__7405 (
            .O(N__36373),
            .I(N__36370));
    Odrv4 I__7404 (
            .O(N__36370),
            .I(\ALU.rshift_15_ns_1_0 ));
    CascadeMux I__7403 (
            .O(N__36367),
            .I(N__36364));
    InMux I__7402 (
            .O(N__36364),
            .I(N__36361));
    LocalMux I__7401 (
            .O(N__36361),
            .I(\ALU.r0_12_prm_2_0_s0_c_RNOZ0 ));
    CascadeMux I__7400 (
            .O(N__36358),
            .I(N__36355));
    InMux I__7399 (
            .O(N__36355),
            .I(N__36352));
    LocalMux I__7398 (
            .O(N__36352),
            .I(\ALU.r0_12_prm_1_6_s1_c_RNOZ0 ));
    CascadeMux I__7397 (
            .O(N__36349),
            .I(\ALU.rshift_3_ns_1_4_cascade_ ));
    InMux I__7396 (
            .O(N__36346),
            .I(N__36343));
    LocalMux I__7395 (
            .O(N__36343),
            .I(N__36340));
    Span4Mux_s2_v I__7394 (
            .O(N__36340),
            .I(N__36337));
    Odrv4 I__7393 (
            .O(N__36337),
            .I(\ALU.r0_12_prm_7_0_s1_c_RNOZ0 ));
    InMux I__7392 (
            .O(N__36334),
            .I(N__36331));
    LocalMux I__7391 (
            .O(N__36331),
            .I(N__36328));
    Span4Mux_s1_v I__7390 (
            .O(N__36328),
            .I(N__36325));
    Span4Mux_h I__7389 (
            .O(N__36325),
            .I(N__36322));
    Span4Mux_h I__7388 (
            .O(N__36322),
            .I(N__36319));
    Odrv4 I__7387 (
            .O(N__36319),
            .I(\ALU.r0_12_prm_6_0_s1_c_RNOZ0 ));
    CascadeMux I__7386 (
            .O(N__36316),
            .I(N__36313));
    InMux I__7385 (
            .O(N__36313),
            .I(N__36309));
    InMux I__7384 (
            .O(N__36312),
            .I(N__36306));
    LocalMux I__7383 (
            .O(N__36309),
            .I(N__36303));
    LocalMux I__7382 (
            .O(N__36306),
            .I(N__36298));
    Span4Mux_s2_v I__7381 (
            .O(N__36303),
            .I(N__36298));
    Span4Mux_h I__7380 (
            .O(N__36298),
            .I(N__36295));
    Odrv4 I__7379 (
            .O(N__36295),
            .I(\ALU.un14_log_0_i_0 ));
    InMux I__7378 (
            .O(N__36292),
            .I(N__36289));
    LocalMux I__7377 (
            .O(N__36289),
            .I(\ALU.r0_12_prm_5_0_s1_c_RNOZ0 ));
    InMux I__7376 (
            .O(N__36286),
            .I(N__36283));
    LocalMux I__7375 (
            .O(N__36283),
            .I(\ALU.r0_12_prm_4_0_s1_c_RNOZ0 ));
    CascadeMux I__7374 (
            .O(N__36280),
            .I(N__36276));
    InMux I__7373 (
            .O(N__36279),
            .I(N__36273));
    InMux I__7372 (
            .O(N__36276),
            .I(N__36270));
    LocalMux I__7371 (
            .O(N__36273),
            .I(\ALU.N_883_i ));
    LocalMux I__7370 (
            .O(N__36270),
            .I(\ALU.N_883_i ));
    InMux I__7369 (
            .O(N__36265),
            .I(N__36262));
    LocalMux I__7368 (
            .O(N__36262),
            .I(\ALU.r0_12_prm_3_15_s0_sf ));
    InMux I__7367 (
            .O(N__36259),
            .I(N__36256));
    LocalMux I__7366 (
            .O(N__36256),
            .I(N__36253));
    Span4Mux_h I__7365 (
            .O(N__36253),
            .I(N__36249));
    InMux I__7364 (
            .O(N__36252),
            .I(N__36245));
    Span4Mux_h I__7363 (
            .O(N__36249),
            .I(N__36242));
    InMux I__7362 (
            .O(N__36248),
            .I(N__36239));
    LocalMux I__7361 (
            .O(N__36245),
            .I(N__36236));
    Span4Mux_v I__7360 (
            .O(N__36242),
            .I(N__36232));
    LocalMux I__7359 (
            .O(N__36239),
            .I(N__36229));
    Span4Mux_v I__7358 (
            .O(N__36236),
            .I(N__36226));
    InMux I__7357 (
            .O(N__36235),
            .I(N__36223));
    Odrv4 I__7356 (
            .O(N__36232),
            .I(\ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9 ));
    Odrv4 I__7355 (
            .O(N__36229),
            .I(\ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9 ));
    Odrv4 I__7354 (
            .O(N__36226),
            .I(\ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9 ));
    LocalMux I__7353 (
            .O(N__36223),
            .I(\ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9 ));
    CascadeMux I__7352 (
            .O(N__36214),
            .I(N__36211));
    InMux I__7351 (
            .O(N__36211),
            .I(N__36208));
    LocalMux I__7350 (
            .O(N__36208),
            .I(N__36205));
    Odrv4 I__7349 (
            .O(N__36205),
            .I(\ALU.r0_12_prm_2_15_s0_c_RNOZ0 ));
    InMux I__7348 (
            .O(N__36202),
            .I(N__36199));
    LocalMux I__7347 (
            .O(N__36199),
            .I(N__36196));
    Odrv12 I__7346 (
            .O(N__36196),
            .I(\ALU.r0_12_prm_1_15_s0_c_RNOZ0 ));
    InMux I__7345 (
            .O(N__36193),
            .I(\ALU.r0_12_s0_15 ));
    InMux I__7344 (
            .O(N__36190),
            .I(N__36187));
    LocalMux I__7343 (
            .O(N__36187),
            .I(N__36184));
    Span4Mux_v I__7342 (
            .O(N__36184),
            .I(N__36181));
    Sp12to4 I__7341 (
            .O(N__36181),
            .I(N__36178));
    Odrv12 I__7340 (
            .O(N__36178),
            .I(\ALU.r0_12_s0_15_THRU_CO ));
    CascadeMux I__7339 (
            .O(N__36175),
            .I(N__36172));
    InMux I__7338 (
            .O(N__36172),
            .I(N__36169));
    LocalMux I__7337 (
            .O(N__36169),
            .I(N__36166));
    Span4Mux_h I__7336 (
            .O(N__36166),
            .I(N__36163));
    Odrv4 I__7335 (
            .O(N__36163),
            .I(\ALU.r5_RNIB8HG5Z0Z_12 ));
    InMux I__7334 (
            .O(N__36160),
            .I(N__36156));
    CascadeMux I__7333 (
            .O(N__36159),
            .I(N__36153));
    LocalMux I__7332 (
            .O(N__36156),
            .I(N__36150));
    InMux I__7331 (
            .O(N__36153),
            .I(N__36147));
    Span4Mux_h I__7330 (
            .O(N__36150),
            .I(N__36142));
    LocalMux I__7329 (
            .O(N__36147),
            .I(N__36142));
    Span4Mux_h I__7328 (
            .O(N__36142),
            .I(N__36137));
    InMux I__7327 (
            .O(N__36141),
            .I(N__36134));
    InMux I__7326 (
            .O(N__36140),
            .I(N__36131));
    Sp12to4 I__7325 (
            .O(N__36137),
            .I(N__36124));
    LocalMux I__7324 (
            .O(N__36134),
            .I(N__36124));
    LocalMux I__7323 (
            .O(N__36131),
            .I(N__36124));
    Span12Mux_v I__7322 (
            .O(N__36124),
            .I(N__36121));
    Odrv12 I__7321 (
            .O(N__36121),
            .I(\ALU.lshift_13 ));
    InMux I__7320 (
            .O(N__36118),
            .I(N__36115));
    LocalMux I__7319 (
            .O(N__36115),
            .I(N__36112));
    Odrv4 I__7318 (
            .O(N__36112),
            .I(\ALU.r0_12_prm_8_13_s1_c_RNOZ0 ));
    InMux I__7317 (
            .O(N__36109),
            .I(N__36105));
    InMux I__7316 (
            .O(N__36108),
            .I(N__36102));
    LocalMux I__7315 (
            .O(N__36105),
            .I(N__36097));
    LocalMux I__7314 (
            .O(N__36102),
            .I(N__36094));
    InMux I__7313 (
            .O(N__36101),
            .I(N__36091));
    InMux I__7312 (
            .O(N__36100),
            .I(N__36088));
    Span4Mux_h I__7311 (
            .O(N__36097),
            .I(N__36081));
    Span4Mux_v I__7310 (
            .O(N__36094),
            .I(N__36081));
    LocalMux I__7309 (
            .O(N__36091),
            .I(N__36081));
    LocalMux I__7308 (
            .O(N__36088),
            .I(N__36078));
    Odrv4 I__7307 (
            .O(N__36081),
            .I(\ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8 ));
    Odrv12 I__7306 (
            .O(N__36078),
            .I(\ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8 ));
    CascadeMux I__7305 (
            .O(N__36073),
            .I(N__36070));
    InMux I__7304 (
            .O(N__36070),
            .I(N__36067));
    LocalMux I__7303 (
            .O(N__36067),
            .I(\ALU.r0_12_prm_1_10_s1_c_RNOZ0 ));
    CascadeMux I__7302 (
            .O(N__36064),
            .I(N__36061));
    InMux I__7301 (
            .O(N__36061),
            .I(N__36058));
    LocalMux I__7300 (
            .O(N__36058),
            .I(N__36055));
    Odrv12 I__7299 (
            .O(N__36055),
            .I(\ALU.r0_12_prm_1_12_s0_c_RNOZ0 ));
    CascadeMux I__7298 (
            .O(N__36052),
            .I(N__36049));
    InMux I__7297 (
            .O(N__36049),
            .I(N__36046));
    LocalMux I__7296 (
            .O(N__36046),
            .I(N__36043));
    Span4Mux_h I__7295 (
            .O(N__36043),
            .I(N__36040));
    Odrv4 I__7294 (
            .O(N__36040),
            .I(\ALU.r0_12_prm_2_14_s0_c_RNOZ0 ));
    InMux I__7293 (
            .O(N__36037),
            .I(N__36034));
    LocalMux I__7292 (
            .O(N__36034),
            .I(\ALU.rshift_15 ));
    InMux I__7291 (
            .O(N__36031),
            .I(N__36028));
    LocalMux I__7290 (
            .O(N__36028),
            .I(N__36024));
    InMux I__7289 (
            .O(N__36027),
            .I(N__36021));
    Span4Mux_v I__7288 (
            .O(N__36024),
            .I(N__36018));
    LocalMux I__7287 (
            .O(N__36021),
            .I(N__36015));
    Span4Mux_h I__7286 (
            .O(N__36018),
            .I(N__36008));
    Span4Mux_h I__7285 (
            .O(N__36015),
            .I(N__36008));
    InMux I__7284 (
            .O(N__36014),
            .I(N__36005));
    InMux I__7283 (
            .O(N__36013),
            .I(N__36002));
    Odrv4 I__7282 (
            .O(N__36008),
            .I(\ALU.lshift_15 ));
    LocalMux I__7281 (
            .O(N__36005),
            .I(\ALU.lshift_15 ));
    LocalMux I__7280 (
            .O(N__36002),
            .I(\ALU.lshift_15 ));
    CascadeMux I__7279 (
            .O(N__35995),
            .I(N__35992));
    InMux I__7278 (
            .O(N__35992),
            .I(N__35989));
    LocalMux I__7277 (
            .O(N__35989),
            .I(\ALU.r0_12_prm_8_15_s0_c_RNOZ0 ));
    InMux I__7276 (
            .O(N__35986),
            .I(N__35983));
    LocalMux I__7275 (
            .O(N__35983),
            .I(N__35979));
    CascadeMux I__7274 (
            .O(N__35982),
            .I(N__35976));
    Span4Mux_v I__7273 (
            .O(N__35979),
            .I(N__35973));
    InMux I__7272 (
            .O(N__35976),
            .I(N__35970));
    Sp12to4 I__7271 (
            .O(N__35973),
            .I(N__35965));
    LocalMux I__7270 (
            .O(N__35970),
            .I(N__35965));
    Odrv12 I__7269 (
            .O(N__35965),
            .I(\ALU.r2_RNI7AQC9_0Z0Z_15 ));
    InMux I__7268 (
            .O(N__35962),
            .I(N__35959));
    LocalMux I__7267 (
            .O(N__35959),
            .I(N__35956));
    Odrv4 I__7266 (
            .O(N__35956),
            .I(\ALU.r0_12_prm_6_15_s0_c_RNOZ0 ));
    CascadeMux I__7265 (
            .O(N__35953),
            .I(N__35950));
    InMux I__7264 (
            .O(N__35950),
            .I(N__35946));
    InMux I__7263 (
            .O(N__35949),
            .I(N__35943));
    LocalMux I__7262 (
            .O(N__35946),
            .I(N__35940));
    LocalMux I__7261 (
            .O(N__35943),
            .I(N__35937));
    Span4Mux_v I__7260 (
            .O(N__35940),
            .I(N__35934));
    Span4Mux_h I__7259 (
            .O(N__35937),
            .I(N__35931));
    Sp12to4 I__7258 (
            .O(N__35934),
            .I(N__35928));
    Sp12to4 I__7257 (
            .O(N__35931),
            .I(N__35923));
    Span12Mux_h I__7256 (
            .O(N__35928),
            .I(N__35923));
    Odrv12 I__7255 (
            .O(N__35923),
            .I(\ALU.un14_log_0_i_15 ));
    InMux I__7254 (
            .O(N__35920),
            .I(N__35917));
    LocalMux I__7253 (
            .O(N__35917),
            .I(N__35914));
    Odrv12 I__7252 (
            .O(N__35914),
            .I(\ALU.r0_12_prm_5_15_s0_c_RNOZ0 ));
    InMux I__7251 (
            .O(N__35911),
            .I(N__35907));
    CascadeMux I__7250 (
            .O(N__35910),
            .I(N__35904));
    LocalMux I__7249 (
            .O(N__35907),
            .I(N__35901));
    InMux I__7248 (
            .O(N__35904),
            .I(N__35898));
    Span4Mux_h I__7247 (
            .O(N__35901),
            .I(N__35895));
    LocalMux I__7246 (
            .O(N__35898),
            .I(N__35892));
    Odrv4 I__7245 (
            .O(N__35895),
            .I(\ALU.r2_RNI7AQC9_1Z0Z_15 ));
    Odrv4 I__7244 (
            .O(N__35892),
            .I(\ALU.r2_RNI7AQC9_1Z0Z_15 ));
    InMux I__7243 (
            .O(N__35887),
            .I(N__35884));
    LocalMux I__7242 (
            .O(N__35884),
            .I(\ALU.r5_RNI5P1F5Z0Z_15 ));
    InMux I__7241 (
            .O(N__35881),
            .I(N__35878));
    LocalMux I__7240 (
            .O(N__35878),
            .I(N__35875));
    Span4Mux_h I__7239 (
            .O(N__35875),
            .I(N__35871));
    CascadeMux I__7238 (
            .O(N__35874),
            .I(N__35868));
    Span4Mux_h I__7237 (
            .O(N__35871),
            .I(N__35865));
    InMux I__7236 (
            .O(N__35868),
            .I(N__35862));
    Odrv4 I__7235 (
            .O(N__35865),
            .I(\ALU.a_i_15 ));
    LocalMux I__7234 (
            .O(N__35862),
            .I(\ALU.a_i_15 ));
    CascadeMux I__7233 (
            .O(N__35857),
            .I(N__35854));
    InMux I__7232 (
            .O(N__35854),
            .I(N__35851));
    LocalMux I__7231 (
            .O(N__35851),
            .I(N__35848));
    Odrv12 I__7230 (
            .O(N__35848),
            .I(\ALU.r0_12_prm_2_10_s0_c_RNOZ0 ));
    CascadeMux I__7229 (
            .O(N__35845),
            .I(N__35841));
    InMux I__7228 (
            .O(N__35844),
            .I(N__35838));
    InMux I__7227 (
            .O(N__35841),
            .I(N__35835));
    LocalMux I__7226 (
            .O(N__35838),
            .I(N__35828));
    LocalMux I__7225 (
            .O(N__35835),
            .I(N__35828));
    InMux I__7224 (
            .O(N__35834),
            .I(N__35825));
    InMux I__7223 (
            .O(N__35833),
            .I(N__35822));
    Span12Mux_v I__7222 (
            .O(N__35828),
            .I(N__35819));
    LocalMux I__7221 (
            .O(N__35825),
            .I(N__35816));
    LocalMux I__7220 (
            .O(N__35822),
            .I(N__35813));
    Odrv12 I__7219 (
            .O(N__35819),
            .I(\ALU.un2_addsub_cry_10_c_RNIS4T7DZ0 ));
    Odrv4 I__7218 (
            .O(N__35816),
            .I(\ALU.un2_addsub_cry_10_c_RNIS4T7DZ0 ));
    Odrv4 I__7217 (
            .O(N__35813),
            .I(\ALU.un2_addsub_cry_10_c_RNIS4T7DZ0 ));
    CascadeMux I__7216 (
            .O(N__35806),
            .I(N__35803));
    InMux I__7215 (
            .O(N__35803),
            .I(N__35800));
    LocalMux I__7214 (
            .O(N__35800),
            .I(N__35797));
    Span4Mux_v I__7213 (
            .O(N__35797),
            .I(N__35794));
    Span4Mux_h I__7212 (
            .O(N__35794),
            .I(N__35791));
    Span4Mux_h I__7211 (
            .O(N__35791),
            .I(N__35788));
    Odrv4 I__7210 (
            .O(N__35788),
            .I(\ALU.r0_12_prm_2_11_s1_c_RNOZ0 ));
    InMux I__7209 (
            .O(N__35785),
            .I(N__35782));
    LocalMux I__7208 (
            .O(N__35782),
            .I(\ALU.r5_RNIAP7U9Z0Z_10 ));
    CascadeMux I__7207 (
            .O(N__35779),
            .I(\ALU.r5_RNIKU3HJZ0Z_10_cascade_ ));
    CascadeMux I__7206 (
            .O(N__35776),
            .I(\ALU.r4_RNIQK1V71Z0Z_5_cascade_ ));
    InMux I__7205 (
            .O(N__35773),
            .I(N__35769));
    InMux I__7204 (
            .O(N__35772),
            .I(N__35765));
    LocalMux I__7203 (
            .O(N__35769),
            .I(N__35762));
    InMux I__7202 (
            .O(N__35768),
            .I(N__35759));
    LocalMux I__7201 (
            .O(N__35765),
            .I(N__35752));
    Span4Mux_v I__7200 (
            .O(N__35762),
            .I(N__35752));
    LocalMux I__7199 (
            .O(N__35759),
            .I(N__35752));
    Span4Mux_v I__7198 (
            .O(N__35752),
            .I(N__35749));
    Span4Mux_h I__7197 (
            .O(N__35749),
            .I(N__35745));
    InMux I__7196 (
            .O(N__35748),
            .I(N__35742));
    Span4Mux_h I__7195 (
            .O(N__35745),
            .I(N__35739));
    LocalMux I__7194 (
            .O(N__35742),
            .I(N__35736));
    Odrv4 I__7193 (
            .O(N__35739),
            .I(\ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09 ));
    Odrv4 I__7192 (
            .O(N__35736),
            .I(\ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09 ));
    CascadeMux I__7191 (
            .O(N__35731),
            .I(N__35728));
    InMux I__7190 (
            .O(N__35728),
            .I(N__35725));
    LocalMux I__7189 (
            .O(N__35725),
            .I(N__35722));
    Span4Mux_v I__7188 (
            .O(N__35722),
            .I(N__35719));
    Span4Mux_h I__7187 (
            .O(N__35719),
            .I(N__35716));
    Odrv4 I__7186 (
            .O(N__35716),
            .I(\ALU.r0_12_prm_1_11_s0_c_RNOZ0 ));
    CascadeMux I__7185 (
            .O(N__35713),
            .I(N__35710));
    InMux I__7184 (
            .O(N__35710),
            .I(N__35707));
    LocalMux I__7183 (
            .O(N__35707),
            .I(N__35704));
    Span4Mux_h I__7182 (
            .O(N__35704),
            .I(N__35701));
    Span4Mux_v I__7181 (
            .O(N__35701),
            .I(N__35698));
    Odrv4 I__7180 (
            .O(N__35698),
            .I(\ALU.r0_12_prm_8_13_s0_c_RNOZ0 ));
    CascadeMux I__7179 (
            .O(N__35695),
            .I(N__35692));
    InMux I__7178 (
            .O(N__35692),
            .I(N__35689));
    LocalMux I__7177 (
            .O(N__35689),
            .I(N__35686));
    Span4Mux_h I__7176 (
            .O(N__35686),
            .I(N__35683));
    Span4Mux_v I__7175 (
            .O(N__35683),
            .I(N__35680));
    Odrv4 I__7174 (
            .O(N__35680),
            .I(\ALU.r0_12_prm_2_12_s0_c_RNOZ0 ));
    CascadeMux I__7173 (
            .O(N__35677),
            .I(N__35674));
    InMux I__7172 (
            .O(N__35674),
            .I(N__35671));
    LocalMux I__7171 (
            .O(N__35671),
            .I(N__35668));
    Odrv4 I__7170 (
            .O(N__35668),
            .I(\ALU.r0_12_prm_1_9_s0_c_RNOZ0 ));
    InMux I__7169 (
            .O(N__35665),
            .I(N__35662));
    LocalMux I__7168 (
            .O(N__35662),
            .I(N__35659));
    Odrv12 I__7167 (
            .O(N__35659),
            .I(\ALU.lshift_3_ns_1_13 ));
    InMux I__7166 (
            .O(N__35656),
            .I(N__35653));
    LocalMux I__7165 (
            .O(N__35653),
            .I(N__35650));
    Span4Mux_v I__7164 (
            .O(N__35650),
            .I(N__35647));
    Span4Mux_h I__7163 (
            .O(N__35647),
            .I(N__35644));
    Odrv4 I__7162 (
            .O(N__35644),
            .I(\ALU.rshift_12 ));
    InMux I__7161 (
            .O(N__35641),
            .I(N__35638));
    LocalMux I__7160 (
            .O(N__35638),
            .I(N__35633));
    InMux I__7159 (
            .O(N__35637),
            .I(N__35629));
    InMux I__7158 (
            .O(N__35636),
            .I(N__35626));
    Span4Mux_h I__7157 (
            .O(N__35633),
            .I(N__35623));
    InMux I__7156 (
            .O(N__35632),
            .I(N__35620));
    LocalMux I__7155 (
            .O(N__35629),
            .I(N__35615));
    LocalMux I__7154 (
            .O(N__35626),
            .I(N__35615));
    Odrv4 I__7153 (
            .O(N__35623),
            .I(\ALU.un2_addsub_cry_9_c_RNIS67KDZ0 ));
    LocalMux I__7152 (
            .O(N__35620),
            .I(\ALU.un2_addsub_cry_9_c_RNIS67KDZ0 ));
    Odrv12 I__7151 (
            .O(N__35615),
            .I(\ALU.un2_addsub_cry_9_c_RNIS67KDZ0 ));
    InMux I__7150 (
            .O(N__35608),
            .I(\ALU.un9_addsub_cry_9 ));
    InMux I__7149 (
            .O(N__35605),
            .I(N__35601));
    CascadeMux I__7148 (
            .O(N__35604),
            .I(N__35598));
    LocalMux I__7147 (
            .O(N__35601),
            .I(N__35595));
    InMux I__7146 (
            .O(N__35598),
            .I(N__35589));
    Span4Mux_v I__7145 (
            .O(N__35595),
            .I(N__35585));
    InMux I__7144 (
            .O(N__35594),
            .I(N__35582));
    CascadeMux I__7143 (
            .O(N__35593),
            .I(N__35574));
    CascadeMux I__7142 (
            .O(N__35592),
            .I(N__35570));
    LocalMux I__7141 (
            .O(N__35589),
            .I(N__35563));
    CascadeMux I__7140 (
            .O(N__35588),
            .I(N__35559));
    Span4Mux_h I__7139 (
            .O(N__35585),
            .I(N__35554));
    LocalMux I__7138 (
            .O(N__35582),
            .I(N__35554));
    InMux I__7137 (
            .O(N__35581),
            .I(N__35551));
    InMux I__7136 (
            .O(N__35580),
            .I(N__35548));
    InMux I__7135 (
            .O(N__35579),
            .I(N__35541));
    InMux I__7134 (
            .O(N__35578),
            .I(N__35541));
    InMux I__7133 (
            .O(N__35577),
            .I(N__35541));
    InMux I__7132 (
            .O(N__35574),
            .I(N__35534));
    InMux I__7131 (
            .O(N__35573),
            .I(N__35534));
    InMux I__7130 (
            .O(N__35570),
            .I(N__35531));
    InMux I__7129 (
            .O(N__35569),
            .I(N__35528));
    InMux I__7128 (
            .O(N__35568),
            .I(N__35521));
    InMux I__7127 (
            .O(N__35567),
            .I(N__35521));
    InMux I__7126 (
            .O(N__35566),
            .I(N__35521));
    Span4Mux_v I__7125 (
            .O(N__35563),
            .I(N__35518));
    InMux I__7124 (
            .O(N__35562),
            .I(N__35515));
    InMux I__7123 (
            .O(N__35559),
            .I(N__35512));
    Span4Mux_h I__7122 (
            .O(N__35554),
            .I(N__35507));
    LocalMux I__7121 (
            .O(N__35551),
            .I(N__35507));
    LocalMux I__7120 (
            .O(N__35548),
            .I(N__35502));
    LocalMux I__7119 (
            .O(N__35541),
            .I(N__35502));
    CascadeMux I__7118 (
            .O(N__35540),
            .I(N__35497));
    InMux I__7117 (
            .O(N__35539),
            .I(N__35493));
    LocalMux I__7116 (
            .O(N__35534),
            .I(N__35490));
    LocalMux I__7115 (
            .O(N__35531),
            .I(N__35483));
    LocalMux I__7114 (
            .O(N__35528),
            .I(N__35483));
    LocalMux I__7113 (
            .O(N__35521),
            .I(N__35483));
    Span4Mux_h I__7112 (
            .O(N__35518),
            .I(N__35478));
    LocalMux I__7111 (
            .O(N__35515),
            .I(N__35478));
    LocalMux I__7110 (
            .O(N__35512),
            .I(N__35473));
    Span4Mux_h I__7109 (
            .O(N__35507),
            .I(N__35473));
    Span12Mux_v I__7108 (
            .O(N__35502),
            .I(N__35470));
    InMux I__7107 (
            .O(N__35501),
            .I(N__35467));
    InMux I__7106 (
            .O(N__35500),
            .I(N__35460));
    InMux I__7105 (
            .O(N__35497),
            .I(N__35460));
    InMux I__7104 (
            .O(N__35496),
            .I(N__35460));
    LocalMux I__7103 (
            .O(N__35493),
            .I(N__35453));
    Span4Mux_v I__7102 (
            .O(N__35490),
            .I(N__35453));
    Span4Mux_v I__7101 (
            .O(N__35483),
            .I(N__35453));
    Span4Mux_h I__7100 (
            .O(N__35478),
            .I(N__35450));
    Span4Mux_v I__7099 (
            .O(N__35473),
            .I(N__35447));
    Odrv12 I__7098 (
            .O(N__35470),
            .I(\ALU.b_11 ));
    LocalMux I__7097 (
            .O(N__35467),
            .I(\ALU.b_11 ));
    LocalMux I__7096 (
            .O(N__35460),
            .I(\ALU.b_11 ));
    Odrv4 I__7095 (
            .O(N__35453),
            .I(\ALU.b_11 ));
    Odrv4 I__7094 (
            .O(N__35450),
            .I(\ALU.b_11 ));
    Odrv4 I__7093 (
            .O(N__35447),
            .I(\ALU.b_11 ));
    InMux I__7092 (
            .O(N__35434),
            .I(\ALU.un9_addsub_cry_10 ));
    InMux I__7091 (
            .O(N__35431),
            .I(\ALU.un9_addsub_cry_11 ));
    InMux I__7090 (
            .O(N__35428),
            .I(N__35421));
    CascadeMux I__7089 (
            .O(N__35427),
            .I(N__35418));
    CascadeMux I__7088 (
            .O(N__35426),
            .I(N__35415));
    CascadeMux I__7087 (
            .O(N__35425),
            .I(N__35412));
    CascadeMux I__7086 (
            .O(N__35424),
            .I(N__35407));
    LocalMux I__7085 (
            .O(N__35421),
            .I(N__35404));
    InMux I__7084 (
            .O(N__35418),
            .I(N__35393));
    InMux I__7083 (
            .O(N__35415),
            .I(N__35393));
    InMux I__7082 (
            .O(N__35412),
            .I(N__35393));
    InMux I__7081 (
            .O(N__35411),
            .I(N__35393));
    InMux I__7080 (
            .O(N__35410),
            .I(N__35393));
    InMux I__7079 (
            .O(N__35407),
            .I(N__35389));
    Span4Mux_v I__7078 (
            .O(N__35404),
            .I(N__35384));
    LocalMux I__7077 (
            .O(N__35393),
            .I(N__35381));
    InMux I__7076 (
            .O(N__35392),
            .I(N__35378));
    LocalMux I__7075 (
            .O(N__35389),
            .I(N__35375));
    InMux I__7074 (
            .O(N__35388),
            .I(N__35368));
    InMux I__7073 (
            .O(N__35387),
            .I(N__35368));
    Span4Mux_h I__7072 (
            .O(N__35384),
            .I(N__35361));
    Span4Mux_v I__7071 (
            .O(N__35381),
            .I(N__35361));
    LocalMux I__7070 (
            .O(N__35378),
            .I(N__35361));
    Span4Mux_v I__7069 (
            .O(N__35375),
            .I(N__35358));
    InMux I__7068 (
            .O(N__35374),
            .I(N__35355));
    InMux I__7067 (
            .O(N__35373),
            .I(N__35352));
    LocalMux I__7066 (
            .O(N__35368),
            .I(N__35349));
    Span4Mux_h I__7065 (
            .O(N__35361),
            .I(N__35344));
    Span4Mux_h I__7064 (
            .O(N__35358),
            .I(N__35341));
    LocalMux I__7063 (
            .O(N__35355),
            .I(N__35338));
    LocalMux I__7062 (
            .O(N__35352),
            .I(N__35335));
    Span4Mux_v I__7061 (
            .O(N__35349),
            .I(N__35332));
    InMux I__7060 (
            .O(N__35348),
            .I(N__35327));
    InMux I__7059 (
            .O(N__35347),
            .I(N__35327));
    Sp12to4 I__7058 (
            .O(N__35344),
            .I(N__35324));
    Span4Mux_h I__7057 (
            .O(N__35341),
            .I(N__35321));
    Span4Mux_v I__7056 (
            .O(N__35338),
            .I(N__35318));
    Span4Mux_s1_h I__7055 (
            .O(N__35335),
            .I(N__35313));
    Span4Mux_v I__7054 (
            .O(N__35332),
            .I(N__35313));
    LocalMux I__7053 (
            .O(N__35327),
            .I(\ALU.b_13 ));
    Odrv12 I__7052 (
            .O(N__35324),
            .I(\ALU.b_13 ));
    Odrv4 I__7051 (
            .O(N__35321),
            .I(\ALU.b_13 ));
    Odrv4 I__7050 (
            .O(N__35318),
            .I(\ALU.b_13 ));
    Odrv4 I__7049 (
            .O(N__35313),
            .I(\ALU.b_13 ));
    InMux I__7048 (
            .O(N__35302),
            .I(N__35297));
    InMux I__7047 (
            .O(N__35301),
            .I(N__35291));
    InMux I__7046 (
            .O(N__35300),
            .I(N__35291));
    LocalMux I__7045 (
            .O(N__35297),
            .I(N__35288));
    InMux I__7044 (
            .O(N__35296),
            .I(N__35285));
    LocalMux I__7043 (
            .O(N__35291),
            .I(N__35282));
    Span4Mux_v I__7042 (
            .O(N__35288),
            .I(N__35279));
    LocalMux I__7041 (
            .O(N__35285),
            .I(N__35274));
    Span4Mux_h I__7040 (
            .O(N__35282),
            .I(N__35274));
    Span4Mux_h I__7039 (
            .O(N__35279),
            .I(N__35269));
    Span4Mux_v I__7038 (
            .O(N__35274),
            .I(N__35269));
    Odrv4 I__7037 (
            .O(N__35269),
            .I(\ALU.un9_addsub_cry_12_c_RNISR30AZ0 ));
    InMux I__7036 (
            .O(N__35266),
            .I(\ALU.un9_addsub_cry_12 ));
    InMux I__7035 (
            .O(N__35263),
            .I(\ALU.un9_addsub_cry_13 ));
    InMux I__7034 (
            .O(N__35260),
            .I(\ALU.un9_addsub_cry_14 ));
    CascadeMux I__7033 (
            .O(N__35257),
            .I(N__35254));
    InMux I__7032 (
            .O(N__35254),
            .I(N__35251));
    LocalMux I__7031 (
            .O(N__35251),
            .I(N__35248));
    Span4Mux_v I__7030 (
            .O(N__35248),
            .I(N__35245));
    Span4Mux_h I__7029 (
            .O(N__35245),
            .I(N__35242));
    Odrv4 I__7028 (
            .O(N__35242),
            .I(\ALU.r0_12_prm_6_10_s0_c_RNOZ0 ));
    CascadeMux I__7027 (
            .O(N__35239),
            .I(N__35236));
    InMux I__7026 (
            .O(N__35236),
            .I(N__35233));
    LocalMux I__7025 (
            .O(N__35233),
            .I(N__35230));
    Span4Mux_h I__7024 (
            .O(N__35230),
            .I(N__35227));
    Span4Mux_v I__7023 (
            .O(N__35227),
            .I(N__35224));
    Odrv4 I__7022 (
            .O(N__35224),
            .I(\ALU.r4_RNI90J9EZ0Z_1 ));
    InMux I__7021 (
            .O(N__35221),
            .I(\ALU.un9_addsub_cry_0 ));
    InMux I__7020 (
            .O(N__35218),
            .I(N__35215));
    LocalMux I__7019 (
            .O(N__35215),
            .I(\ALU.r4_RNI468UDZ0Z_2 ));
    InMux I__7018 (
            .O(N__35212),
            .I(\ALU.un9_addsub_cry_1 ));
    CascadeMux I__7017 (
            .O(N__35209),
            .I(N__35206));
    InMux I__7016 (
            .O(N__35206),
            .I(N__35203));
    LocalMux I__7015 (
            .O(N__35203),
            .I(N__35200));
    Span4Mux_v I__7014 (
            .O(N__35200),
            .I(N__35197));
    Odrv4 I__7013 (
            .O(N__35197),
            .I(\ALU.r4_RNIUU8UDZ0Z_3 ));
    InMux I__7012 (
            .O(N__35194),
            .I(\ALU.un9_addsub_cry_2 ));
    InMux I__7011 (
            .O(N__35191),
            .I(N__35188));
    LocalMux I__7010 (
            .O(N__35188),
            .I(N__35185));
    Odrv4 I__7009 (
            .O(N__35185),
            .I(\ALU.r4_RNIQK1EDZ0Z_4 ));
    InMux I__7008 (
            .O(N__35182),
            .I(\ALU.un9_addsub_cry_3 ));
    InMux I__7007 (
            .O(N__35179),
            .I(\ALU.un9_addsub_cry_4 ));
    InMux I__7006 (
            .O(N__35176),
            .I(\ALU.un9_addsub_cry_5 ));
    InMux I__7005 (
            .O(N__35173),
            .I(\ALU.un9_addsub_cry_6 ));
    InMux I__7004 (
            .O(N__35170),
            .I(bfn_11_9_0_));
    InMux I__7003 (
            .O(N__35167),
            .I(\ALU.un9_addsub_cry_8 ));
    CascadeMux I__7002 (
            .O(N__35164),
            .I(\ALU.r5_RNI9S2TIZ0Z_11_cascade_ ));
    CascadeMux I__7001 (
            .O(N__35161),
            .I(\ALU.lshift_15_ns_1_13_cascade_ ));
    InMux I__7000 (
            .O(N__35158),
            .I(N__35155));
    LocalMux I__6999 (
            .O(N__35155),
            .I(N__35152));
    Odrv4 I__6998 (
            .O(N__35152),
            .I(\ALU.un9_addsub_axb_2 ));
    CascadeMux I__6997 (
            .O(N__35149),
            .I(N__35146));
    InMux I__6996 (
            .O(N__35146),
            .I(N__35142));
    InMux I__6995 (
            .O(N__35145),
            .I(N__35139));
    LocalMux I__6994 (
            .O(N__35142),
            .I(N__35136));
    LocalMux I__6993 (
            .O(N__35139),
            .I(N__35133));
    Span4Mux_h I__6992 (
            .O(N__35136),
            .I(N__35130));
    Span4Mux_h I__6991 (
            .O(N__35133),
            .I(N__35125));
    Span4Mux_v I__6990 (
            .O(N__35130),
            .I(N__35125));
    Span4Mux_v I__6989 (
            .O(N__35125),
            .I(N__35122));
    Span4Mux_h I__6988 (
            .O(N__35122),
            .I(N__35119));
    Odrv4 I__6987 (
            .O(N__35119),
            .I(\ALU.un14_log_0_i_11 ));
    InMux I__6986 (
            .O(N__35116),
            .I(N__35110));
    InMux I__6985 (
            .O(N__35115),
            .I(N__35110));
    LocalMux I__6984 (
            .O(N__35110),
            .I(N__35107));
    Span4Mux_h I__6983 (
            .O(N__35107),
            .I(N__35104));
    Odrv4 I__6982 (
            .O(N__35104),
            .I(\ALU.a6_b_0 ));
    CascadeMux I__6981 (
            .O(N__35101),
            .I(\ALU.lshift_3_ns_1_8_cascade_ ));
    CascadeMux I__6980 (
            .O(N__35098),
            .I(\ALU.r4_RNILIPV9Z0Z_6_cascade_ ));
    CascadeMux I__6979 (
            .O(N__35095),
            .I(\ALU.r4_RNI1G9PKZ0Z_6_cascade_ ));
    CascadeMux I__6978 (
            .O(N__35092),
            .I(N__35089));
    InMux I__6977 (
            .O(N__35089),
            .I(N__35086));
    LocalMux I__6976 (
            .O(N__35086),
            .I(N__35083));
    Span4Mux_h I__6975 (
            .O(N__35083),
            .I(N__35079));
    InMux I__6974 (
            .O(N__35082),
            .I(N__35076));
    Span4Mux_h I__6973 (
            .O(N__35079),
            .I(N__35073));
    LocalMux I__6972 (
            .O(N__35076),
            .I(N__35070));
    Span4Mux_v I__6971 (
            .O(N__35073),
            .I(N__35066));
    Span4Mux_v I__6970 (
            .O(N__35070),
            .I(N__35063));
    InMux I__6969 (
            .O(N__35069),
            .I(N__35060));
    Odrv4 I__6968 (
            .O(N__35066),
            .I(r0_1));
    Odrv4 I__6967 (
            .O(N__35063),
            .I(r0_1));
    LocalMux I__6966 (
            .O(N__35060),
            .I(r0_1));
    InMux I__6965 (
            .O(N__35053),
            .I(N__35050));
    LocalMux I__6964 (
            .O(N__35050),
            .I(N__35046));
    InMux I__6963 (
            .O(N__35049),
            .I(N__35043));
    Span4Mux_h I__6962 (
            .O(N__35046),
            .I(N__35037));
    LocalMux I__6961 (
            .O(N__35043),
            .I(N__35037));
    InMux I__6960 (
            .O(N__35042),
            .I(N__35034));
    Span4Mux_h I__6959 (
            .O(N__35037),
            .I(N__35031));
    LocalMux I__6958 (
            .O(N__35034),
            .I(r0_3));
    Odrv4 I__6957 (
            .O(N__35031),
            .I(r0_3));
    InMux I__6956 (
            .O(N__35026),
            .I(N__35022));
    InMux I__6955 (
            .O(N__35025),
            .I(N__35019));
    LocalMux I__6954 (
            .O(N__35022),
            .I(N__35013));
    LocalMux I__6953 (
            .O(N__35019),
            .I(N__35013));
    InMux I__6952 (
            .O(N__35018),
            .I(N__35010));
    Span4Mux_v I__6951 (
            .O(N__35013),
            .I(N__35004));
    LocalMux I__6950 (
            .O(N__35010),
            .I(N__35004));
    InMux I__6949 (
            .O(N__35009),
            .I(N__35001));
    Span4Mux_v I__6948 (
            .O(N__35004),
            .I(N__34997));
    LocalMux I__6947 (
            .O(N__35001),
            .I(N__34994));
    InMux I__6946 (
            .O(N__35000),
            .I(N__34991));
    Span4Mux_v I__6945 (
            .O(N__34997),
            .I(N__34988));
    Sp12to4 I__6944 (
            .O(N__34994),
            .I(N__34983));
    LocalMux I__6943 (
            .O(N__34991),
            .I(N__34980));
    Span4Mux_h I__6942 (
            .O(N__34988),
            .I(N__34977));
    InMux I__6941 (
            .O(N__34987),
            .I(N__34974));
    InMux I__6940 (
            .O(N__34986),
            .I(N__34971));
    Span12Mux_v I__6939 (
            .O(N__34983),
            .I(N__34967));
    Span12Mux_s10_h I__6938 (
            .O(N__34980),
            .I(N__34964));
    Span4Mux_h I__6937 (
            .O(N__34977),
            .I(N__34959));
    LocalMux I__6936 (
            .O(N__34974),
            .I(N__34959));
    LocalMux I__6935 (
            .O(N__34971),
            .I(N__34956));
    InMux I__6934 (
            .O(N__34970),
            .I(N__34953));
    Odrv12 I__6933 (
            .O(N__34967),
            .I(\ALU.r0_12_0 ));
    Odrv12 I__6932 (
            .O(N__34964),
            .I(\ALU.r0_12_0 ));
    Odrv4 I__6931 (
            .O(N__34959),
            .I(\ALU.r0_12_0 ));
    Odrv4 I__6930 (
            .O(N__34956),
            .I(\ALU.r0_12_0 ));
    LocalMux I__6929 (
            .O(N__34953),
            .I(\ALU.r0_12_0 ));
    InMux I__6928 (
            .O(N__34942),
            .I(N__34936));
    InMux I__6927 (
            .O(N__34941),
            .I(N__34936));
    LocalMux I__6926 (
            .O(N__34936),
            .I(N__34933));
    Span4Mux_h I__6925 (
            .O(N__34933),
            .I(N__34929));
    InMux I__6924 (
            .O(N__34932),
            .I(N__34926));
    Odrv4 I__6923 (
            .O(N__34929),
            .I(r0_0));
    LocalMux I__6922 (
            .O(N__34926),
            .I(r0_0));
    CascadeMux I__6921 (
            .O(N__34921),
            .I(N__34918));
    InMux I__6920 (
            .O(N__34918),
            .I(N__34915));
    LocalMux I__6919 (
            .O(N__34915),
            .I(\ALU.r0_12_prm_5_0_s0_c_RNOZ0 ));
    CascadeMux I__6918 (
            .O(N__34912),
            .I(N__34909));
    InMux I__6917 (
            .O(N__34909),
            .I(N__34906));
    LocalMux I__6916 (
            .O(N__34906),
            .I(N__34903));
    Span4Mux_s2_v I__6915 (
            .O(N__34903),
            .I(N__34900));
    Span4Mux_h I__6914 (
            .O(N__34900),
            .I(N__34897));
    Odrv4 I__6913 (
            .O(N__34897),
            .I(\ALU.r2_RNIKG5N5Z0Z_0 ));
    CascadeMux I__6912 (
            .O(N__34894),
            .I(N__34891));
    InMux I__6911 (
            .O(N__34891),
            .I(N__34888));
    LocalMux I__6910 (
            .O(N__34888),
            .I(N__34885));
    Odrv4 I__6909 (
            .O(N__34885),
            .I(\ALU.r0_12_prm_3_0_s0_c_RNOZ0 ));
    CascadeMux I__6908 (
            .O(N__34882),
            .I(N__34879));
    InMux I__6907 (
            .O(N__34879),
            .I(N__34876));
    LocalMux I__6906 (
            .O(N__34876),
            .I(N__34873));
    Span4Mux_h I__6905 (
            .O(N__34873),
            .I(N__34870));
    Odrv4 I__6904 (
            .O(N__34870),
            .I(\ALU.r0_12_prm_1_0_s0_c_RNOZ0 ));
    InMux I__6903 (
            .O(N__34867),
            .I(N__34864));
    LocalMux I__6902 (
            .O(N__34864),
            .I(N__34861));
    Odrv4 I__6901 (
            .O(N__34861),
            .I(\ALU.rshift_0 ));
    InMux I__6900 (
            .O(N__34858),
            .I(bfn_11_4_0_));
    InMux I__6899 (
            .O(N__34855),
            .I(N__34848));
    InMux I__6898 (
            .O(N__34854),
            .I(N__34848));
    CascadeMux I__6897 (
            .O(N__34853),
            .I(N__34845));
    LocalMux I__6896 (
            .O(N__34848),
            .I(N__34842));
    InMux I__6895 (
            .O(N__34845),
            .I(N__34839));
    Span4Mux_v I__6894 (
            .O(N__34842),
            .I(N__34836));
    LocalMux I__6893 (
            .O(N__34839),
            .I(N__34833));
    Span4Mux_h I__6892 (
            .O(N__34836),
            .I(N__34828));
    Span4Mux_v I__6891 (
            .O(N__34833),
            .I(N__34828));
    Odrv4 I__6890 (
            .O(N__34828),
            .I(r1_0));
    InMux I__6889 (
            .O(N__34825),
            .I(\ALU.r0_12_s1_6 ));
    CascadeMux I__6888 (
            .O(N__34822),
            .I(\ALU.lshift_6_cascade_ ));
    InMux I__6887 (
            .O(N__34819),
            .I(N__34816));
    LocalMux I__6886 (
            .O(N__34816),
            .I(\ALU.r0_12_prm_8_6_s1_c_RNOZ0 ));
    CascadeMux I__6885 (
            .O(N__34813),
            .I(N__34810));
    InMux I__6884 (
            .O(N__34810),
            .I(N__34807));
    LocalMux I__6883 (
            .O(N__34807),
            .I(N__34804));
    Odrv4 I__6882 (
            .O(N__34804),
            .I(\ALU.r0_12_prm_7_0_s0_c_RNOZ0 ));
    CascadeMux I__6881 (
            .O(N__34801),
            .I(N__34798));
    InMux I__6880 (
            .O(N__34798),
            .I(N__34795));
    LocalMux I__6879 (
            .O(N__34795),
            .I(N__34792));
    Odrv4 I__6878 (
            .O(N__34792),
            .I(\ALU.r0_12_prm_6_0_s0_c_RNOZ0 ));
    CascadeMux I__6877 (
            .O(N__34789),
            .I(N__34786));
    InMux I__6876 (
            .O(N__34786),
            .I(N__34783));
    LocalMux I__6875 (
            .O(N__34783),
            .I(\ALU.r0_12_prm_7_6_s1_c_RNOZ0 ));
    InMux I__6874 (
            .O(N__34780),
            .I(N__34777));
    LocalMux I__6873 (
            .O(N__34777),
            .I(\ALU.r0_12_prm_6_6_s1_c_RNOZ0 ));
    InMux I__6872 (
            .O(N__34774),
            .I(N__34771));
    LocalMux I__6871 (
            .O(N__34771),
            .I(N__34768));
    Odrv4 I__6870 (
            .O(N__34768),
            .I(\ALU.r0_12_prm_5_6_s1_c_RNOZ0 ));
    InMux I__6869 (
            .O(N__34765),
            .I(N__34762));
    LocalMux I__6868 (
            .O(N__34762),
            .I(N__34759));
    Span4Mux_h I__6867 (
            .O(N__34759),
            .I(N__34756));
    Odrv4 I__6866 (
            .O(N__34756),
            .I(\ALU.r0_12_prm_4_6_s1_c_RNOZ0 ));
    CascadeMux I__6865 (
            .O(N__34753),
            .I(N__34750));
    InMux I__6864 (
            .O(N__34750),
            .I(N__34747));
    LocalMux I__6863 (
            .O(N__34747),
            .I(\ALU.r0_12_prm_2_6_s1_c_RNOZ0 ));
    InMux I__6862 (
            .O(N__34744),
            .I(N__34741));
    LocalMux I__6861 (
            .O(N__34741),
            .I(\ALU.r0_12_prm_6_10_s1_c_RNOZ0 ));
    CascadeMux I__6860 (
            .O(N__34738),
            .I(N__34734));
    InMux I__6859 (
            .O(N__34737),
            .I(N__34731));
    InMux I__6858 (
            .O(N__34734),
            .I(N__34728));
    LocalMux I__6857 (
            .O(N__34731),
            .I(N__34725));
    LocalMux I__6856 (
            .O(N__34728),
            .I(N__34722));
    Span4Mux_v I__6855 (
            .O(N__34725),
            .I(N__34719));
    Span4Mux_v I__6854 (
            .O(N__34722),
            .I(N__34716));
    Odrv4 I__6853 (
            .O(N__34719),
            .I(\ALU.un14_log_0_i_10 ));
    Odrv4 I__6852 (
            .O(N__34716),
            .I(\ALU.un14_log_0_i_10 ));
    InMux I__6851 (
            .O(N__34711),
            .I(N__34708));
    LocalMux I__6850 (
            .O(N__34708),
            .I(\ALU.r0_12_prm_5_10_s1_c_RNOZ0 ));
    CascadeMux I__6849 (
            .O(N__34705),
            .I(N__34702));
    InMux I__6848 (
            .O(N__34702),
            .I(N__34699));
    LocalMux I__6847 (
            .O(N__34699),
            .I(N__34695));
    InMux I__6846 (
            .O(N__34698),
            .I(N__34692));
    Span4Mux_h I__6845 (
            .O(N__34695),
            .I(N__34689));
    LocalMux I__6844 (
            .O(N__34692),
            .I(N__34684));
    Span4Mux_v I__6843 (
            .O(N__34689),
            .I(N__34684));
    Odrv4 I__6842 (
            .O(N__34684),
            .I(\ALU.r5_RNIUF9K8_1Z0Z_10 ));
    InMux I__6841 (
            .O(N__34681),
            .I(N__34678));
    LocalMux I__6840 (
            .O(N__34678),
            .I(\ALU.r0_12_prm_4_10_s1_c_RNOZ0 ));
    CascadeMux I__6839 (
            .O(N__34675),
            .I(N__34672));
    InMux I__6838 (
            .O(N__34672),
            .I(N__34669));
    LocalMux I__6837 (
            .O(N__34669),
            .I(N__34666));
    Span4Mux_h I__6836 (
            .O(N__34666),
            .I(N__34662));
    InMux I__6835 (
            .O(N__34665),
            .I(N__34659));
    Span4Mux_v I__6834 (
            .O(N__34662),
            .I(N__34656));
    LocalMux I__6833 (
            .O(N__34659),
            .I(\ALU.a_i_10 ));
    Odrv4 I__6832 (
            .O(N__34656),
            .I(\ALU.a_i_10 ));
    CascadeMux I__6831 (
            .O(N__34651),
            .I(N__34648));
    InMux I__6830 (
            .O(N__34648),
            .I(N__34645));
    LocalMux I__6829 (
            .O(N__34645),
            .I(\ALU.r0_12_prm_2_10_s1_c_RNOZ0 ));
    InMux I__6828 (
            .O(N__34642),
            .I(\ALU.r0_12_s1_10 ));
    InMux I__6827 (
            .O(N__34639),
            .I(N__34636));
    LocalMux I__6826 (
            .O(N__34636),
            .I(N__34633));
    Span4Mux_h I__6825 (
            .O(N__34633),
            .I(N__34630));
    Span4Mux_v I__6824 (
            .O(N__34630),
            .I(N__34627));
    Odrv4 I__6823 (
            .O(N__34627),
            .I(\ALU.r0_12_s1_10_THRU_CO ));
    CascadeMux I__6822 (
            .O(N__34624),
            .I(N__34621));
    InMux I__6821 (
            .O(N__34621),
            .I(N__34618));
    LocalMux I__6820 (
            .O(N__34618),
            .I(N__34615));
    Odrv12 I__6819 (
            .O(N__34615),
            .I(\ALU.r0_12_prm_1_13_s0_c_RNOZ0 ));
    CascadeMux I__6818 (
            .O(N__34612),
            .I(N__34609));
    InMux I__6817 (
            .O(N__34609),
            .I(N__34606));
    LocalMux I__6816 (
            .O(N__34606),
            .I(N__34603));
    Span4Mux_h I__6815 (
            .O(N__34603),
            .I(N__34600));
    Odrv4 I__6814 (
            .O(N__34600),
            .I(\ALU.r5_RNI27VE5Z0Z_10 ));
    InMux I__6813 (
            .O(N__34597),
            .I(N__34593));
    CascadeMux I__6812 (
            .O(N__34596),
            .I(N__34590));
    LocalMux I__6811 (
            .O(N__34593),
            .I(N__34586));
    InMux I__6810 (
            .O(N__34590),
            .I(N__34583));
    InMux I__6809 (
            .O(N__34589),
            .I(N__34580));
    Span4Mux_v I__6808 (
            .O(N__34586),
            .I(N__34576));
    LocalMux I__6807 (
            .O(N__34583),
            .I(N__34571));
    LocalMux I__6806 (
            .O(N__34580),
            .I(N__34571));
    InMux I__6805 (
            .O(N__34579),
            .I(N__34568));
    Span4Mux_h I__6804 (
            .O(N__34576),
            .I(N__34563));
    Span4Mux_v I__6803 (
            .O(N__34571),
            .I(N__34563));
    LocalMux I__6802 (
            .O(N__34568),
            .I(N__34560));
    Odrv4 I__6801 (
            .O(N__34563),
            .I(\ALU.un2_addsub_cry_12_c_RNI74A7EZ0 ));
    Odrv12 I__6800 (
            .O(N__34560),
            .I(\ALU.un2_addsub_cry_12_c_RNI74A7EZ0 ));
    InMux I__6799 (
            .O(N__34555),
            .I(N__34552));
    LocalMux I__6798 (
            .O(N__34552),
            .I(\ALU.r0_12_prm_2_13_s1_c_RNOZ0 ));
    InMux I__6797 (
            .O(N__34549),
            .I(N__34546));
    LocalMux I__6796 (
            .O(N__34546),
            .I(N__34543));
    Span4Mux_h I__6795 (
            .O(N__34543),
            .I(N__34540));
    Span4Mux_h I__6794 (
            .O(N__34540),
            .I(N__34537));
    Odrv4 I__6793 (
            .O(N__34537),
            .I(\ALU.rshift_11 ));
    InMux I__6792 (
            .O(N__34534),
            .I(N__34531));
    LocalMux I__6791 (
            .O(N__34531),
            .I(N__34528));
    Span12Mux_v I__6790 (
            .O(N__34528),
            .I(N__34525));
    Odrv12 I__6789 (
            .O(N__34525),
            .I(\ALU.r0_12_prm_8_10_s1_c_RNOZ0Z_1 ));
    InMux I__6788 (
            .O(N__34522),
            .I(N__34519));
    LocalMux I__6787 (
            .O(N__34519),
            .I(N__34516));
    Odrv4 I__6786 (
            .O(N__34516),
            .I(\ALU.r0_12_prm_7_10_s1_c_RNOZ0 ));
    InMux I__6785 (
            .O(N__34513),
            .I(N__34509));
    CascadeMux I__6784 (
            .O(N__34512),
            .I(N__34506));
    LocalMux I__6783 (
            .O(N__34509),
            .I(N__34503));
    InMux I__6782 (
            .O(N__34506),
            .I(N__34500));
    Span4Mux_h I__6781 (
            .O(N__34503),
            .I(N__34497));
    LocalMux I__6780 (
            .O(N__34500),
            .I(N__34494));
    Odrv4 I__6779 (
            .O(N__34497),
            .I(\ALU.r5_RNIUF9K8_0Z0Z_10 ));
    Odrv4 I__6778 (
            .O(N__34494),
            .I(\ALU.r5_RNIUF9K8_0Z0Z_10 ));
    InMux I__6777 (
            .O(N__34489),
            .I(N__34486));
    LocalMux I__6776 (
            .O(N__34486),
            .I(N__34483));
    Odrv12 I__6775 (
            .O(N__34483),
            .I(\ALU.N_884_i ));
    CascadeMux I__6774 (
            .O(N__34480),
            .I(N__34477));
    InMux I__6773 (
            .O(N__34477),
            .I(N__34474));
    LocalMux I__6772 (
            .O(N__34474),
            .I(N__34471));
    Span4Mux_v I__6771 (
            .O(N__34471),
            .I(N__34468));
    Odrv4 I__6770 (
            .O(N__34468),
            .I(\ALU.r0_12_prm_8_12_s0_c_RNOZ0 ));
    CascadeMux I__6769 (
            .O(N__34465),
            .I(\ALU.lshift_3_ns_1_3_cascade_ ));
    InMux I__6768 (
            .O(N__34462),
            .I(N__34458));
    InMux I__6767 (
            .O(N__34461),
            .I(N__34455));
    LocalMux I__6766 (
            .O(N__34458),
            .I(N__34450));
    LocalMux I__6765 (
            .O(N__34455),
            .I(N__34450));
    Odrv12 I__6764 (
            .O(N__34450),
            .I(\ALU.r4_RNI1RK3KZ0Z_9 ));
    CascadeMux I__6763 (
            .O(N__34447),
            .I(\ALU.r4_RNIOK1781Z0Z_9_cascade_ ));
    InMux I__6762 (
            .O(N__34444),
            .I(N__34440));
    InMux I__6761 (
            .O(N__34443),
            .I(N__34437));
    LocalMux I__6760 (
            .O(N__34440),
            .I(N__34434));
    LocalMux I__6759 (
            .O(N__34437),
            .I(N__34431));
    Span4Mux_h I__6758 (
            .O(N__34434),
            .I(N__34428));
    Span4Mux_h I__6757 (
            .O(N__34431),
            .I(N__34425));
    Span4Mux_h I__6756 (
            .O(N__34428),
            .I(N__34418));
    Span4Mux_h I__6755 (
            .O(N__34425),
            .I(N__34418));
    InMux I__6754 (
            .O(N__34424),
            .I(N__34415));
    InMux I__6753 (
            .O(N__34423),
            .I(N__34412));
    Odrv4 I__6752 (
            .O(N__34418),
            .I(\ALU.lshift_11 ));
    LocalMux I__6751 (
            .O(N__34415),
            .I(\ALU.lshift_11 ));
    LocalMux I__6750 (
            .O(N__34412),
            .I(\ALU.lshift_11 ));
    InMux I__6749 (
            .O(N__34405),
            .I(N__34402));
    LocalMux I__6748 (
            .O(N__34402),
            .I(N__34398));
    InMux I__6747 (
            .O(N__34401),
            .I(N__34395));
    Span4Mux_h I__6746 (
            .O(N__34398),
            .I(N__34392));
    LocalMux I__6745 (
            .O(N__34395),
            .I(N__34388));
    Span4Mux_v I__6744 (
            .O(N__34392),
            .I(N__34385));
    InMux I__6743 (
            .O(N__34391),
            .I(N__34382));
    Span12Mux_s10_v I__6742 (
            .O(N__34388),
            .I(N__34379));
    Span4Mux_h I__6741 (
            .O(N__34385),
            .I(N__34374));
    LocalMux I__6740 (
            .O(N__34382),
            .I(N__34374));
    Odrv12 I__6739 (
            .O(N__34379),
            .I(r4_9));
    Odrv4 I__6738 (
            .O(N__34374),
            .I(r4_9));
    InMux I__6737 (
            .O(N__34369),
            .I(N__34365));
    InMux I__6736 (
            .O(N__34368),
            .I(N__34362));
    LocalMux I__6735 (
            .O(N__34365),
            .I(N__34358));
    LocalMux I__6734 (
            .O(N__34362),
            .I(N__34355));
    InMux I__6733 (
            .O(N__34361),
            .I(N__34352));
    Span4Mux_h I__6732 (
            .O(N__34358),
            .I(N__34349));
    Span4Mux_h I__6731 (
            .O(N__34355),
            .I(N__34346));
    LocalMux I__6730 (
            .O(N__34352),
            .I(N__34343));
    Span4Mux_h I__6729 (
            .O(N__34349),
            .I(N__34338));
    Span4Mux_v I__6728 (
            .O(N__34346),
            .I(N__34338));
    Odrv4 I__6727 (
            .O(N__34343),
            .I(r4_1));
    Odrv4 I__6726 (
            .O(N__34338),
            .I(r4_1));
    InMux I__6725 (
            .O(N__34333),
            .I(N__34330));
    LocalMux I__6724 (
            .O(N__34330),
            .I(N__34326));
    InMux I__6723 (
            .O(N__34329),
            .I(N__34322));
    Span4Mux_v I__6722 (
            .O(N__34326),
            .I(N__34319));
    InMux I__6721 (
            .O(N__34325),
            .I(N__34316));
    LocalMux I__6720 (
            .O(N__34322),
            .I(N__34313));
    Span4Mux_h I__6719 (
            .O(N__34319),
            .I(N__34310));
    LocalMux I__6718 (
            .O(N__34316),
            .I(N__34305));
    Span4Mux_h I__6717 (
            .O(N__34313),
            .I(N__34305));
    Odrv4 I__6716 (
            .O(N__34310),
            .I(r4_2));
    Odrv4 I__6715 (
            .O(N__34305),
            .I(r4_2));
    InMux I__6714 (
            .O(N__34300),
            .I(N__34297));
    LocalMux I__6713 (
            .O(N__34297),
            .I(N__34294));
    Span4Mux_v I__6712 (
            .O(N__34294),
            .I(N__34291));
    Span4Mux_h I__6711 (
            .O(N__34291),
            .I(N__34286));
    InMux I__6710 (
            .O(N__34290),
            .I(N__34283));
    InMux I__6709 (
            .O(N__34289),
            .I(N__34280));
    Span4Mux_h I__6708 (
            .O(N__34286),
            .I(N__34277));
    LocalMux I__6707 (
            .O(N__34283),
            .I(N__34274));
    LocalMux I__6706 (
            .O(N__34280),
            .I(N__34271));
    Span4Mux_h I__6705 (
            .O(N__34277),
            .I(N__34268));
    Span4Mux_h I__6704 (
            .O(N__34274),
            .I(N__34263));
    Span4Mux_v I__6703 (
            .O(N__34271),
            .I(N__34263));
    Odrv4 I__6702 (
            .O(N__34268),
            .I(r4_4));
    Odrv4 I__6701 (
            .O(N__34263),
            .I(r4_4));
    InMux I__6700 (
            .O(N__34258),
            .I(N__34255));
    LocalMux I__6699 (
            .O(N__34255),
            .I(N__34252));
    Span4Mux_h I__6698 (
            .O(N__34252),
            .I(N__34249));
    Span4Mux_v I__6697 (
            .O(N__34249),
            .I(N__34246));
    Span4Mux_h I__6696 (
            .O(N__34246),
            .I(N__34243));
    Span4Mux_h I__6695 (
            .O(N__34243),
            .I(N__34240));
    Odrv4 I__6694 (
            .O(N__34240),
            .I(\ALU.r5_RNIVF7TIZ0Z_13 ));
    CascadeMux I__6693 (
            .O(N__34237),
            .I(\ALU.lshift_15_ns_1_15_cascade_ ));
    InMux I__6692 (
            .O(N__34234),
            .I(N__34231));
    LocalMux I__6691 (
            .O(N__34231),
            .I(N__34228));
    Span4Mux_h I__6690 (
            .O(N__34228),
            .I(N__34225));
    Span4Mux_h I__6689 (
            .O(N__34225),
            .I(N__34222));
    Span4Mux_h I__6688 (
            .O(N__34222),
            .I(N__34219));
    Odrv4 I__6687 (
            .O(N__34219),
            .I(\ALU.r0_12_prm_8_11_s1_c_RNOZ0Z_1 ));
    InMux I__6686 (
            .O(N__34216),
            .I(N__34213));
    LocalMux I__6685 (
            .O(N__34213),
            .I(N__34210));
    Span4Mux_h I__6684 (
            .O(N__34210),
            .I(N__34207));
    Span4Mux_h I__6683 (
            .O(N__34207),
            .I(N__34204));
    Odrv4 I__6682 (
            .O(N__34204),
            .I(\ALU.r0_12_prm_2_11_s0_c_RNOZ0 ));
    CascadeMux I__6681 (
            .O(N__34201),
            .I(N__34198));
    InMux I__6680 (
            .O(N__34198),
            .I(N__34195));
    LocalMux I__6679 (
            .O(N__34195),
            .I(N__34192));
    Odrv4 I__6678 (
            .O(N__34192),
            .I(\ALU.r0_12_prm_1_10_s0_c_RNOZ0 ));
    CascadeMux I__6677 (
            .O(N__34189),
            .I(N__34186));
    InMux I__6676 (
            .O(N__34186),
            .I(N__34183));
    LocalMux I__6675 (
            .O(N__34183),
            .I(N__34180));
    Span4Mux_h I__6674 (
            .O(N__34180),
            .I(N__34177));
    Span4Mux_h I__6673 (
            .O(N__34177),
            .I(N__34174));
    Odrv4 I__6672 (
            .O(N__34174),
            .I(\ALU.r5_RNIUF9K8_2Z0Z_10 ));
    InMux I__6671 (
            .O(N__34171),
            .I(\ALU.un2_addsub_cry_9 ));
    CascadeMux I__6670 (
            .O(N__34168),
            .I(N__34165));
    InMux I__6669 (
            .O(N__34165),
            .I(N__34162));
    LocalMux I__6668 (
            .O(N__34162),
            .I(N__34159));
    Span4Mux_v I__6667 (
            .O(N__34159),
            .I(N__34156));
    Span4Mux_h I__6666 (
            .O(N__34156),
            .I(N__34153));
    Span4Mux_h I__6665 (
            .O(N__34153),
            .I(N__34150));
    Odrv4 I__6664 (
            .O(N__34150),
            .I(\ALU.r5_RNIE0AK8_2Z0Z_11 ));
    InMux I__6663 (
            .O(N__34147),
            .I(\ALU.un2_addsub_cry_10 ));
    CascadeMux I__6662 (
            .O(N__34144),
            .I(N__34141));
    InMux I__6661 (
            .O(N__34141),
            .I(N__34138));
    LocalMux I__6660 (
            .O(N__34138),
            .I(N__34135));
    Odrv12 I__6659 (
            .O(N__34135),
            .I(\ALU.r5_RNISP2L9_2Z0Z_12 ));
    InMux I__6658 (
            .O(N__34132),
            .I(\ALU.un2_addsub_cry_11 ));
    CascadeMux I__6657 (
            .O(N__34129),
            .I(N__34126));
    InMux I__6656 (
            .O(N__34126),
            .I(N__34123));
    LocalMux I__6655 (
            .O(N__34123),
            .I(N__34120));
    Span4Mux_h I__6654 (
            .O(N__34120),
            .I(N__34117));
    Span4Mux_h I__6653 (
            .O(N__34117),
            .I(N__34114));
    Odrv4 I__6652 (
            .O(N__34114),
            .I(\ALU.r5_RNID2JJ9_2Z0Z_13 ));
    InMux I__6651 (
            .O(N__34111),
            .I(\ALU.un2_addsub_cry_12 ));
    CascadeMux I__6650 (
            .O(N__34108),
            .I(N__34105));
    InMux I__6649 (
            .O(N__34105),
            .I(N__34102));
    LocalMux I__6648 (
            .O(N__34102),
            .I(N__34099));
    Odrv12 I__6647 (
            .O(N__34099),
            .I(\ALU.r2_RNINPPC9_2Z0Z_14 ));
    InMux I__6646 (
            .O(N__34096),
            .I(\ALU.un2_addsub_cry_13 ));
    InMux I__6645 (
            .O(N__34093),
            .I(\ALU.un2_addsub_cry_14 ));
    InMux I__6644 (
            .O(N__34090),
            .I(N__34084));
    InMux I__6643 (
            .O(N__34089),
            .I(N__34084));
    LocalMux I__6642 (
            .O(N__34084),
            .I(N__34080));
    InMux I__6641 (
            .O(N__34083),
            .I(N__34077));
    Span4Mux_h I__6640 (
            .O(N__34080),
            .I(N__34072));
    LocalMux I__6639 (
            .O(N__34077),
            .I(N__34072));
    Odrv4 I__6638 (
            .O(N__34072),
            .I(r4_7));
    InMux I__6637 (
            .O(N__34069),
            .I(N__34066));
    LocalMux I__6636 (
            .O(N__34066),
            .I(N__34062));
    InMux I__6635 (
            .O(N__34065),
            .I(N__34059));
    Span4Mux_s2_v I__6634 (
            .O(N__34062),
            .I(N__34056));
    LocalMux I__6633 (
            .O(N__34059),
            .I(N__34052));
    Span4Mux_h I__6632 (
            .O(N__34056),
            .I(N__34049));
    InMux I__6631 (
            .O(N__34055),
            .I(N__34046));
    Span4Mux_h I__6630 (
            .O(N__34052),
            .I(N__34043));
    Span4Mux_v I__6629 (
            .O(N__34049),
            .I(N__34038));
    LocalMux I__6628 (
            .O(N__34046),
            .I(N__34038));
    Odrv4 I__6627 (
            .O(N__34043),
            .I(r4_8));
    Odrv4 I__6626 (
            .O(N__34038),
            .I(r4_8));
    InMux I__6625 (
            .O(N__34033),
            .I(N__34028));
    InMux I__6624 (
            .O(N__34032),
            .I(N__34023));
    InMux I__6623 (
            .O(N__34031),
            .I(N__34019));
    LocalMux I__6622 (
            .O(N__34028),
            .I(N__34016));
    InMux I__6621 (
            .O(N__34027),
            .I(N__34011));
    InMux I__6620 (
            .O(N__34026),
            .I(N__34008));
    LocalMux I__6619 (
            .O(N__34023),
            .I(N__34005));
    InMux I__6618 (
            .O(N__34022),
            .I(N__34002));
    LocalMux I__6617 (
            .O(N__34019),
            .I(N__33997));
    Span4Mux_v I__6616 (
            .O(N__34016),
            .I(N__33997));
    InMux I__6615 (
            .O(N__34015),
            .I(N__33994));
    InMux I__6614 (
            .O(N__34014),
            .I(N__33991));
    LocalMux I__6613 (
            .O(N__34011),
            .I(N__33988));
    LocalMux I__6612 (
            .O(N__34008),
            .I(N__33983));
    Span4Mux_v I__6611 (
            .O(N__34005),
            .I(N__33983));
    LocalMux I__6610 (
            .O(N__34002),
            .I(N__33978));
    Span4Mux_h I__6609 (
            .O(N__33997),
            .I(N__33978));
    LocalMux I__6608 (
            .O(N__33994),
            .I(N__33969));
    LocalMux I__6607 (
            .O(N__33991),
            .I(N__33969));
    Span4Mux_v I__6606 (
            .O(N__33988),
            .I(N__33969));
    Span4Mux_h I__6605 (
            .O(N__33983),
            .I(N__33969));
    Odrv4 I__6604 (
            .O(N__33978),
            .I(\ALU.r0_12_9 ));
    Odrv4 I__6603 (
            .O(N__33969),
            .I(\ALU.r0_12_9 ));
    InMux I__6602 (
            .O(N__33964),
            .I(\ALU.un2_addsub_cry_0 ));
    InMux I__6601 (
            .O(N__33961),
            .I(N__33958));
    LocalMux I__6600 (
            .O(N__33958),
            .I(N__33955));
    Span4Mux_v I__6599 (
            .O(N__33955),
            .I(N__33952));
    Odrv4 I__6598 (
            .O(N__33952),
            .I(\ALU.r4_RNIUM9JCZ0Z_2 ));
    CascadeMux I__6597 (
            .O(N__33949),
            .I(N__33946));
    InMux I__6596 (
            .O(N__33946),
            .I(N__33943));
    LocalMux I__6595 (
            .O(N__33943),
            .I(N__33940));
    Span4Mux_v I__6594 (
            .O(N__33940),
            .I(N__33937));
    Span4Mux_v I__6593 (
            .O(N__33937),
            .I(N__33933));
    InMux I__6592 (
            .O(N__33936),
            .I(N__33930));
    Odrv4 I__6591 (
            .O(N__33933),
            .I(\ALU.b_i_2 ));
    LocalMux I__6590 (
            .O(N__33930),
            .I(\ALU.b_i_2 ));
    InMux I__6589 (
            .O(N__33925),
            .I(\ALU.un2_addsub_cry_1 ));
    InMux I__6588 (
            .O(N__33922),
            .I(N__33919));
    LocalMux I__6587 (
            .O(N__33919),
            .I(N__33916));
    Sp12to4 I__6586 (
            .O(N__33916),
            .I(N__33913));
    Odrv12 I__6585 (
            .O(N__33913),
            .I(\ALU.r4_RNINFAJCZ0Z_3 ));
    CascadeMux I__6584 (
            .O(N__33910),
            .I(N__33907));
    InMux I__6583 (
            .O(N__33907),
            .I(N__33904));
    LocalMux I__6582 (
            .O(N__33904),
            .I(N__33901));
    Span12Mux_h I__6581 (
            .O(N__33901),
            .I(N__33898));
    Odrv12 I__6580 (
            .O(N__33898),
            .I(\ALU.b_i_3 ));
    InMux I__6579 (
            .O(N__33895),
            .I(\ALU.un2_addsub_cry_2 ));
    InMux I__6578 (
            .O(N__33892),
            .I(N__33889));
    LocalMux I__6577 (
            .O(N__33889),
            .I(N__33886));
    Odrv12 I__6576 (
            .O(N__33886),
            .I(\ALU.r4_RNI20C8CZ0Z_4 ));
    CascadeMux I__6575 (
            .O(N__33883),
            .I(N__33879));
    InMux I__6574 (
            .O(N__33882),
            .I(N__33876));
    InMux I__6573 (
            .O(N__33879),
            .I(N__33873));
    LocalMux I__6572 (
            .O(N__33876),
            .I(N__33870));
    LocalMux I__6571 (
            .O(N__33873),
            .I(N__33867));
    Span4Mux_h I__6570 (
            .O(N__33870),
            .I(N__33864));
    Span4Mux_h I__6569 (
            .O(N__33867),
            .I(N__33859));
    Span4Mux_v I__6568 (
            .O(N__33864),
            .I(N__33859));
    Odrv4 I__6567 (
            .O(N__33859),
            .I(\ALU.b_i_4 ));
    InMux I__6566 (
            .O(N__33856),
            .I(\ALU.un2_addsub_cry_3 ));
    CascadeMux I__6565 (
            .O(N__33853),
            .I(N__33850));
    InMux I__6564 (
            .O(N__33850),
            .I(N__33847));
    LocalMux I__6563 (
            .O(N__33847),
            .I(N__33844));
    Span4Mux_v I__6562 (
            .O(N__33844),
            .I(N__33841));
    Sp12to4 I__6561 (
            .O(N__33841),
            .I(N__33838));
    Odrv12 I__6560 (
            .O(N__33838),
            .I(\ALU.r4_RNI8B628_1Z0Z_5 ));
    InMux I__6559 (
            .O(N__33835),
            .I(\ALU.un2_addsub_cry_4 ));
    CascadeMux I__6558 (
            .O(N__33832),
            .I(N__33829));
    InMux I__6557 (
            .O(N__33829),
            .I(N__33826));
    LocalMux I__6556 (
            .O(N__33826),
            .I(N__33823));
    Span4Mux_v I__6555 (
            .O(N__33823),
            .I(N__33820));
    Span4Mux_h I__6554 (
            .O(N__33820),
            .I(N__33817));
    Span4Mux_v I__6553 (
            .O(N__33817),
            .I(N__33814));
    Span4Mux_s3_v I__6552 (
            .O(N__33814),
            .I(N__33811));
    Odrv4 I__6551 (
            .O(N__33811),
            .I(\ALU.r4_RNI2BKQ8_1Z0Z_6 ));
    InMux I__6550 (
            .O(N__33808),
            .I(\ALU.un2_addsub_cry_5 ));
    InMux I__6549 (
            .O(N__33805),
            .I(\ALU.un2_addsub_cry_6 ));
    CascadeMux I__6548 (
            .O(N__33802),
            .I(N__33799));
    InMux I__6547 (
            .O(N__33799),
            .I(N__33796));
    LocalMux I__6546 (
            .O(N__33796),
            .I(N__33793));
    Odrv12 I__6545 (
            .O(N__33793),
            .I(\ALU.r4_RNIKUMQ8_1Z0Z_8 ));
    InMux I__6544 (
            .O(N__33790),
            .I(bfn_10_10_0_));
    InMux I__6543 (
            .O(N__33787),
            .I(\ALU.un2_addsub_cry_8 ));
    InMux I__6542 (
            .O(N__33784),
            .I(N__33780));
    InMux I__6541 (
            .O(N__33783),
            .I(N__33777));
    LocalMux I__6540 (
            .O(N__33780),
            .I(N__33774));
    LocalMux I__6539 (
            .O(N__33777),
            .I(N__33771));
    Span4Mux_v I__6538 (
            .O(N__33774),
            .I(N__33767));
    Span4Mux_h I__6537 (
            .O(N__33771),
            .I(N__33764));
    InMux I__6536 (
            .O(N__33770),
            .I(N__33761));
    Span4Mux_h I__6535 (
            .O(N__33767),
            .I(N__33758));
    Span4Mux_v I__6534 (
            .O(N__33764),
            .I(N__33753));
    LocalMux I__6533 (
            .O(N__33761),
            .I(N__33753));
    Span4Mux_v I__6532 (
            .O(N__33758),
            .I(N__33748));
    Span4Mux_h I__6531 (
            .O(N__33753),
            .I(N__33748));
    Odrv4 I__6530 (
            .O(N__33748),
            .I(r5_6));
    InMux I__6529 (
            .O(N__33745),
            .I(N__33739));
    InMux I__6528 (
            .O(N__33744),
            .I(N__33739));
    LocalMux I__6527 (
            .O(N__33739),
            .I(N__33735));
    InMux I__6526 (
            .O(N__33738),
            .I(N__33732));
    Odrv4 I__6525 (
            .O(N__33735),
            .I(r5_7));
    LocalMux I__6524 (
            .O(N__33732),
            .I(r5_7));
    CascadeMux I__6523 (
            .O(N__33727),
            .I(N__33724));
    InMux I__6522 (
            .O(N__33724),
            .I(N__33721));
    LocalMux I__6521 (
            .O(N__33721),
            .I(N__33718));
    Span4Mux_s2_v I__6520 (
            .O(N__33718),
            .I(N__33713));
    InMux I__6519 (
            .O(N__33717),
            .I(N__33710));
    InMux I__6518 (
            .O(N__33716),
            .I(N__33707));
    Span4Mux_h I__6517 (
            .O(N__33713),
            .I(N__33704));
    LocalMux I__6516 (
            .O(N__33710),
            .I(N__33699));
    LocalMux I__6515 (
            .O(N__33707),
            .I(N__33699));
    Span4Mux_v I__6514 (
            .O(N__33704),
            .I(N__33696));
    Odrv12 I__6513 (
            .O(N__33699),
            .I(r5_8));
    Odrv4 I__6512 (
            .O(N__33696),
            .I(r5_8));
    InMux I__6511 (
            .O(N__33691),
            .I(N__33688));
    LocalMux I__6510 (
            .O(N__33688),
            .I(N__33684));
    InMux I__6509 (
            .O(N__33687),
            .I(N__33681));
    Span4Mux_h I__6508 (
            .O(N__33684),
            .I(N__33677));
    LocalMux I__6507 (
            .O(N__33681),
            .I(N__33674));
    InMux I__6506 (
            .O(N__33680),
            .I(N__33671));
    Odrv4 I__6505 (
            .O(N__33677),
            .I(r5_9));
    Odrv12 I__6504 (
            .O(N__33674),
            .I(r5_9));
    LocalMux I__6503 (
            .O(N__33671),
            .I(r5_9));
    InMux I__6502 (
            .O(N__33664),
            .I(N__33660));
    InMux I__6501 (
            .O(N__33663),
            .I(N__33657));
    LocalMux I__6500 (
            .O(N__33660),
            .I(N__33654));
    LocalMux I__6499 (
            .O(N__33657),
            .I(N__33650));
    Span4Mux_v I__6498 (
            .O(N__33654),
            .I(N__33647));
    InMux I__6497 (
            .O(N__33653),
            .I(N__33644));
    Span4Mux_h I__6496 (
            .O(N__33650),
            .I(N__33641));
    Odrv4 I__6495 (
            .O(N__33647),
            .I(r5_1));
    LocalMux I__6494 (
            .O(N__33644),
            .I(r5_1));
    Odrv4 I__6493 (
            .O(N__33641),
            .I(r5_1));
    InMux I__6492 (
            .O(N__33634),
            .I(N__33631));
    LocalMux I__6491 (
            .O(N__33631),
            .I(N__33628));
    Span4Mux_v I__6490 (
            .O(N__33628),
            .I(N__33623));
    InMux I__6489 (
            .O(N__33627),
            .I(N__33620));
    InMux I__6488 (
            .O(N__33626),
            .I(N__33617));
    Odrv4 I__6487 (
            .O(N__33623),
            .I(r5_2));
    LocalMux I__6486 (
            .O(N__33620),
            .I(r5_2));
    LocalMux I__6485 (
            .O(N__33617),
            .I(r5_2));
    InMux I__6484 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__6483 (
            .O(N__33607),
            .I(N__33604));
    Span4Mux_v I__6482 (
            .O(N__33604),
            .I(N__33600));
    CascadeMux I__6481 (
            .O(N__33603),
            .I(N__33597));
    Span4Mux_h I__6480 (
            .O(N__33600),
            .I(N__33594));
    InMux I__6479 (
            .O(N__33597),
            .I(N__33591));
    Span4Mux_v I__6478 (
            .O(N__33594),
            .I(N__33586));
    LocalMux I__6477 (
            .O(N__33591),
            .I(N__33586));
    Span4Mux_h I__6476 (
            .O(N__33586),
            .I(N__33582));
    InMux I__6475 (
            .O(N__33585),
            .I(N__33579));
    Odrv4 I__6474 (
            .O(N__33582),
            .I(r5_3));
    LocalMux I__6473 (
            .O(N__33579),
            .I(r5_3));
    InMux I__6472 (
            .O(N__33574),
            .I(N__33571));
    LocalMux I__6471 (
            .O(N__33571),
            .I(N__33568));
    Span4Mux_v I__6470 (
            .O(N__33568),
            .I(N__33565));
    Span4Mux_h I__6469 (
            .O(N__33565),
            .I(N__33562));
    Span4Mux_h I__6468 (
            .O(N__33562),
            .I(N__33557));
    InMux I__6467 (
            .O(N__33561),
            .I(N__33554));
    InMux I__6466 (
            .O(N__33560),
            .I(N__33551));
    Odrv4 I__6465 (
            .O(N__33557),
            .I(r5_4));
    LocalMux I__6464 (
            .O(N__33554),
            .I(r5_4));
    LocalMux I__6463 (
            .O(N__33551),
            .I(r5_4));
    CascadeMux I__6462 (
            .O(N__33544),
            .I(N__33541));
    InMux I__6461 (
            .O(N__33541),
            .I(N__33538));
    LocalMux I__6460 (
            .O(N__33538),
            .I(N__33535));
    Span4Mux_v I__6459 (
            .O(N__33535),
            .I(N__33532));
    Span4Mux_v I__6458 (
            .O(N__33532),
            .I(N__33529));
    Span4Mux_h I__6457 (
            .O(N__33529),
            .I(N__33526));
    Odrv4 I__6456 (
            .O(N__33526),
            .I(\ALU.r4_RNIUES39Z0Z_1 ));
    InMux I__6455 (
            .O(N__33523),
            .I(N__33520));
    LocalMux I__6454 (
            .O(N__33520),
            .I(N__33517));
    Span4Mux_h I__6453 (
            .O(N__33517),
            .I(N__33514));
    Odrv4 I__6452 (
            .O(N__33514),
            .I(\ALU.b_3_ns_1_0 ));
    InMux I__6451 (
            .O(N__33511),
            .I(N__33508));
    LocalMux I__6450 (
            .O(N__33508),
            .I(N__33504));
    InMux I__6449 (
            .O(N__33507),
            .I(N__33501));
    Span4Mux_h I__6448 (
            .O(N__33504),
            .I(N__33498));
    LocalMux I__6447 (
            .O(N__33501),
            .I(N__33494));
    Span4Mux_h I__6446 (
            .O(N__33498),
            .I(N__33491));
    InMux I__6445 (
            .O(N__33497),
            .I(N__33488));
    Span4Mux_h I__6444 (
            .O(N__33494),
            .I(N__33485));
    Odrv4 I__6443 (
            .O(N__33491),
            .I(r0_4));
    LocalMux I__6442 (
            .O(N__33488),
            .I(r0_4));
    Odrv4 I__6441 (
            .O(N__33485),
            .I(r0_4));
    InMux I__6440 (
            .O(N__33478),
            .I(N__33475));
    LocalMux I__6439 (
            .O(N__33475),
            .I(N__33472));
    Span4Mux_v I__6438 (
            .O(N__33472),
            .I(N__33469));
    Span4Mux_h I__6437 (
            .O(N__33469),
            .I(N__33464));
    CascadeMux I__6436 (
            .O(N__33468),
            .I(N__33461));
    InMux I__6435 (
            .O(N__33467),
            .I(N__33458));
    Span4Mux_h I__6434 (
            .O(N__33464),
            .I(N__33455));
    InMux I__6433 (
            .O(N__33461),
            .I(N__33452));
    LocalMux I__6432 (
            .O(N__33458),
            .I(N__33449));
    Odrv4 I__6431 (
            .O(N__33455),
            .I(r1_4));
    LocalMux I__6430 (
            .O(N__33452),
            .I(r1_4));
    Odrv12 I__6429 (
            .O(N__33449),
            .I(r1_4));
    CascadeMux I__6428 (
            .O(N__33442),
            .I(\ALU.b_3_ns_1_4_cascade_ ));
    InMux I__6427 (
            .O(N__33439),
            .I(N__33435));
    InMux I__6426 (
            .O(N__33438),
            .I(N__33432));
    LocalMux I__6425 (
            .O(N__33435),
            .I(N__33429));
    LocalMux I__6424 (
            .O(N__33432),
            .I(N__33426));
    Span4Mux_v I__6423 (
            .O(N__33429),
            .I(N__33421));
    Span4Mux_v I__6422 (
            .O(N__33426),
            .I(N__33421));
    Odrv4 I__6421 (
            .O(N__33421),
            .I(\ALU.r4_RNISLNE1Z0Z_4 ));
    InMux I__6420 (
            .O(N__33418),
            .I(N__33415));
    LocalMux I__6419 (
            .O(N__33415),
            .I(N__33412));
    Span4Mux_h I__6418 (
            .O(N__33412),
            .I(N__33408));
    InMux I__6417 (
            .O(N__33411),
            .I(N__33404));
    Span4Mux_h I__6416 (
            .O(N__33408),
            .I(N__33401));
    InMux I__6415 (
            .O(N__33407),
            .I(N__33398));
    LocalMux I__6414 (
            .O(N__33404),
            .I(N__33395));
    Odrv4 I__6413 (
            .O(N__33401),
            .I(r0_2));
    LocalMux I__6412 (
            .O(N__33398),
            .I(r0_2));
    Odrv4 I__6411 (
            .O(N__33395),
            .I(r0_2));
    InMux I__6410 (
            .O(N__33388),
            .I(N__33385));
    LocalMux I__6409 (
            .O(N__33385),
            .I(N__33381));
    CascadeMux I__6408 (
            .O(N__33384),
            .I(N__33377));
    Span4Mux_v I__6407 (
            .O(N__33381),
            .I(N__33374));
    CascadeMux I__6406 (
            .O(N__33380),
            .I(N__33371));
    InMux I__6405 (
            .O(N__33377),
            .I(N__33368));
    Span4Mux_h I__6404 (
            .O(N__33374),
            .I(N__33365));
    InMux I__6403 (
            .O(N__33371),
            .I(N__33362));
    LocalMux I__6402 (
            .O(N__33368),
            .I(N__33359));
    Odrv4 I__6401 (
            .O(N__33365),
            .I(r1_2));
    LocalMux I__6400 (
            .O(N__33362),
            .I(r1_2));
    Odrv12 I__6399 (
            .O(N__33359),
            .I(r1_2));
    CascadeMux I__6398 (
            .O(N__33352),
            .I(\ALU.b_3_ns_1_2_cascade_ ));
    InMux I__6397 (
            .O(N__33349),
            .I(N__33344));
    InMux I__6396 (
            .O(N__33348),
            .I(N__33341));
    InMux I__6395 (
            .O(N__33347),
            .I(N__33337));
    LocalMux I__6394 (
            .O(N__33344),
            .I(N__33334));
    LocalMux I__6393 (
            .O(N__33341),
            .I(N__33331));
    InMux I__6392 (
            .O(N__33340),
            .I(N__33328));
    LocalMux I__6391 (
            .O(N__33337),
            .I(N__33325));
    Span4Mux_h I__6390 (
            .O(N__33334),
            .I(N__33322));
    Span12Mux_s8_h I__6389 (
            .O(N__33331),
            .I(N__33319));
    LocalMux I__6388 (
            .O(N__33328),
            .I(N__33316));
    Span4Mux_h I__6387 (
            .O(N__33325),
            .I(N__33313));
    Odrv4 I__6386 (
            .O(N__33322),
            .I(\ALU.r4_RNIKDNE1Z0Z_2 ));
    Odrv12 I__6385 (
            .O(N__33319),
            .I(\ALU.r4_RNIKDNE1Z0Z_2 ));
    Odrv4 I__6384 (
            .O(N__33316),
            .I(\ALU.r4_RNIKDNE1Z0Z_2 ));
    Odrv4 I__6383 (
            .O(N__33313),
            .I(\ALU.r4_RNIKDNE1Z0Z_2 ));
    CascadeMux I__6382 (
            .O(N__33304),
            .I(N__33300));
    InMux I__6381 (
            .O(N__33303),
            .I(N__33292));
    InMux I__6380 (
            .O(N__33300),
            .I(N__33285));
    InMux I__6379 (
            .O(N__33299),
            .I(N__33276));
    InMux I__6378 (
            .O(N__33298),
            .I(N__33276));
    InMux I__6377 (
            .O(N__33297),
            .I(N__33276));
    InMux I__6376 (
            .O(N__33296),
            .I(N__33276));
    InMux I__6375 (
            .O(N__33295),
            .I(N__33273));
    LocalMux I__6374 (
            .O(N__33292),
            .I(N__33270));
    InMux I__6373 (
            .O(N__33291),
            .I(N__33261));
    InMux I__6372 (
            .O(N__33290),
            .I(N__33261));
    InMux I__6371 (
            .O(N__33289),
            .I(N__33261));
    InMux I__6370 (
            .O(N__33288),
            .I(N__33261));
    LocalMux I__6369 (
            .O(N__33285),
            .I(N__33258));
    LocalMux I__6368 (
            .O(N__33276),
            .I(N__33255));
    LocalMux I__6367 (
            .O(N__33273),
            .I(b_fastZ0Z_2));
    Odrv4 I__6366 (
            .O(N__33270),
            .I(b_fastZ0Z_2));
    LocalMux I__6365 (
            .O(N__33261),
            .I(b_fastZ0Z_2));
    Odrv4 I__6364 (
            .O(N__33258),
            .I(b_fastZ0Z_2));
    Odrv12 I__6363 (
            .O(N__33255),
            .I(b_fastZ0Z_2));
    InMux I__6362 (
            .O(N__33244),
            .I(N__33241));
    LocalMux I__6361 (
            .O(N__33241),
            .I(N__33238));
    Span4Mux_v I__6360 (
            .O(N__33238),
            .I(N__33234));
    CascadeMux I__6359 (
            .O(N__33237),
            .I(N__33230));
    Sp12to4 I__6358 (
            .O(N__33234),
            .I(N__33227));
    CascadeMux I__6357 (
            .O(N__33233),
            .I(N__33224));
    InMux I__6356 (
            .O(N__33230),
            .I(N__33221));
    Span12Mux_s8_h I__6355 (
            .O(N__33227),
            .I(N__33218));
    InMux I__6354 (
            .O(N__33224),
            .I(N__33215));
    LocalMux I__6353 (
            .O(N__33221),
            .I(N__33212));
    Odrv12 I__6352 (
            .O(N__33218),
            .I(r1_3));
    LocalMux I__6351 (
            .O(N__33215),
            .I(r1_3));
    Odrv4 I__6350 (
            .O(N__33212),
            .I(r1_3));
    InMux I__6349 (
            .O(N__33205),
            .I(N__33197));
    InMux I__6348 (
            .O(N__33204),
            .I(N__33197));
    InMux I__6347 (
            .O(N__33203),
            .I(N__33194));
    InMux I__6346 (
            .O(N__33202),
            .I(N__33191));
    LocalMux I__6345 (
            .O(N__33197),
            .I(N__33188));
    LocalMux I__6344 (
            .O(N__33194),
            .I(N__33185));
    LocalMux I__6343 (
            .O(N__33191),
            .I(N__33178));
    Span4Mux_v I__6342 (
            .O(N__33188),
            .I(N__33175));
    Span4Mux_h I__6341 (
            .O(N__33185),
            .I(N__33171));
    InMux I__6340 (
            .O(N__33184),
            .I(N__33168));
    InMux I__6339 (
            .O(N__33183),
            .I(N__33161));
    InMux I__6338 (
            .O(N__33182),
            .I(N__33161));
    InMux I__6337 (
            .O(N__33181),
            .I(N__33161));
    Span4Mux_h I__6336 (
            .O(N__33178),
            .I(N__33156));
    Span4Mux_h I__6335 (
            .O(N__33175),
            .I(N__33156));
    InMux I__6334 (
            .O(N__33174),
            .I(N__33153));
    Odrv4 I__6333 (
            .O(N__33171),
            .I(b_fastZ0Z_0));
    LocalMux I__6332 (
            .O(N__33168),
            .I(b_fastZ0Z_0));
    LocalMux I__6331 (
            .O(N__33161),
            .I(b_fastZ0Z_0));
    Odrv4 I__6330 (
            .O(N__33156),
            .I(b_fastZ0Z_0));
    LocalMux I__6329 (
            .O(N__33153),
            .I(b_fastZ0Z_0));
    InMux I__6328 (
            .O(N__33142),
            .I(N__33132));
    InMux I__6327 (
            .O(N__33141),
            .I(N__33127));
    InMux I__6326 (
            .O(N__33140),
            .I(N__33127));
    InMux I__6325 (
            .O(N__33139),
            .I(N__33124));
    InMux I__6324 (
            .O(N__33138),
            .I(N__33121));
    InMux I__6323 (
            .O(N__33137),
            .I(N__33114));
    InMux I__6322 (
            .O(N__33136),
            .I(N__33114));
    InMux I__6321 (
            .O(N__33135),
            .I(N__33114));
    LocalMux I__6320 (
            .O(N__33132),
            .I(N__33108));
    LocalMux I__6319 (
            .O(N__33127),
            .I(N__33105));
    LocalMux I__6318 (
            .O(N__33124),
            .I(N__33102));
    LocalMux I__6317 (
            .O(N__33121),
            .I(N__33097));
    LocalMux I__6316 (
            .O(N__33114),
            .I(N__33097));
    InMux I__6315 (
            .O(N__33113),
            .I(N__33094));
    InMux I__6314 (
            .O(N__33112),
            .I(N__33091));
    InMux I__6313 (
            .O(N__33111),
            .I(N__33088));
    Span4Mux_v I__6312 (
            .O(N__33108),
            .I(N__33083));
    Span4Mux_h I__6311 (
            .O(N__33105),
            .I(N__33083));
    Span4Mux_h I__6310 (
            .O(N__33102),
            .I(N__33080));
    Span4Mux_h I__6309 (
            .O(N__33097),
            .I(N__33077));
    LocalMux I__6308 (
            .O(N__33094),
            .I(b_2_repZ0Z1));
    LocalMux I__6307 (
            .O(N__33091),
            .I(b_2_repZ0Z1));
    LocalMux I__6306 (
            .O(N__33088),
            .I(b_2_repZ0Z1));
    Odrv4 I__6305 (
            .O(N__33083),
            .I(b_2_repZ0Z1));
    Odrv4 I__6304 (
            .O(N__33080),
            .I(b_2_repZ0Z1));
    Odrv4 I__6303 (
            .O(N__33077),
            .I(b_2_repZ0Z1));
    InMux I__6302 (
            .O(N__33064),
            .I(N__33061));
    LocalMux I__6301 (
            .O(N__33061),
            .I(N__33058));
    Span4Mux_v I__6300 (
            .O(N__33058),
            .I(N__33053));
    InMux I__6299 (
            .O(N__33057),
            .I(N__33048));
    InMux I__6298 (
            .O(N__33056),
            .I(N__33048));
    Span4Mux_h I__6297 (
            .O(N__33053),
            .I(N__33045));
    LocalMux I__6296 (
            .O(N__33048),
            .I(r4_3));
    Odrv4 I__6295 (
            .O(N__33045),
            .I(r4_3));
    CascadeMux I__6294 (
            .O(N__33040),
            .I(\ALU.b_3_ns_1_3_cascade_ ));
    InMux I__6293 (
            .O(N__33037),
            .I(N__33031));
    InMux I__6292 (
            .O(N__33036),
            .I(N__33031));
    LocalMux I__6291 (
            .O(N__33031),
            .I(N__33027));
    InMux I__6290 (
            .O(N__33030),
            .I(N__33024));
    Span4Mux_v I__6289 (
            .O(N__33027),
            .I(N__33021));
    LocalMux I__6288 (
            .O(N__33024),
            .I(N__33018));
    Span4Mux_h I__6287 (
            .O(N__33021),
            .I(N__33013));
    Span4Mux_v I__6286 (
            .O(N__33018),
            .I(N__33013));
    Odrv4 I__6285 (
            .O(N__33013),
            .I(\ALU.r4_RNIOHNE1Z0Z_3 ));
    InMux I__6284 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__6283 (
            .O(N__33007),
            .I(N__33004));
    Span4Mux_v I__6282 (
            .O(N__33004),
            .I(N__33001));
    Span4Mux_v I__6281 (
            .O(N__33001),
            .I(N__32998));
    Odrv4 I__6280 (
            .O(N__32998),
            .I(\ALU.rshift_10 ));
    InMux I__6279 (
            .O(N__32995),
            .I(N__32992));
    LocalMux I__6278 (
            .O(N__32992),
            .I(N__32989));
    Span4Mux_h I__6277 (
            .O(N__32989),
            .I(N__32986));
    Odrv4 I__6276 (
            .O(N__32986),
            .I(\ALU.madd_76_0 ));
    CascadeMux I__6275 (
            .O(N__32983),
            .I(\ALU.lshift_3_ns_1_11_cascade_ ));
    CascadeMux I__6274 (
            .O(N__32980),
            .I(N__32977));
    InMux I__6273 (
            .O(N__32977),
            .I(N__32974));
    LocalMux I__6272 (
            .O(N__32974),
            .I(\ALU.un9_addsub_axb_4 ));
    InMux I__6271 (
            .O(N__32971),
            .I(N__32968));
    LocalMux I__6270 (
            .O(N__32968),
            .I(N__32965));
    Span4Mux_h I__6269 (
            .O(N__32965),
            .I(N__32962));
    Odrv4 I__6268 (
            .O(N__32962),
            .I(\ALU.lshift_3_ns_1_9 ));
    InMux I__6267 (
            .O(N__32959),
            .I(N__32956));
    LocalMux I__6266 (
            .O(N__32956),
            .I(N__32951));
    InMux I__6265 (
            .O(N__32955),
            .I(N__32948));
    InMux I__6264 (
            .O(N__32954),
            .I(N__32945));
    Span4Mux_h I__6263 (
            .O(N__32951),
            .I(N__32940));
    LocalMux I__6262 (
            .O(N__32948),
            .I(N__32940));
    LocalMux I__6261 (
            .O(N__32945),
            .I(r1_1));
    Odrv4 I__6260 (
            .O(N__32940),
            .I(r1_1));
    InMux I__6259 (
            .O(N__32935),
            .I(N__32932));
    LocalMux I__6258 (
            .O(N__32932),
            .I(N__32929));
    Span4Mux_h I__6257 (
            .O(N__32929),
            .I(N__32926));
    Odrv4 I__6256 (
            .O(N__32926),
            .I(\ALU.r0_RNIE5LHZ0Z_1 ));
    CascadeMux I__6255 (
            .O(N__32923),
            .I(\ALU.rshift_3_ns_1_3_cascade_ ));
    CascadeMux I__6254 (
            .O(N__32920),
            .I(\ALU.r0_12_prm_8_3_c_RNOZ0Z_3_cascade_ ));
    InMux I__6253 (
            .O(N__32917),
            .I(N__32914));
    LocalMux I__6252 (
            .O(N__32914),
            .I(N__32911));
    Span4Mux_v I__6251 (
            .O(N__32911),
            .I(N__32907));
    InMux I__6250 (
            .O(N__32910),
            .I(N__32904));
    Span4Mux_v I__6249 (
            .O(N__32907),
            .I(N__32901));
    LocalMux I__6248 (
            .O(N__32904),
            .I(\ALU.r5_RNI67NNKZ0Z_10 ));
    Odrv4 I__6247 (
            .O(N__32901),
            .I(\ALU.r5_RNI67NNKZ0Z_10 ));
    InMux I__6246 (
            .O(N__32896),
            .I(N__32888));
    CascadeMux I__6245 (
            .O(N__32895),
            .I(N__32884));
    CascadeMux I__6244 (
            .O(N__32894),
            .I(N__32880));
    InMux I__6243 (
            .O(N__32893),
            .I(N__32877));
    InMux I__6242 (
            .O(N__32892),
            .I(N__32874));
    InMux I__6241 (
            .O(N__32891),
            .I(N__32871));
    LocalMux I__6240 (
            .O(N__32888),
            .I(N__32868));
    InMux I__6239 (
            .O(N__32887),
            .I(N__32865));
    InMux I__6238 (
            .O(N__32884),
            .I(N__32856));
    InMux I__6237 (
            .O(N__32883),
            .I(N__32856));
    InMux I__6236 (
            .O(N__32880),
            .I(N__32853));
    LocalMux I__6235 (
            .O(N__32877),
            .I(N__32842));
    LocalMux I__6234 (
            .O(N__32874),
            .I(N__32842));
    LocalMux I__6233 (
            .O(N__32871),
            .I(N__32842));
    Span4Mux_v I__6232 (
            .O(N__32868),
            .I(N__32842));
    LocalMux I__6231 (
            .O(N__32865),
            .I(N__32842));
    CascadeMux I__6230 (
            .O(N__32864),
            .I(N__32838));
    CascadeMux I__6229 (
            .O(N__32863),
            .I(N__32835));
    InMux I__6228 (
            .O(N__32862),
            .I(N__32831));
    InMux I__6227 (
            .O(N__32861),
            .I(N__32827));
    LocalMux I__6226 (
            .O(N__32856),
            .I(N__32824));
    LocalMux I__6225 (
            .O(N__32853),
            .I(N__32821));
    Span4Mux_v I__6224 (
            .O(N__32842),
            .I(N__32818));
    CascadeMux I__6223 (
            .O(N__32841),
            .I(N__32812));
    InMux I__6222 (
            .O(N__32838),
            .I(N__32807));
    InMux I__6221 (
            .O(N__32835),
            .I(N__32807));
    InMux I__6220 (
            .O(N__32834),
            .I(N__32804));
    LocalMux I__6219 (
            .O(N__32831),
            .I(N__32801));
    InMux I__6218 (
            .O(N__32830),
            .I(N__32798));
    LocalMux I__6217 (
            .O(N__32827),
            .I(N__32795));
    Span4Mux_s2_h I__6216 (
            .O(N__32824),
            .I(N__32788));
    Span4Mux_v I__6215 (
            .O(N__32821),
            .I(N__32788));
    Span4Mux_s2_h I__6214 (
            .O(N__32818),
            .I(N__32788));
    InMux I__6213 (
            .O(N__32817),
            .I(N__32781));
    InMux I__6212 (
            .O(N__32816),
            .I(N__32781));
    InMux I__6211 (
            .O(N__32815),
            .I(N__32781));
    InMux I__6210 (
            .O(N__32812),
            .I(N__32778));
    LocalMux I__6209 (
            .O(N__32807),
            .I(N__32775));
    LocalMux I__6208 (
            .O(N__32804),
            .I(N__32768));
    Span12Mux_h I__6207 (
            .O(N__32801),
            .I(N__32768));
    LocalMux I__6206 (
            .O(N__32798),
            .I(N__32768));
    Span4Mux_h I__6205 (
            .O(N__32795),
            .I(N__32763));
    Span4Mux_h I__6204 (
            .O(N__32788),
            .I(N__32763));
    LocalMux I__6203 (
            .O(N__32781),
            .I(bZ0Z_1));
    LocalMux I__6202 (
            .O(N__32778),
            .I(bZ0Z_1));
    Odrv12 I__6201 (
            .O(N__32775),
            .I(bZ0Z_1));
    Odrv12 I__6200 (
            .O(N__32768),
            .I(bZ0Z_1));
    Odrv4 I__6199 (
            .O(N__32763),
            .I(bZ0Z_1));
    InMux I__6198 (
            .O(N__32752),
            .I(N__32749));
    LocalMux I__6197 (
            .O(N__32749),
            .I(N__32745));
    InMux I__6196 (
            .O(N__32748),
            .I(N__32741));
    Span4Mux_v I__6195 (
            .O(N__32745),
            .I(N__32738));
    InMux I__6194 (
            .O(N__32744),
            .I(N__32735));
    LocalMux I__6193 (
            .O(N__32741),
            .I(N__32732));
    Span4Mux_h I__6192 (
            .O(N__32738),
            .I(N__32729));
    LocalMux I__6191 (
            .O(N__32735),
            .I(N__32726));
    Odrv12 I__6190 (
            .O(N__32732),
            .I(\ALU.r6_RNI6TET1Z0Z_0 ));
    Odrv4 I__6189 (
            .O(N__32729),
            .I(\ALU.r6_RNI6TET1Z0Z_0 ));
    Odrv4 I__6188 (
            .O(N__32726),
            .I(\ALU.r6_RNI6TET1Z0Z_0 ));
    InMux I__6187 (
            .O(N__32719),
            .I(N__32715));
    InMux I__6186 (
            .O(N__32718),
            .I(N__32712));
    LocalMux I__6185 (
            .O(N__32715),
            .I(N__32709));
    LocalMux I__6184 (
            .O(N__32712),
            .I(N__32705));
    Span4Mux_h I__6183 (
            .O(N__32709),
            .I(N__32702));
    InMux I__6182 (
            .O(N__32708),
            .I(N__32699));
    Odrv12 I__6181 (
            .O(N__32705),
            .I(\ALU.r4_RNIC5NE1Z0Z_0 ));
    Odrv4 I__6180 (
            .O(N__32702),
            .I(\ALU.r4_RNIC5NE1Z0Z_0 ));
    LocalMux I__6179 (
            .O(N__32699),
            .I(\ALU.r4_RNIC5NE1Z0Z_0 ));
    InMux I__6178 (
            .O(N__32692),
            .I(N__32686));
    InMux I__6177 (
            .O(N__32691),
            .I(N__32686));
    LocalMux I__6176 (
            .O(N__32686),
            .I(N__32681));
    InMux I__6175 (
            .O(N__32685),
            .I(N__32678));
    InMux I__6174 (
            .O(N__32684),
            .I(N__32672));
    Span4Mux_s1_v I__6173 (
            .O(N__32681),
            .I(N__32667));
    LocalMux I__6172 (
            .O(N__32678),
            .I(N__32667));
    InMux I__6171 (
            .O(N__32677),
            .I(N__32660));
    InMux I__6170 (
            .O(N__32676),
            .I(N__32660));
    InMux I__6169 (
            .O(N__32675),
            .I(N__32657));
    LocalMux I__6168 (
            .O(N__32672),
            .I(N__32652));
    Span4Mux_h I__6167 (
            .O(N__32667),
            .I(N__32649));
    InMux I__6166 (
            .O(N__32666),
            .I(N__32646));
    InMux I__6165 (
            .O(N__32665),
            .I(N__32643));
    LocalMux I__6164 (
            .O(N__32660),
            .I(N__32638));
    LocalMux I__6163 (
            .O(N__32657),
            .I(N__32638));
    InMux I__6162 (
            .O(N__32656),
            .I(N__32635));
    InMux I__6161 (
            .O(N__32655),
            .I(N__32632));
    Span4Mux_v I__6160 (
            .O(N__32652),
            .I(N__32629));
    Span4Mux_v I__6159 (
            .O(N__32649),
            .I(N__32624));
    LocalMux I__6158 (
            .O(N__32646),
            .I(N__32624));
    LocalMux I__6157 (
            .O(N__32643),
            .I(N__32621));
    Span4Mux_h I__6156 (
            .O(N__32638),
            .I(N__32616));
    LocalMux I__6155 (
            .O(N__32635),
            .I(N__32616));
    LocalMux I__6154 (
            .O(N__32632),
            .I(N__32613));
    Sp12to4 I__6153 (
            .O(N__32629),
            .I(N__32610));
    Span4Mux_h I__6152 (
            .O(N__32624),
            .I(N__32605));
    Span4Mux_v I__6151 (
            .O(N__32621),
            .I(N__32605));
    Span4Mux_h I__6150 (
            .O(N__32616),
            .I(N__32602));
    Odrv12 I__6149 (
            .O(N__32613),
            .I(\ALU.r6_RNIBF8D2Z0Z_2 ));
    Odrv12 I__6148 (
            .O(N__32610),
            .I(\ALU.r6_RNIBF8D2Z0Z_2 ));
    Odrv4 I__6147 (
            .O(N__32605),
            .I(\ALU.r6_RNIBF8D2Z0Z_2 ));
    Odrv4 I__6146 (
            .O(N__32602),
            .I(\ALU.r6_RNIBF8D2Z0Z_2 ));
    InMux I__6145 (
            .O(N__32593),
            .I(N__32586));
    CascadeMux I__6144 (
            .O(N__32592),
            .I(N__32583));
    CascadeMux I__6143 (
            .O(N__32591),
            .I(N__32580));
    InMux I__6142 (
            .O(N__32590),
            .I(N__32575));
    InMux I__6141 (
            .O(N__32589),
            .I(N__32571));
    LocalMux I__6140 (
            .O(N__32586),
            .I(N__32567));
    InMux I__6139 (
            .O(N__32583),
            .I(N__32564));
    InMux I__6138 (
            .O(N__32580),
            .I(N__32559));
    InMux I__6137 (
            .O(N__32579),
            .I(N__32559));
    InMux I__6136 (
            .O(N__32578),
            .I(N__32556));
    LocalMux I__6135 (
            .O(N__32575),
            .I(N__32553));
    InMux I__6134 (
            .O(N__32574),
            .I(N__32550));
    LocalMux I__6133 (
            .O(N__32571),
            .I(N__32545));
    InMux I__6132 (
            .O(N__32570),
            .I(N__32542));
    Span4Mux_v I__6131 (
            .O(N__32567),
            .I(N__32537));
    LocalMux I__6130 (
            .O(N__32564),
            .I(N__32537));
    LocalMux I__6129 (
            .O(N__32559),
            .I(N__32534));
    LocalMux I__6128 (
            .O(N__32556),
            .I(N__32531));
    Span4Mux_h I__6127 (
            .O(N__32553),
            .I(N__32526));
    LocalMux I__6126 (
            .O(N__32550),
            .I(N__32526));
    InMux I__6125 (
            .O(N__32549),
            .I(N__32521));
    InMux I__6124 (
            .O(N__32548),
            .I(N__32521));
    Span4Mux_v I__6123 (
            .O(N__32545),
            .I(N__32518));
    LocalMux I__6122 (
            .O(N__32542),
            .I(N__32515));
    Span4Mux_h I__6121 (
            .O(N__32537),
            .I(N__32510));
    Span4Mux_v I__6120 (
            .O(N__32534),
            .I(N__32510));
    Span4Mux_h I__6119 (
            .O(N__32531),
            .I(N__32507));
    Span4Mux_v I__6118 (
            .O(N__32526),
            .I(N__32504));
    LocalMux I__6117 (
            .O(N__32521),
            .I(N__32501));
    Span4Mux_h I__6116 (
            .O(N__32518),
            .I(N__32498));
    Span12Mux_s8_h I__6115 (
            .O(N__32515),
            .I(N__32495));
    Span4Mux_v I__6114 (
            .O(N__32510),
            .I(N__32492));
    Span4Mux_h I__6113 (
            .O(N__32507),
            .I(N__32487));
    Span4Mux_h I__6112 (
            .O(N__32504),
            .I(N__32487));
    Odrv12 I__6111 (
            .O(N__32501),
            .I(\ALU.r4_RNIHM992Z0Z_2 ));
    Odrv4 I__6110 (
            .O(N__32498),
            .I(\ALU.r4_RNIHM992Z0Z_2 ));
    Odrv12 I__6109 (
            .O(N__32495),
            .I(\ALU.r4_RNIHM992Z0Z_2 ));
    Odrv4 I__6108 (
            .O(N__32492),
            .I(\ALU.r4_RNIHM992Z0Z_2 ));
    Odrv4 I__6107 (
            .O(N__32487),
            .I(\ALU.r4_RNIHM992Z0Z_2 ));
    InMux I__6106 (
            .O(N__32476),
            .I(N__32473));
    LocalMux I__6105 (
            .O(N__32473),
            .I(N__32465));
    InMux I__6104 (
            .O(N__32472),
            .I(N__32461));
    InMux I__6103 (
            .O(N__32471),
            .I(N__32457));
    InMux I__6102 (
            .O(N__32470),
            .I(N__32454));
    InMux I__6101 (
            .O(N__32469),
            .I(N__32448));
    InMux I__6100 (
            .O(N__32468),
            .I(N__32448));
    Span4Mux_s1_v I__6099 (
            .O(N__32465),
            .I(N__32444));
    InMux I__6098 (
            .O(N__32464),
            .I(N__32441));
    LocalMux I__6097 (
            .O(N__32461),
            .I(N__32438));
    InMux I__6096 (
            .O(N__32460),
            .I(N__32435));
    LocalMux I__6095 (
            .O(N__32457),
            .I(N__32432));
    LocalMux I__6094 (
            .O(N__32454),
            .I(N__32429));
    InMux I__6093 (
            .O(N__32453),
            .I(N__32426));
    LocalMux I__6092 (
            .O(N__32448),
            .I(N__32423));
    InMux I__6091 (
            .O(N__32447),
            .I(N__32420));
    Span4Mux_v I__6090 (
            .O(N__32444),
            .I(N__32417));
    LocalMux I__6089 (
            .O(N__32441),
            .I(N__32414));
    Span4Mux_s2_v I__6088 (
            .O(N__32438),
            .I(N__32407));
    LocalMux I__6087 (
            .O(N__32435),
            .I(N__32407));
    Span4Mux_h I__6086 (
            .O(N__32432),
            .I(N__32407));
    Span4Mux_h I__6085 (
            .O(N__32429),
            .I(N__32402));
    LocalMux I__6084 (
            .O(N__32426),
            .I(N__32402));
    Span4Mux_v I__6083 (
            .O(N__32423),
            .I(N__32397));
    LocalMux I__6082 (
            .O(N__32420),
            .I(N__32397));
    Span4Mux_v I__6081 (
            .O(N__32417),
            .I(N__32394));
    Span4Mux_h I__6080 (
            .O(N__32414),
            .I(N__32389));
    Span4Mux_v I__6079 (
            .O(N__32407),
            .I(N__32389));
    Span4Mux_v I__6078 (
            .O(N__32402),
            .I(N__32384));
    Span4Mux_h I__6077 (
            .O(N__32397),
            .I(N__32384));
    Odrv4 I__6076 (
            .O(N__32394),
            .I(\ALU.r6_RNI403D2Z0Z_4 ));
    Odrv4 I__6075 (
            .O(N__32389),
            .I(\ALU.r6_RNI403D2Z0Z_4 ));
    Odrv4 I__6074 (
            .O(N__32384),
            .I(\ALU.r6_RNI403D2Z0Z_4 ));
    InMux I__6073 (
            .O(N__32377),
            .I(N__32369));
    InMux I__6072 (
            .O(N__32376),
            .I(N__32366));
    InMux I__6071 (
            .O(N__32375),
            .I(N__32363));
    CascadeMux I__6070 (
            .O(N__32374),
            .I(N__32357));
    InMux I__6069 (
            .O(N__32373),
            .I(N__32354));
    InMux I__6068 (
            .O(N__32372),
            .I(N__32351));
    LocalMux I__6067 (
            .O(N__32369),
            .I(N__32345));
    LocalMux I__6066 (
            .O(N__32366),
            .I(N__32345));
    LocalMux I__6065 (
            .O(N__32363),
            .I(N__32342));
    InMux I__6064 (
            .O(N__32362),
            .I(N__32339));
    InMux I__6063 (
            .O(N__32361),
            .I(N__32336));
    InMux I__6062 (
            .O(N__32360),
            .I(N__32331));
    InMux I__6061 (
            .O(N__32357),
            .I(N__32331));
    LocalMux I__6060 (
            .O(N__32354),
            .I(N__32328));
    LocalMux I__6059 (
            .O(N__32351),
            .I(N__32325));
    InMux I__6058 (
            .O(N__32350),
            .I(N__32322));
    Span4Mux_v I__6057 (
            .O(N__32345),
            .I(N__32319));
    Span4Mux_h I__6056 (
            .O(N__32342),
            .I(N__32312));
    LocalMux I__6055 (
            .O(N__32339),
            .I(N__32312));
    LocalMux I__6054 (
            .O(N__32336),
            .I(N__32312));
    LocalMux I__6053 (
            .O(N__32331),
            .I(N__32309));
    Span4Mux_h I__6052 (
            .O(N__32328),
            .I(N__32306));
    Span4Mux_v I__6051 (
            .O(N__32325),
            .I(N__32303));
    LocalMux I__6050 (
            .O(N__32322),
            .I(N__32300));
    Span4Mux_h I__6049 (
            .O(N__32319),
            .I(N__32295));
    Span4Mux_v I__6048 (
            .O(N__32312),
            .I(N__32295));
    Span4Mux_h I__6047 (
            .O(N__32309),
            .I(N__32290));
    Span4Mux_v I__6046 (
            .O(N__32306),
            .I(N__32290));
    Span4Mux_h I__6045 (
            .O(N__32303),
            .I(N__32283));
    Span4Mux_v I__6044 (
            .O(N__32300),
            .I(N__32283));
    Span4Mux_v I__6043 (
            .O(N__32295),
            .I(N__32283));
    Odrv4 I__6042 (
            .O(N__32290),
            .I(\ALU.r4_RNIQU992Z0Z_4 ));
    Odrv4 I__6041 (
            .O(N__32283),
            .I(\ALU.r4_RNIQU992Z0Z_4 ));
    CascadeMux I__6040 (
            .O(N__32278),
            .I(N__32273));
    CascadeMux I__6039 (
            .O(N__32277),
            .I(N__32269));
    CascadeMux I__6038 (
            .O(N__32276),
            .I(N__32266));
    InMux I__6037 (
            .O(N__32273),
            .I(N__32258));
    CascadeMux I__6036 (
            .O(N__32272),
            .I(N__32254));
    InMux I__6035 (
            .O(N__32269),
            .I(N__32249));
    InMux I__6034 (
            .O(N__32266),
            .I(N__32249));
    CascadeMux I__6033 (
            .O(N__32265),
            .I(N__32246));
    CascadeMux I__6032 (
            .O(N__32264),
            .I(N__32242));
    CascadeMux I__6031 (
            .O(N__32263),
            .I(N__32239));
    CascadeMux I__6030 (
            .O(N__32262),
            .I(N__32233));
    CascadeMux I__6029 (
            .O(N__32261),
            .I(N__32230));
    LocalMux I__6028 (
            .O(N__32258),
            .I(N__32225));
    CascadeMux I__6027 (
            .O(N__32257),
            .I(N__32220));
    InMux I__6026 (
            .O(N__32254),
            .I(N__32217));
    LocalMux I__6025 (
            .O(N__32249),
            .I(N__32214));
    InMux I__6024 (
            .O(N__32246),
            .I(N__32211));
    InMux I__6023 (
            .O(N__32245),
            .I(N__32206));
    InMux I__6022 (
            .O(N__32242),
            .I(N__32206));
    InMux I__6021 (
            .O(N__32239),
            .I(N__32203));
    CascadeMux I__6020 (
            .O(N__32238),
            .I(N__32196));
    CascadeMux I__6019 (
            .O(N__32237),
            .I(N__32193));
    CascadeMux I__6018 (
            .O(N__32236),
            .I(N__32190));
    InMux I__6017 (
            .O(N__32233),
            .I(N__32187));
    InMux I__6016 (
            .O(N__32230),
            .I(N__32182));
    CascadeMux I__6015 (
            .O(N__32229),
            .I(N__32179));
    CascadeMux I__6014 (
            .O(N__32228),
            .I(N__32175));
    Span4Mux_s2_h I__6013 (
            .O(N__32225),
            .I(N__32170));
    InMux I__6012 (
            .O(N__32224),
            .I(N__32163));
    InMux I__6011 (
            .O(N__32223),
            .I(N__32163));
    InMux I__6010 (
            .O(N__32220),
            .I(N__32163));
    LocalMux I__6009 (
            .O(N__32217),
            .I(N__32156));
    Span4Mux_s2_v I__6008 (
            .O(N__32214),
            .I(N__32156));
    LocalMux I__6007 (
            .O(N__32211),
            .I(N__32149));
    LocalMux I__6006 (
            .O(N__32206),
            .I(N__32149));
    LocalMux I__6005 (
            .O(N__32203),
            .I(N__32149));
    CascadeMux I__6004 (
            .O(N__32202),
            .I(N__32146));
    CascadeMux I__6003 (
            .O(N__32201),
            .I(N__32143));
    CascadeMux I__6002 (
            .O(N__32200),
            .I(N__32140));
    InMux I__6001 (
            .O(N__32199),
            .I(N__32133));
    InMux I__6000 (
            .O(N__32196),
            .I(N__32133));
    InMux I__5999 (
            .O(N__32193),
            .I(N__32133));
    InMux I__5998 (
            .O(N__32190),
            .I(N__32130));
    LocalMux I__5997 (
            .O(N__32187),
            .I(N__32126));
    CascadeMux I__5996 (
            .O(N__32186),
            .I(N__32123));
    CascadeMux I__5995 (
            .O(N__32185),
            .I(N__32120));
    LocalMux I__5994 (
            .O(N__32182),
            .I(N__32117));
    InMux I__5993 (
            .O(N__32179),
            .I(N__32110));
    InMux I__5992 (
            .O(N__32178),
            .I(N__32110));
    InMux I__5991 (
            .O(N__32175),
            .I(N__32110));
    CascadeMux I__5990 (
            .O(N__32174),
            .I(N__32107));
    CascadeMux I__5989 (
            .O(N__32173),
            .I(N__32103));
    Span4Mux_h I__5988 (
            .O(N__32170),
            .I(N__32099));
    LocalMux I__5987 (
            .O(N__32163),
            .I(N__32096));
    InMux I__5986 (
            .O(N__32162),
            .I(N__32091));
    InMux I__5985 (
            .O(N__32161),
            .I(N__32091));
    Span4Mux_v I__5984 (
            .O(N__32156),
            .I(N__32086));
    Span4Mux_v I__5983 (
            .O(N__32149),
            .I(N__32086));
    InMux I__5982 (
            .O(N__32146),
            .I(N__32083));
    InMux I__5981 (
            .O(N__32143),
            .I(N__32078));
    InMux I__5980 (
            .O(N__32140),
            .I(N__32078));
    LocalMux I__5979 (
            .O(N__32133),
            .I(N__32075));
    LocalMux I__5978 (
            .O(N__32130),
            .I(N__32072));
    InMux I__5977 (
            .O(N__32129),
            .I(N__32069));
    Span4Mux_v I__5976 (
            .O(N__32126),
            .I(N__32066));
    InMux I__5975 (
            .O(N__32123),
            .I(N__32063));
    InMux I__5974 (
            .O(N__32120),
            .I(N__32060));
    Span4Mux_s1_v I__5973 (
            .O(N__32117),
            .I(N__32055));
    LocalMux I__5972 (
            .O(N__32110),
            .I(N__32055));
    InMux I__5971 (
            .O(N__32107),
            .I(N__32050));
    InMux I__5970 (
            .O(N__32106),
            .I(N__32050));
    InMux I__5969 (
            .O(N__32103),
            .I(N__32045));
    InMux I__5968 (
            .O(N__32102),
            .I(N__32045));
    Span4Mux_v I__5967 (
            .O(N__32099),
            .I(N__32037));
    Span4Mux_v I__5966 (
            .O(N__32096),
            .I(N__32037));
    LocalMux I__5965 (
            .O(N__32091),
            .I(N__32034));
    Sp12to4 I__5964 (
            .O(N__32086),
            .I(N__32031));
    LocalMux I__5963 (
            .O(N__32083),
            .I(N__32026));
    LocalMux I__5962 (
            .O(N__32078),
            .I(N__32026));
    Span4Mux_v I__5961 (
            .O(N__32075),
            .I(N__32023));
    Span4Mux_h I__5960 (
            .O(N__32072),
            .I(N__32014));
    LocalMux I__5959 (
            .O(N__32069),
            .I(N__32014));
    Span4Mux_h I__5958 (
            .O(N__32066),
            .I(N__32014));
    LocalMux I__5957 (
            .O(N__32063),
            .I(N__32014));
    LocalMux I__5956 (
            .O(N__32060),
            .I(N__32011));
    Span4Mux_h I__5955 (
            .O(N__32055),
            .I(N__32004));
    LocalMux I__5954 (
            .O(N__32050),
            .I(N__32004));
    LocalMux I__5953 (
            .O(N__32045),
            .I(N__32004));
    InMux I__5952 (
            .O(N__32044),
            .I(N__31997));
    InMux I__5951 (
            .O(N__32043),
            .I(N__31997));
    InMux I__5950 (
            .O(N__32042),
            .I(N__31997));
    Span4Mux_h I__5949 (
            .O(N__32037),
            .I(N__31994));
    Sp12to4 I__5948 (
            .O(N__32034),
            .I(N__31987));
    Span12Mux_h I__5947 (
            .O(N__32031),
            .I(N__31987));
    Span12Mux_s5_h I__5946 (
            .O(N__32026),
            .I(N__31987));
    Span4Mux_h I__5945 (
            .O(N__32023),
            .I(N__31982));
    Span4Mux_v I__5944 (
            .O(N__32014),
            .I(N__31982));
    Span4Mux_v I__5943 (
            .O(N__32011),
            .I(N__31977));
    Span4Mux_v I__5942 (
            .O(N__32004),
            .I(N__31977));
    LocalMux I__5941 (
            .O(N__31997),
            .I(aZ0Z_1));
    Odrv4 I__5940 (
            .O(N__31994),
            .I(aZ0Z_1));
    Odrv12 I__5939 (
            .O(N__31987),
            .I(aZ0Z_1));
    Odrv4 I__5938 (
            .O(N__31982),
            .I(aZ0Z_1));
    Odrv4 I__5937 (
            .O(N__31977),
            .I(aZ0Z_1));
    CascadeMux I__5936 (
            .O(N__31966),
            .I(\ALU.un2_addsub_axb_4_cascade_ ));
    InMux I__5935 (
            .O(N__31963),
            .I(N__31960));
    LocalMux I__5934 (
            .O(N__31960),
            .I(N__31957));
    Odrv12 I__5933 (
            .O(N__31957),
            .I(\ALU.un9_addsub_axb_3 ));
    InMux I__5932 (
            .O(N__31954),
            .I(N__31951));
    LocalMux I__5931 (
            .O(N__31951),
            .I(N__31948));
    Span4Mux_v I__5930 (
            .O(N__31948),
            .I(N__31945));
    Span4Mux_h I__5929 (
            .O(N__31945),
            .I(N__31942));
    Span4Mux_h I__5928 (
            .O(N__31942),
            .I(N__31939));
    Odrv4 I__5927 (
            .O(N__31939),
            .I(\ALU.madd_490_5 ));
    InMux I__5926 (
            .O(N__31936),
            .I(N__31931));
    InMux I__5925 (
            .O(N__31935),
            .I(N__31928));
    InMux I__5924 (
            .O(N__31934),
            .I(N__31925));
    LocalMux I__5923 (
            .O(N__31931),
            .I(N__31918));
    LocalMux I__5922 (
            .O(N__31928),
            .I(N__31915));
    LocalMux I__5921 (
            .O(N__31925),
            .I(N__31912));
    InMux I__5920 (
            .O(N__31924),
            .I(N__31908));
    InMux I__5919 (
            .O(N__31923),
            .I(N__31903));
    InMux I__5918 (
            .O(N__31922),
            .I(N__31903));
    InMux I__5917 (
            .O(N__31921),
            .I(N__31898));
    Span4Mux_h I__5916 (
            .O(N__31918),
            .I(N__31893));
    Span4Mux_s1_v I__5915 (
            .O(N__31915),
            .I(N__31893));
    Span4Mux_v I__5914 (
            .O(N__31912),
            .I(N__31890));
    InMux I__5913 (
            .O(N__31911),
            .I(N__31887));
    LocalMux I__5912 (
            .O(N__31908),
            .I(N__31882));
    LocalMux I__5911 (
            .O(N__31903),
            .I(N__31882));
    InMux I__5910 (
            .O(N__31902),
            .I(N__31879));
    InMux I__5909 (
            .O(N__31901),
            .I(N__31876));
    LocalMux I__5908 (
            .O(N__31898),
            .I(N__31873));
    Span4Mux_v I__5907 (
            .O(N__31893),
            .I(N__31870));
    Span4Mux_h I__5906 (
            .O(N__31890),
            .I(N__31863));
    LocalMux I__5905 (
            .O(N__31887),
            .I(N__31863));
    Span4Mux_h I__5904 (
            .O(N__31882),
            .I(N__31863));
    LocalMux I__5903 (
            .O(N__31879),
            .I(N__31858));
    LocalMux I__5902 (
            .O(N__31876),
            .I(N__31858));
    Span4Mux_v I__5901 (
            .O(N__31873),
            .I(N__31853));
    Span4Mux_v I__5900 (
            .O(N__31870),
            .I(N__31853));
    Span4Mux_v I__5899 (
            .O(N__31863),
            .I(N__31850));
    Span4Mux_v I__5898 (
            .O(N__31858),
            .I(N__31847));
    Odrv4 I__5897 (
            .O(N__31853),
            .I(\ALU.r6_RNIFJ8D2Z0Z_3 ));
    Odrv4 I__5896 (
            .O(N__31850),
            .I(\ALU.r6_RNIFJ8D2Z0Z_3 ));
    Odrv4 I__5895 (
            .O(N__31847),
            .I(\ALU.r6_RNIFJ8D2Z0Z_3 ));
    CascadeMux I__5894 (
            .O(N__31840),
            .I(N__31836));
    InMux I__5893 (
            .O(N__31839),
            .I(N__31830));
    InMux I__5892 (
            .O(N__31836),
            .I(N__31825));
    InMux I__5891 (
            .O(N__31835),
            .I(N__31819));
    InMux I__5890 (
            .O(N__31834),
            .I(N__31819));
    CascadeMux I__5889 (
            .O(N__31833),
            .I(N__31816));
    LocalMux I__5888 (
            .O(N__31830),
            .I(N__31813));
    InMux I__5887 (
            .O(N__31829),
            .I(N__31810));
    InMux I__5886 (
            .O(N__31828),
            .I(N__31807));
    LocalMux I__5885 (
            .O(N__31825),
            .I(N__31804));
    InMux I__5884 (
            .O(N__31824),
            .I(N__31801));
    LocalMux I__5883 (
            .O(N__31819),
            .I(N__31798));
    InMux I__5882 (
            .O(N__31816),
            .I(N__31793));
    Span4Mux_v I__5881 (
            .O(N__31813),
            .I(N__31788));
    LocalMux I__5880 (
            .O(N__31810),
            .I(N__31788));
    LocalMux I__5879 (
            .O(N__31807),
            .I(N__31785));
    Span4Mux_s3_v I__5878 (
            .O(N__31804),
            .I(N__31782));
    LocalMux I__5877 (
            .O(N__31801),
            .I(N__31779));
    Span4Mux_v I__5876 (
            .O(N__31798),
            .I(N__31776));
    InMux I__5875 (
            .O(N__31797),
            .I(N__31771));
    InMux I__5874 (
            .O(N__31796),
            .I(N__31771));
    LocalMux I__5873 (
            .O(N__31793),
            .I(N__31768));
    Span4Mux_h I__5872 (
            .O(N__31788),
            .I(N__31765));
    Span4Mux_s3_v I__5871 (
            .O(N__31785),
            .I(N__31760));
    Span4Mux_h I__5870 (
            .O(N__31782),
            .I(N__31760));
    Span4Mux_v I__5869 (
            .O(N__31779),
            .I(N__31755));
    Span4Mux_h I__5868 (
            .O(N__31776),
            .I(N__31755));
    LocalMux I__5867 (
            .O(N__31771),
            .I(N__31752));
    Odrv12 I__5866 (
            .O(N__31768),
            .I(\ALU.r4_RNIMQ992Z0Z_3 ));
    Odrv4 I__5865 (
            .O(N__31765),
            .I(\ALU.r4_RNIMQ992Z0Z_3 ));
    Odrv4 I__5864 (
            .O(N__31760),
            .I(\ALU.r4_RNIMQ992Z0Z_3 ));
    Odrv4 I__5863 (
            .O(N__31755),
            .I(\ALU.r4_RNIMQ992Z0Z_3 ));
    Odrv12 I__5862 (
            .O(N__31752),
            .I(\ALU.r4_RNIMQ992Z0Z_3 ));
    InMux I__5861 (
            .O(N__31741),
            .I(N__31735));
    CascadeMux I__5860 (
            .O(N__31740),
            .I(N__31732));
    InMux I__5859 (
            .O(N__31739),
            .I(N__31726));
    InMux I__5858 (
            .O(N__31738),
            .I(N__31726));
    LocalMux I__5857 (
            .O(N__31735),
            .I(N__31723));
    InMux I__5856 (
            .O(N__31732),
            .I(N__31714));
    InMux I__5855 (
            .O(N__31731),
            .I(N__31714));
    LocalMux I__5854 (
            .O(N__31726),
            .I(N__31711));
    Span4Mux_v I__5853 (
            .O(N__31723),
            .I(N__31708));
    InMux I__5852 (
            .O(N__31722),
            .I(N__31701));
    InMux I__5851 (
            .O(N__31721),
            .I(N__31701));
    InMux I__5850 (
            .O(N__31720),
            .I(N__31701));
    InMux I__5849 (
            .O(N__31719),
            .I(N__31698));
    LocalMux I__5848 (
            .O(N__31714),
            .I(N__31695));
    Span4Mux_s3_v I__5847 (
            .O(N__31711),
            .I(N__31692));
    Span4Mux_h I__5846 (
            .O(N__31708),
            .I(N__31687));
    LocalMux I__5845 (
            .O(N__31701),
            .I(N__31687));
    LocalMux I__5844 (
            .O(N__31698),
            .I(N__31684));
    Span4Mux_s3_v I__5843 (
            .O(N__31695),
            .I(N__31681));
    Span4Mux_v I__5842 (
            .O(N__31692),
            .I(N__31678));
    Span4Mux_h I__5841 (
            .O(N__31687),
            .I(N__31675));
    Odrv12 I__5840 (
            .O(N__31684),
            .I(\ALU.r4_RNIDI992Z0Z_1 ));
    Odrv4 I__5839 (
            .O(N__31681),
            .I(\ALU.r4_RNIDI992Z0Z_1 ));
    Odrv4 I__5838 (
            .O(N__31678),
            .I(\ALU.r4_RNIDI992Z0Z_1 ));
    Odrv4 I__5837 (
            .O(N__31675),
            .I(\ALU.r4_RNIDI992Z0Z_1 ));
    InMux I__5836 (
            .O(N__31666),
            .I(N__31661));
    InMux I__5835 (
            .O(N__31665),
            .I(N__31656));
    InMux I__5834 (
            .O(N__31664),
            .I(N__31656));
    LocalMux I__5833 (
            .O(N__31661),
            .I(N__31652));
    LocalMux I__5832 (
            .O(N__31656),
            .I(N__31649));
    InMux I__5831 (
            .O(N__31655),
            .I(N__31644));
    Span4Mux_s1_v I__5830 (
            .O(N__31652),
            .I(N__31641));
    Span4Mux_s1_v I__5829 (
            .O(N__31649),
            .I(N__31638));
    InMux I__5828 (
            .O(N__31648),
            .I(N__31633));
    InMux I__5827 (
            .O(N__31647),
            .I(N__31633));
    LocalMux I__5826 (
            .O(N__31644),
            .I(N__31627));
    Span4Mux_v I__5825 (
            .O(N__31641),
            .I(N__31622));
    Span4Mux_v I__5824 (
            .O(N__31638),
            .I(N__31622));
    LocalMux I__5823 (
            .O(N__31633),
            .I(N__31619));
    InMux I__5822 (
            .O(N__31632),
            .I(N__31612));
    InMux I__5821 (
            .O(N__31631),
            .I(N__31612));
    InMux I__5820 (
            .O(N__31630),
            .I(N__31612));
    Span4Mux_h I__5819 (
            .O(N__31627),
            .I(N__31609));
    Span4Mux_h I__5818 (
            .O(N__31622),
            .I(N__31606));
    Span12Mux_s8_v I__5817 (
            .O(N__31619),
            .I(N__31603));
    LocalMux I__5816 (
            .O(N__31612),
            .I(N__31600));
    Odrv4 I__5815 (
            .O(N__31609),
            .I(\ALU.r6_RNI7B8D2Z0Z_1 ));
    Odrv4 I__5814 (
            .O(N__31606),
            .I(\ALU.r6_RNI7B8D2Z0Z_1 ));
    Odrv12 I__5813 (
            .O(N__31603),
            .I(\ALU.r6_RNI7B8D2Z0Z_1 ));
    Odrv12 I__5812 (
            .O(N__31600),
            .I(\ALU.r6_RNI7B8D2Z0Z_1 ));
    InMux I__5811 (
            .O(N__31591),
            .I(N__31582));
    InMux I__5810 (
            .O(N__31590),
            .I(N__31582));
    InMux I__5809 (
            .O(N__31589),
            .I(N__31582));
    LocalMux I__5808 (
            .O(N__31582),
            .I(N__31579));
    Odrv4 I__5807 (
            .O(N__31579),
            .I(\ALU.a1_b_3 ));
    CascadeMux I__5806 (
            .O(N__31576),
            .I(N__31572));
    CascadeMux I__5805 (
            .O(N__31575),
            .I(N__31569));
    InMux I__5804 (
            .O(N__31572),
            .I(N__31564));
    InMux I__5803 (
            .O(N__31569),
            .I(N__31564));
    LocalMux I__5802 (
            .O(N__31564),
            .I(N__31560));
    InMux I__5801 (
            .O(N__31563),
            .I(N__31557));
    Span4Mux_s1_v I__5800 (
            .O(N__31560),
            .I(N__31554));
    LocalMux I__5799 (
            .O(N__31557),
            .I(N__31551));
    Span4Mux_s2_h I__5798 (
            .O(N__31554),
            .I(N__31548));
    Span4Mux_h I__5797 (
            .O(N__31551),
            .I(N__31543));
    Span4Mux_h I__5796 (
            .O(N__31548),
            .I(N__31543));
    Odrv4 I__5795 (
            .O(N__31543),
            .I(\ALU.madd_135_0 ));
    InMux I__5794 (
            .O(N__31540),
            .I(N__31537));
    LocalMux I__5793 (
            .O(N__31537),
            .I(N__31534));
    Odrv4 I__5792 (
            .O(N__31534),
            .I(\ALU.lshift_3_ns_1_6 ));
    InMux I__5791 (
            .O(N__31531),
            .I(N__31528));
    LocalMux I__5790 (
            .O(N__31528),
            .I(N__31525));
    Span4Mux_s3_v I__5789 (
            .O(N__31525),
            .I(N__31522));
    Span4Mux_h I__5788 (
            .O(N__31522),
            .I(N__31519));
    Odrv4 I__5787 (
            .O(N__31519),
            .I(\ALU.lshift_3_ns_1_7 ));
    InMux I__5786 (
            .O(N__31516),
            .I(\ALU.r0_12_s1_13 ));
    InMux I__5785 (
            .O(N__31513),
            .I(N__31510));
    LocalMux I__5784 (
            .O(N__31510),
            .I(N__31507));
    Odrv12 I__5783 (
            .O(N__31507),
            .I(\ALU.r0_12_s1_13_THRU_CO ));
    CascadeMux I__5782 (
            .O(N__31504),
            .I(N__31501));
    InMux I__5781 (
            .O(N__31501),
            .I(N__31498));
    LocalMux I__5780 (
            .O(N__31498),
            .I(\ALU.r0_12_prm_1_13_s1_c_RNOZ0 ));
    CascadeMux I__5779 (
            .O(N__31495),
            .I(\ALU.rshift_3_ns_1_2_cascade_ ));
    InMux I__5778 (
            .O(N__31492),
            .I(N__31489));
    LocalMux I__5777 (
            .O(N__31489),
            .I(N__31486));
    Span4Mux_h I__5776 (
            .O(N__31486),
            .I(N__31483));
    Span4Mux_h I__5775 (
            .O(N__31483),
            .I(N__31480));
    Odrv4 I__5774 (
            .O(N__31480),
            .I(\ALU.r0_12_prm_7_13_s1_c_RNOZ0 ));
    CascadeMux I__5773 (
            .O(N__31477),
            .I(N__31473));
    InMux I__5772 (
            .O(N__31476),
            .I(N__31470));
    InMux I__5771 (
            .O(N__31473),
            .I(N__31467));
    LocalMux I__5770 (
            .O(N__31470),
            .I(N__31464));
    LocalMux I__5769 (
            .O(N__31467),
            .I(N__31461));
    Span4Mux_v I__5768 (
            .O(N__31464),
            .I(N__31458));
    Span4Mux_v I__5767 (
            .O(N__31461),
            .I(N__31455));
    Span4Mux_h I__5766 (
            .O(N__31458),
            .I(N__31452));
    Sp12to4 I__5765 (
            .O(N__31455),
            .I(N__31449));
    Odrv4 I__5764 (
            .O(N__31452),
            .I(\ALU.r5_RNID2JJ9_0Z0Z_13 ));
    Odrv12 I__5763 (
            .O(N__31449),
            .I(\ALU.r5_RNID2JJ9_0Z0Z_13 ));
    InMux I__5762 (
            .O(N__31444),
            .I(N__31441));
    LocalMux I__5761 (
            .O(N__31441),
            .I(N__31438));
    Span4Mux_h I__5760 (
            .O(N__31438),
            .I(N__31435));
    Odrv4 I__5759 (
            .O(N__31435),
            .I(\ALU.r0_12_prm_6_13_s1_c_RNOZ0 ));
    InMux I__5758 (
            .O(N__31432),
            .I(N__31429));
    LocalMux I__5757 (
            .O(N__31429),
            .I(N__31425));
    CascadeMux I__5756 (
            .O(N__31428),
            .I(N__31422));
    Span4Mux_h I__5755 (
            .O(N__31425),
            .I(N__31419));
    InMux I__5754 (
            .O(N__31422),
            .I(N__31416));
    Odrv4 I__5753 (
            .O(N__31419),
            .I(\ALU.un14_log_0_i_13 ));
    LocalMux I__5752 (
            .O(N__31416),
            .I(\ALU.un14_log_0_i_13 ));
    InMux I__5751 (
            .O(N__31411),
            .I(N__31408));
    LocalMux I__5750 (
            .O(N__31408),
            .I(N__31405));
    Span4Mux_h I__5749 (
            .O(N__31405),
            .I(N__31402));
    Odrv4 I__5748 (
            .O(N__31402),
            .I(\ALU.r0_12_prm_5_13_s1_c_RNOZ0 ));
    CascadeMux I__5747 (
            .O(N__31399),
            .I(N__31395));
    CascadeMux I__5746 (
            .O(N__31398),
            .I(N__31392));
    InMux I__5745 (
            .O(N__31395),
            .I(N__31389));
    InMux I__5744 (
            .O(N__31392),
            .I(N__31386));
    LocalMux I__5743 (
            .O(N__31389),
            .I(N__31383));
    LocalMux I__5742 (
            .O(N__31386),
            .I(N__31378));
    Span4Mux_h I__5741 (
            .O(N__31383),
            .I(N__31378));
    Span4Mux_h I__5740 (
            .O(N__31378),
            .I(N__31375));
    Odrv4 I__5739 (
            .O(N__31375),
            .I(\ALU.r5_RNID2JJ9_1Z0Z_13 ));
    InMux I__5738 (
            .O(N__31372),
            .I(N__31369));
    LocalMux I__5737 (
            .O(N__31369),
            .I(N__31366));
    Span4Mux_h I__5736 (
            .O(N__31366),
            .I(N__31363));
    Odrv4 I__5735 (
            .O(N__31363),
            .I(\ALU.r0_12_prm_4_13_s1_c_RNOZ0 ));
    CascadeMux I__5734 (
            .O(N__31360),
            .I(N__31356));
    InMux I__5733 (
            .O(N__31359),
            .I(N__31353));
    InMux I__5732 (
            .O(N__31356),
            .I(N__31350));
    LocalMux I__5731 (
            .O(N__31353),
            .I(N__31345));
    LocalMux I__5730 (
            .O(N__31350),
            .I(N__31345));
    Odrv4 I__5729 (
            .O(N__31345),
            .I(\ALU.a_i_13 ));
    InMux I__5728 (
            .O(N__31342),
            .I(N__31339));
    LocalMux I__5727 (
            .O(N__31339),
            .I(\ALU.rshift_10_ns_1_3 ));
    CascadeMux I__5726 (
            .O(N__31336),
            .I(\ALU.r5_RNI465TIZ0Z_13_cascade_ ));
    InMux I__5725 (
            .O(N__31333),
            .I(N__31330));
    LocalMux I__5724 (
            .O(N__31330),
            .I(N__31327));
    Span4Mux_v I__5723 (
            .O(N__31327),
            .I(N__31324));
    Span4Mux_v I__5722 (
            .O(N__31324),
            .I(N__31321));
    Odrv4 I__5721 (
            .O(N__31321),
            .I(\ALU.r5_RNIOL1S71Z0Z_10 ));
    CascadeMux I__5720 (
            .O(N__31318),
            .I(N__31315));
    InMux I__5719 (
            .O(N__31315),
            .I(N__31312));
    LocalMux I__5718 (
            .O(N__31312),
            .I(N__31309));
    Span4Mux_h I__5717 (
            .O(N__31309),
            .I(N__31306));
    Odrv4 I__5716 (
            .O(N__31306),
            .I(\ALU.r0_12_prm_5_12_s0_c_RNOZ0 ));
    CascadeMux I__5715 (
            .O(N__31303),
            .I(N__31300));
    InMux I__5714 (
            .O(N__31300),
            .I(N__31297));
    LocalMux I__5713 (
            .O(N__31297),
            .I(N__31294));
    Span4Mux_v I__5712 (
            .O(N__31294),
            .I(N__31291));
    Span4Mux_h I__5711 (
            .O(N__31291),
            .I(N__31288));
    Odrv4 I__5710 (
            .O(N__31288),
            .I(\ALU.r0_12_prm_8_11_s0_c_RNOZ0 ));
    CascadeMux I__5709 (
            .O(N__31285),
            .I(N__31282));
    InMux I__5708 (
            .O(N__31282),
            .I(N__31279));
    LocalMux I__5707 (
            .O(N__31279),
            .I(N__31276));
    Span4Mux_h I__5706 (
            .O(N__31276),
            .I(N__31273));
    Odrv4 I__5705 (
            .O(N__31273),
            .I(\ALU.r0_12_prm_7_12_s0_c_RNOZ0 ));
    CascadeMux I__5704 (
            .O(N__31270),
            .I(N__31267));
    InMux I__5703 (
            .O(N__31267),
            .I(N__31264));
    LocalMux I__5702 (
            .O(N__31264),
            .I(N__31261));
    Span4Mux_v I__5701 (
            .O(N__31261),
            .I(N__31258));
    Span4Mux_h I__5700 (
            .O(N__31258),
            .I(N__31255));
    Sp12to4 I__5699 (
            .O(N__31255),
            .I(N__31252));
    Odrv12 I__5698 (
            .O(N__31252),
            .I(\ALU.r0_12_prm_6_12_s0_c_RNOZ0 ));
    CascadeMux I__5697 (
            .O(N__31249),
            .I(N__31246));
    InMux I__5696 (
            .O(N__31246),
            .I(N__31243));
    LocalMux I__5695 (
            .O(N__31243),
            .I(N__31240));
    Span4Mux_h I__5694 (
            .O(N__31240),
            .I(N__31237));
    Odrv4 I__5693 (
            .O(N__31237),
            .I(\ALU.r0_12_prm_2_15_s1_c_RNOZ0 ));
    CascadeMux I__5692 (
            .O(N__31234),
            .I(N__31231));
    InMux I__5691 (
            .O(N__31231),
            .I(N__31228));
    LocalMux I__5690 (
            .O(N__31228),
            .I(N__31225));
    Span4Mux_v I__5689 (
            .O(N__31225),
            .I(N__31222));
    Span4Mux_h I__5688 (
            .O(N__31222),
            .I(N__31219));
    Odrv4 I__5687 (
            .O(N__31219),
            .I(\ALU.r0_12_prm_2_13_s0_c_RNOZ0 ));
    CascadeMux I__5686 (
            .O(N__31216),
            .I(N__31213));
    InMux I__5685 (
            .O(N__31213),
            .I(N__31210));
    LocalMux I__5684 (
            .O(N__31210),
            .I(N__31207));
    Span4Mux_h I__5683 (
            .O(N__31207),
            .I(N__31204));
    Odrv4 I__5682 (
            .O(N__31204),
            .I(\ALU.r0_12_prm_1_14_s0_c_RNOZ0 ));
    CascadeMux I__5681 (
            .O(N__31201),
            .I(N__31198));
    InMux I__5680 (
            .O(N__31198),
            .I(N__31195));
    LocalMux I__5679 (
            .O(N__31195),
            .I(N__31192));
    Span4Mux_h I__5678 (
            .O(N__31192),
            .I(N__31189));
    Odrv4 I__5677 (
            .O(N__31189),
            .I(\ALU.r0_12_prm_8_15_s1_c_RNOZ0 ));
    InMux I__5676 (
            .O(N__31186),
            .I(N__31183));
    LocalMux I__5675 (
            .O(N__31183),
            .I(\ALU.r0_12_prm_3_9_s0_sf ));
    CascadeMux I__5674 (
            .O(N__31180),
            .I(N__31177));
    InMux I__5673 (
            .O(N__31177),
            .I(N__31174));
    LocalMux I__5672 (
            .O(N__31174),
            .I(N__31171));
    Span4Mux_h I__5671 (
            .O(N__31171),
            .I(N__31168));
    Span4Mux_h I__5670 (
            .O(N__31168),
            .I(N__31165));
    Odrv4 I__5669 (
            .O(N__31165),
            .I(\ALU.r0_12_prm_2_9_s0_c_RNOZ0 ));
    InMux I__5668 (
            .O(N__31162),
            .I(N__31159));
    LocalMux I__5667 (
            .O(N__31159),
            .I(N__31156));
    Span4Mux_v I__5666 (
            .O(N__31156),
            .I(N__31153));
    Odrv4 I__5665 (
            .O(N__31153),
            .I(\ALU.mult_9 ));
    InMux I__5664 (
            .O(N__31150),
            .I(\ALU.r0_12_s0_9 ));
    InMux I__5663 (
            .O(N__31147),
            .I(N__31143));
    InMux I__5662 (
            .O(N__31146),
            .I(N__31140));
    LocalMux I__5661 (
            .O(N__31143),
            .I(N__31135));
    LocalMux I__5660 (
            .O(N__31140),
            .I(N__31135));
    Span4Mux_h I__5659 (
            .O(N__31135),
            .I(N__31131));
    InMux I__5658 (
            .O(N__31134),
            .I(N__31128));
    Span4Mux_h I__5657 (
            .O(N__31131),
            .I(N__31123));
    LocalMux I__5656 (
            .O(N__31128),
            .I(N__31123));
    Odrv4 I__5655 (
            .O(N__31123),
            .I(r0_9));
    CascadeMux I__5654 (
            .O(N__31120),
            .I(N__31117));
    InMux I__5653 (
            .O(N__31117),
            .I(N__31114));
    LocalMux I__5652 (
            .O(N__31114),
            .I(N__31111));
    Span4Mux_v I__5651 (
            .O(N__31111),
            .I(N__31108));
    Span4Mux_h I__5650 (
            .O(N__31108),
            .I(N__31105));
    Span4Mux_v I__5649 (
            .O(N__31105),
            .I(N__31102));
    Odrv4 I__5648 (
            .O(N__31102),
            .I(\ALU.r0_12_prm_8_11_s1_c_RNOZ0 ));
    CascadeMux I__5647 (
            .O(N__31099),
            .I(\ALU.a_3_ns_1_4_cascade_ ));
    InMux I__5646 (
            .O(N__31096),
            .I(N__31092));
    CascadeMux I__5645 (
            .O(N__31095),
            .I(N__31089));
    LocalMux I__5644 (
            .O(N__31092),
            .I(N__31081));
    InMux I__5643 (
            .O(N__31089),
            .I(N__31072));
    InMux I__5642 (
            .O(N__31088),
            .I(N__31072));
    InMux I__5641 (
            .O(N__31087),
            .I(N__31072));
    InMux I__5640 (
            .O(N__31086),
            .I(N__31072));
    CascadeMux I__5639 (
            .O(N__31085),
            .I(N__31069));
    CascadeMux I__5638 (
            .O(N__31084),
            .I(N__31063));
    Span4Mux_s1_h I__5637 (
            .O(N__31081),
            .I(N__31057));
    LocalMux I__5636 (
            .O(N__31072),
            .I(N__31054));
    InMux I__5635 (
            .O(N__31069),
            .I(N__31047));
    InMux I__5634 (
            .O(N__31068),
            .I(N__31047));
    InMux I__5633 (
            .O(N__31067),
            .I(N__31047));
    InMux I__5632 (
            .O(N__31066),
            .I(N__31044));
    InMux I__5631 (
            .O(N__31063),
            .I(N__31041));
    InMux I__5630 (
            .O(N__31062),
            .I(N__31038));
    InMux I__5629 (
            .O(N__31061),
            .I(N__31033));
    InMux I__5628 (
            .O(N__31060),
            .I(N__31033));
    Span4Mux_h I__5627 (
            .O(N__31057),
            .I(N__31028));
    Span4Mux_h I__5626 (
            .O(N__31054),
            .I(N__31028));
    LocalMux I__5625 (
            .O(N__31047),
            .I(N__31025));
    LocalMux I__5624 (
            .O(N__31044),
            .I(a_fastZ0Z_2));
    LocalMux I__5623 (
            .O(N__31041),
            .I(a_fastZ0Z_2));
    LocalMux I__5622 (
            .O(N__31038),
            .I(a_fastZ0Z_2));
    LocalMux I__5621 (
            .O(N__31033),
            .I(a_fastZ0Z_2));
    Odrv4 I__5620 (
            .O(N__31028),
            .I(a_fastZ0Z_2));
    Odrv4 I__5619 (
            .O(N__31025),
            .I(a_fastZ0Z_2));
    CascadeMux I__5618 (
            .O(N__31012),
            .I(N__31007));
    InMux I__5617 (
            .O(N__31011),
            .I(N__31004));
    InMux I__5616 (
            .O(N__31010),
            .I(N__31001));
    InMux I__5615 (
            .O(N__31007),
            .I(N__30998));
    LocalMux I__5614 (
            .O(N__31004),
            .I(N__30995));
    LocalMux I__5613 (
            .O(N__31001),
            .I(N__30990));
    LocalMux I__5612 (
            .O(N__30998),
            .I(N__30990));
    Span4Mux_h I__5611 (
            .O(N__30995),
            .I(N__30987));
    Span4Mux_h I__5610 (
            .O(N__30990),
            .I(N__30984));
    Odrv4 I__5609 (
            .O(N__30987),
            .I(r1_9));
    Odrv4 I__5608 (
            .O(N__30984),
            .I(r1_9));
    InMux I__5607 (
            .O(N__30979),
            .I(N__30965));
    InMux I__5606 (
            .O(N__30978),
            .I(N__30965));
    InMux I__5605 (
            .O(N__30977),
            .I(N__30958));
    InMux I__5604 (
            .O(N__30976),
            .I(N__30958));
    InMux I__5603 (
            .O(N__30975),
            .I(N__30958));
    InMux I__5602 (
            .O(N__30974),
            .I(N__30947));
    InMux I__5601 (
            .O(N__30973),
            .I(N__30947));
    InMux I__5600 (
            .O(N__30972),
            .I(N__30947));
    InMux I__5599 (
            .O(N__30971),
            .I(N__30947));
    InMux I__5598 (
            .O(N__30970),
            .I(N__30947));
    LocalMux I__5597 (
            .O(N__30965),
            .I(N__30944));
    LocalMux I__5596 (
            .O(N__30958),
            .I(a_fastZ0Z_0));
    LocalMux I__5595 (
            .O(N__30947),
            .I(a_fastZ0Z_0));
    Odrv4 I__5594 (
            .O(N__30944),
            .I(a_fastZ0Z_0));
    InMux I__5593 (
            .O(N__30937),
            .I(N__30931));
    InMux I__5592 (
            .O(N__30936),
            .I(N__30931));
    LocalMux I__5591 (
            .O(N__30931),
            .I(N__30921));
    InMux I__5590 (
            .O(N__30930),
            .I(N__30916));
    InMux I__5589 (
            .O(N__30929),
            .I(N__30916));
    InMux I__5588 (
            .O(N__30928),
            .I(N__30909));
    InMux I__5587 (
            .O(N__30927),
            .I(N__30906));
    InMux I__5586 (
            .O(N__30926),
            .I(N__30903));
    InMux I__5585 (
            .O(N__30925),
            .I(N__30900));
    InMux I__5584 (
            .O(N__30924),
            .I(N__30897));
    Span4Mux_v I__5583 (
            .O(N__30921),
            .I(N__30894));
    LocalMux I__5582 (
            .O(N__30916),
            .I(N__30891));
    InMux I__5581 (
            .O(N__30915),
            .I(N__30880));
    InMux I__5580 (
            .O(N__30914),
            .I(N__30880));
    InMux I__5579 (
            .O(N__30913),
            .I(N__30875));
    InMux I__5578 (
            .O(N__30912),
            .I(N__30875));
    LocalMux I__5577 (
            .O(N__30909),
            .I(N__30872));
    LocalMux I__5576 (
            .O(N__30906),
            .I(N__30867));
    LocalMux I__5575 (
            .O(N__30903),
            .I(N__30867));
    LocalMux I__5574 (
            .O(N__30900),
            .I(N__30862));
    LocalMux I__5573 (
            .O(N__30897),
            .I(N__30862));
    Span4Mux_v I__5572 (
            .O(N__30894),
            .I(N__30857));
    Span4Mux_v I__5571 (
            .O(N__30891),
            .I(N__30857));
    InMux I__5570 (
            .O(N__30890),
            .I(N__30852));
    InMux I__5569 (
            .O(N__30889),
            .I(N__30852));
    InMux I__5568 (
            .O(N__30888),
            .I(N__30845));
    InMux I__5567 (
            .O(N__30887),
            .I(N__30845));
    InMux I__5566 (
            .O(N__30886),
            .I(N__30845));
    InMux I__5565 (
            .O(N__30885),
            .I(N__30842));
    LocalMux I__5564 (
            .O(N__30880),
            .I(N__30833));
    LocalMux I__5563 (
            .O(N__30875),
            .I(N__30833));
    Span4Mux_h I__5562 (
            .O(N__30872),
            .I(N__30833));
    Span4Mux_h I__5561 (
            .O(N__30867),
            .I(N__30833));
    Span4Mux_v I__5560 (
            .O(N__30862),
            .I(N__30828));
    Span4Mux_h I__5559 (
            .O(N__30857),
            .I(N__30828));
    LocalMux I__5558 (
            .O(N__30852),
            .I(a_2_repZ0Z2));
    LocalMux I__5557 (
            .O(N__30845),
            .I(a_2_repZ0Z2));
    LocalMux I__5556 (
            .O(N__30842),
            .I(a_2_repZ0Z2));
    Odrv4 I__5555 (
            .O(N__30833),
            .I(a_2_repZ0Z2));
    Odrv4 I__5554 (
            .O(N__30828),
            .I(a_2_repZ0Z2));
    CascadeMux I__5553 (
            .O(N__30817),
            .I(\ALU.a_3_ns_1_9_cascade_ ));
    InMux I__5552 (
            .O(N__30814),
            .I(N__30808));
    InMux I__5551 (
            .O(N__30813),
            .I(N__30805));
    InMux I__5550 (
            .O(N__30812),
            .I(N__30802));
    InMux I__5549 (
            .O(N__30811),
            .I(N__30799));
    LocalMux I__5548 (
            .O(N__30808),
            .I(N__30796));
    LocalMux I__5547 (
            .O(N__30805),
            .I(N__30791));
    LocalMux I__5546 (
            .O(N__30802),
            .I(N__30791));
    LocalMux I__5545 (
            .O(N__30799),
            .I(N__30788));
    Span4Mux_v I__5544 (
            .O(N__30796),
            .I(N__30785));
    Span4Mux_h I__5543 (
            .O(N__30791),
            .I(N__30782));
    Span4Mux_h I__5542 (
            .O(N__30788),
            .I(N__30779));
    Span4Mux_h I__5541 (
            .O(N__30785),
            .I(N__30774));
    Span4Mux_v I__5540 (
            .O(N__30782),
            .I(N__30774));
    Odrv4 I__5539 (
            .O(N__30779),
            .I(\ALU.r4_RNIEJA92Z0Z_9 ));
    Odrv4 I__5538 (
            .O(N__30774),
            .I(\ALU.r4_RNIEJA92Z0Z_9 ));
    CascadeMux I__5537 (
            .O(N__30769),
            .I(N__30766));
    InMux I__5536 (
            .O(N__30766),
            .I(N__30763));
    LocalMux I__5535 (
            .O(N__30763),
            .I(N__30760));
    Span4Mux_h I__5534 (
            .O(N__30760),
            .I(N__30757));
    Span4Mux_v I__5533 (
            .O(N__30757),
            .I(N__30754));
    Odrv4 I__5532 (
            .O(N__30754),
            .I(\ALU.r0_12_prm_6_9_s0_c_RNOZ0 ));
    InMux I__5531 (
            .O(N__30751),
            .I(N__30748));
    LocalMux I__5530 (
            .O(N__30748),
            .I(N__30745));
    Span4Mux_v I__5529 (
            .O(N__30745),
            .I(N__30742));
    Span4Mux_h I__5528 (
            .O(N__30742),
            .I(N__30737));
    InMux I__5527 (
            .O(N__30741),
            .I(N__30732));
    InMux I__5526 (
            .O(N__30740),
            .I(N__30732));
    Odrv4 I__5525 (
            .O(N__30737),
            .I(r0_7));
    LocalMux I__5524 (
            .O(N__30732),
            .I(r0_7));
    CascadeMux I__5523 (
            .O(N__30727),
            .I(\ALU.a_3_ns_1_7_cascade_ ));
    InMux I__5522 (
            .O(N__30724),
            .I(N__30719));
    InMux I__5521 (
            .O(N__30723),
            .I(N__30716));
    InMux I__5520 (
            .O(N__30722),
            .I(N__30712));
    LocalMux I__5519 (
            .O(N__30719),
            .I(N__30708));
    LocalMux I__5518 (
            .O(N__30716),
            .I(N__30705));
    InMux I__5517 (
            .O(N__30715),
            .I(N__30702));
    LocalMux I__5516 (
            .O(N__30712),
            .I(N__30699));
    InMux I__5515 (
            .O(N__30711),
            .I(N__30696));
    Span4Mux_h I__5514 (
            .O(N__30708),
            .I(N__30693));
    Span4Mux_h I__5513 (
            .O(N__30705),
            .I(N__30688));
    LocalMux I__5512 (
            .O(N__30702),
            .I(N__30688));
    Span4Mux_v I__5511 (
            .O(N__30699),
            .I(N__30685));
    LocalMux I__5510 (
            .O(N__30696),
            .I(N__30682));
    Span4Mux_h I__5509 (
            .O(N__30693),
            .I(N__30679));
    Span4Mux_h I__5508 (
            .O(N__30688),
            .I(N__30676));
    Span4Mux_h I__5507 (
            .O(N__30685),
            .I(N__30671));
    Span4Mux_v I__5506 (
            .O(N__30682),
            .I(N__30671));
    Odrv4 I__5505 (
            .O(N__30679),
            .I(\ALU.r4_RNI6BA92Z0Z_7 ));
    Odrv4 I__5504 (
            .O(N__30676),
            .I(\ALU.r4_RNI6BA92Z0Z_7 ));
    Odrv4 I__5503 (
            .O(N__30671),
            .I(\ALU.r4_RNI6BA92Z0Z_7 ));
    CascadeMux I__5502 (
            .O(N__30664),
            .I(N__30660));
    CascadeMux I__5501 (
            .O(N__30663),
            .I(N__30657));
    InMux I__5500 (
            .O(N__30660),
            .I(N__30653));
    InMux I__5499 (
            .O(N__30657),
            .I(N__30650));
    InMux I__5498 (
            .O(N__30656),
            .I(N__30647));
    LocalMux I__5497 (
            .O(N__30653),
            .I(N__30644));
    LocalMux I__5496 (
            .O(N__30650),
            .I(N__30641));
    LocalMux I__5495 (
            .O(N__30647),
            .I(N__30638));
    Span12Mux_s10_v I__5494 (
            .O(N__30644),
            .I(N__30635));
    Span4Mux_h I__5493 (
            .O(N__30641),
            .I(N__30632));
    Odrv4 I__5492 (
            .O(N__30638),
            .I(r1_8));
    Odrv12 I__5491 (
            .O(N__30635),
            .I(r1_8));
    Odrv4 I__5490 (
            .O(N__30632),
            .I(r1_8));
    CascadeMux I__5489 (
            .O(N__30625),
            .I(\ALU.a_3_ns_1_8_cascade_ ));
    InMux I__5488 (
            .O(N__30622),
            .I(N__30618));
    CascadeMux I__5487 (
            .O(N__30621),
            .I(N__30615));
    LocalMux I__5486 (
            .O(N__30618),
            .I(N__30610));
    InMux I__5485 (
            .O(N__30615),
            .I(N__30605));
    InMux I__5484 (
            .O(N__30614),
            .I(N__30605));
    InMux I__5483 (
            .O(N__30613),
            .I(N__30602));
    Span4Mux_v I__5482 (
            .O(N__30610),
            .I(N__30599));
    LocalMux I__5481 (
            .O(N__30605),
            .I(N__30594));
    LocalMux I__5480 (
            .O(N__30602),
            .I(N__30594));
    Span4Mux_h I__5479 (
            .O(N__30599),
            .I(N__30591));
    Span4Mux_h I__5478 (
            .O(N__30594),
            .I(N__30588));
    Odrv4 I__5477 (
            .O(N__30591),
            .I(\ALU.r4_RNIAFA92Z0Z_8 ));
    Odrv4 I__5476 (
            .O(N__30588),
            .I(\ALU.r4_RNIAFA92Z0Z_8 ));
    InMux I__5475 (
            .O(N__30583),
            .I(N__30580));
    LocalMux I__5474 (
            .O(N__30580),
            .I(N__30577));
    Odrv4 I__5473 (
            .O(N__30577),
            .I(\ALU.a_3_ns_1_3 ));
    CascadeMux I__5472 (
            .O(N__30574),
            .I(\ALU.a_3_ns_1_2_cascade_ ));
    InMux I__5471 (
            .O(N__30571),
            .I(N__30564));
    InMux I__5470 (
            .O(N__30570),
            .I(N__30560));
    InMux I__5469 (
            .O(N__30569),
            .I(N__30554));
    InMux I__5468 (
            .O(N__30568),
            .I(N__30550));
    InMux I__5467 (
            .O(N__30567),
            .I(N__30547));
    LocalMux I__5466 (
            .O(N__30564),
            .I(N__30544));
    CascadeMux I__5465 (
            .O(N__30563),
            .I(N__30538));
    LocalMux I__5464 (
            .O(N__30560),
            .I(N__30535));
    InMux I__5463 (
            .O(N__30559),
            .I(N__30528));
    InMux I__5462 (
            .O(N__30558),
            .I(N__30528));
    InMux I__5461 (
            .O(N__30557),
            .I(N__30528));
    LocalMux I__5460 (
            .O(N__30554),
            .I(N__30525));
    InMux I__5459 (
            .O(N__30553),
            .I(N__30522));
    LocalMux I__5458 (
            .O(N__30550),
            .I(N__30515));
    LocalMux I__5457 (
            .O(N__30547),
            .I(N__30515));
    Span4Mux_v I__5456 (
            .O(N__30544),
            .I(N__30515));
    InMux I__5455 (
            .O(N__30543),
            .I(N__30506));
    InMux I__5454 (
            .O(N__30542),
            .I(N__30506));
    InMux I__5453 (
            .O(N__30541),
            .I(N__30506));
    InMux I__5452 (
            .O(N__30538),
            .I(N__30506));
    Span4Mux_h I__5451 (
            .O(N__30535),
            .I(N__30503));
    LocalMux I__5450 (
            .O(N__30528),
            .I(N__30498));
    Span4Mux_h I__5449 (
            .O(N__30525),
            .I(N__30498));
    LocalMux I__5448 (
            .O(N__30522),
            .I(a_2_repZ0Z1));
    Odrv4 I__5447 (
            .O(N__30515),
            .I(a_2_repZ0Z1));
    LocalMux I__5446 (
            .O(N__30506),
            .I(a_2_repZ0Z1));
    Odrv4 I__5445 (
            .O(N__30503),
            .I(a_2_repZ0Z1));
    Odrv4 I__5444 (
            .O(N__30498),
            .I(a_2_repZ0Z1));
    InMux I__5443 (
            .O(N__30487),
            .I(N__30484));
    LocalMux I__5442 (
            .O(N__30484),
            .I(N__30481));
    Span4Mux_h I__5441 (
            .O(N__30481),
            .I(N__30476));
    InMux I__5440 (
            .O(N__30480),
            .I(N__30473));
    CascadeMux I__5439 (
            .O(N__30479),
            .I(N__30470));
    Span4Mux_h I__5438 (
            .O(N__30476),
            .I(N__30465));
    LocalMux I__5437 (
            .O(N__30473),
            .I(N__30465));
    InMux I__5436 (
            .O(N__30470),
            .I(N__30462));
    Span4Mux_v I__5435 (
            .O(N__30465),
            .I(N__30459));
    LocalMux I__5434 (
            .O(N__30462),
            .I(N__30456));
    Odrv4 I__5433 (
            .O(N__30459),
            .I(r1_15));
    Odrv4 I__5432 (
            .O(N__30456),
            .I(r1_15));
    InMux I__5431 (
            .O(N__30451),
            .I(N__30448));
    LocalMux I__5430 (
            .O(N__30448),
            .I(N__30444));
    InMux I__5429 (
            .O(N__30447),
            .I(N__30441));
    Span4Mux_h I__5428 (
            .O(N__30444),
            .I(N__30438));
    LocalMux I__5427 (
            .O(N__30441),
            .I(N__30435));
    Span4Mux_v I__5426 (
            .O(N__30438),
            .I(N__30429));
    Span4Mux_h I__5425 (
            .O(N__30435),
            .I(N__30429));
    InMux I__5424 (
            .O(N__30434),
            .I(N__30426));
    Odrv4 I__5423 (
            .O(N__30429),
            .I(r5_15));
    LocalMux I__5422 (
            .O(N__30426),
            .I(r5_15));
    CascadeMux I__5421 (
            .O(N__30421),
            .I(TXbuffer_18_10_ns_1_7_cascade_));
    CascadeMux I__5420 (
            .O(N__30418),
            .I(N__30411));
    CascadeMux I__5419 (
            .O(N__30417),
            .I(N__30408));
    CascadeMux I__5418 (
            .O(N__30416),
            .I(N__30405));
    CascadeMux I__5417 (
            .O(N__30415),
            .I(N__30402));
    CascadeMux I__5416 (
            .O(N__30414),
            .I(N__30399));
    InMux I__5415 (
            .O(N__30411),
            .I(N__30389));
    InMux I__5414 (
            .O(N__30408),
            .I(N__30389));
    InMux I__5413 (
            .O(N__30405),
            .I(N__30381));
    InMux I__5412 (
            .O(N__30402),
            .I(N__30381));
    InMux I__5411 (
            .O(N__30399),
            .I(N__30378));
    CascadeMux I__5410 (
            .O(N__30398),
            .I(N__30375));
    CascadeMux I__5409 (
            .O(N__30397),
            .I(N__30372));
    CascadeMux I__5408 (
            .O(N__30396),
            .I(N__30368));
    CascadeMux I__5407 (
            .O(N__30395),
            .I(N__30365));
    CascadeMux I__5406 (
            .O(N__30394),
            .I(N__30361));
    LocalMux I__5405 (
            .O(N__30389),
            .I(N__30356));
    CascadeMux I__5404 (
            .O(N__30388),
            .I(N__30351));
    CascadeMux I__5403 (
            .O(N__30387),
            .I(N__30348));
    InMux I__5402 (
            .O(N__30386),
            .I(N__30345));
    LocalMux I__5401 (
            .O(N__30381),
            .I(N__30340));
    LocalMux I__5400 (
            .O(N__30378),
            .I(N__30340));
    InMux I__5399 (
            .O(N__30375),
            .I(N__30337));
    InMux I__5398 (
            .O(N__30372),
            .I(N__30331));
    InMux I__5397 (
            .O(N__30371),
            .I(N__30331));
    InMux I__5396 (
            .O(N__30368),
            .I(N__30328));
    InMux I__5395 (
            .O(N__30365),
            .I(N__30325));
    CascadeMux I__5394 (
            .O(N__30364),
            .I(N__30321));
    InMux I__5393 (
            .O(N__30361),
            .I(N__30318));
    CascadeMux I__5392 (
            .O(N__30360),
            .I(N__30314));
    CascadeMux I__5391 (
            .O(N__30359),
            .I(N__30311));
    Span4Mux_v I__5390 (
            .O(N__30356),
            .I(N__30306));
    CascadeMux I__5389 (
            .O(N__30355),
            .I(N__30300));
    CascadeMux I__5388 (
            .O(N__30354),
            .I(N__30297));
    InMux I__5387 (
            .O(N__30351),
            .I(N__30292));
    InMux I__5386 (
            .O(N__30348),
            .I(N__30292));
    LocalMux I__5385 (
            .O(N__30345),
            .I(N__30285));
    Span4Mux_h I__5384 (
            .O(N__30340),
            .I(N__30285));
    LocalMux I__5383 (
            .O(N__30337),
            .I(N__30285));
    CascadeMux I__5382 (
            .O(N__30336),
            .I(N__30282));
    LocalMux I__5381 (
            .O(N__30331),
            .I(N__30276));
    LocalMux I__5380 (
            .O(N__30328),
            .I(N__30276));
    LocalMux I__5379 (
            .O(N__30325),
            .I(N__30273));
    CascadeMux I__5378 (
            .O(N__30324),
            .I(N__30270));
    InMux I__5377 (
            .O(N__30321),
            .I(N__30265));
    LocalMux I__5376 (
            .O(N__30318),
            .I(N__30262));
    InMux I__5375 (
            .O(N__30317),
            .I(N__30259));
    InMux I__5374 (
            .O(N__30314),
            .I(N__30256));
    InMux I__5373 (
            .O(N__30311),
            .I(N__30253));
    CascadeMux I__5372 (
            .O(N__30310),
            .I(N__30250));
    InMux I__5371 (
            .O(N__30309),
            .I(N__30247));
    Span4Mux_h I__5370 (
            .O(N__30306),
            .I(N__30244));
    InMux I__5369 (
            .O(N__30305),
            .I(N__30241));
    CascadeMux I__5368 (
            .O(N__30304),
            .I(N__30237));
    InMux I__5367 (
            .O(N__30303),
            .I(N__30230));
    InMux I__5366 (
            .O(N__30300),
            .I(N__30230));
    InMux I__5365 (
            .O(N__30297),
            .I(N__30230));
    LocalMux I__5364 (
            .O(N__30292),
            .I(N__30225));
    Span4Mux_h I__5363 (
            .O(N__30285),
            .I(N__30225));
    InMux I__5362 (
            .O(N__30282),
            .I(N__30220));
    InMux I__5361 (
            .O(N__30281),
            .I(N__30220));
    Span4Mux_h I__5360 (
            .O(N__30276),
            .I(N__30215));
    Span4Mux_v I__5359 (
            .O(N__30273),
            .I(N__30215));
    InMux I__5358 (
            .O(N__30270),
            .I(N__30210));
    InMux I__5357 (
            .O(N__30269),
            .I(N__30210));
    CascadeMux I__5356 (
            .O(N__30268),
            .I(N__30205));
    LocalMux I__5355 (
            .O(N__30265),
            .I(N__30202));
    Span4Mux_v I__5354 (
            .O(N__30262),
            .I(N__30193));
    LocalMux I__5353 (
            .O(N__30259),
            .I(N__30193));
    LocalMux I__5352 (
            .O(N__30256),
            .I(N__30193));
    LocalMux I__5351 (
            .O(N__30253),
            .I(N__30193));
    InMux I__5350 (
            .O(N__30250),
            .I(N__30190));
    LocalMux I__5349 (
            .O(N__30247),
            .I(N__30183));
    Sp12to4 I__5348 (
            .O(N__30244),
            .I(N__30183));
    LocalMux I__5347 (
            .O(N__30241),
            .I(N__30183));
    InMux I__5346 (
            .O(N__30240),
            .I(N__30178));
    InMux I__5345 (
            .O(N__30237),
            .I(N__30178));
    LocalMux I__5344 (
            .O(N__30230),
            .I(N__30175));
    Span4Mux_s1_h I__5343 (
            .O(N__30225),
            .I(N__30172));
    LocalMux I__5342 (
            .O(N__30220),
            .I(N__30167));
    Span4Mux_h I__5341 (
            .O(N__30215),
            .I(N__30167));
    LocalMux I__5340 (
            .O(N__30210),
            .I(N__30164));
    InMux I__5339 (
            .O(N__30209),
            .I(N__30161));
    InMux I__5338 (
            .O(N__30208),
            .I(N__30156));
    InMux I__5337 (
            .O(N__30205),
            .I(N__30156));
    Span4Mux_h I__5336 (
            .O(N__30202),
            .I(N__30153));
    Span4Mux_h I__5335 (
            .O(N__30193),
            .I(N__30150));
    LocalMux I__5334 (
            .O(N__30190),
            .I(N__30145));
    Span12Mux_h I__5333 (
            .O(N__30183),
            .I(N__30145));
    LocalMux I__5332 (
            .O(N__30178),
            .I(N__30138));
    Span4Mux_h I__5331 (
            .O(N__30175),
            .I(N__30138));
    Span4Mux_v I__5330 (
            .O(N__30172),
            .I(N__30138));
    Span4Mux_v I__5329 (
            .O(N__30167),
            .I(N__30135));
    Odrv12 I__5328 (
            .O(N__30164),
            .I(clkdivZ0Z_7));
    LocalMux I__5327 (
            .O(N__30161),
            .I(clkdivZ0Z_7));
    LocalMux I__5326 (
            .O(N__30156),
            .I(clkdivZ0Z_7));
    Odrv4 I__5325 (
            .O(N__30153),
            .I(clkdivZ0Z_7));
    Odrv4 I__5324 (
            .O(N__30150),
            .I(clkdivZ0Z_7));
    Odrv12 I__5323 (
            .O(N__30145),
            .I(clkdivZ0Z_7));
    Odrv4 I__5322 (
            .O(N__30138),
            .I(clkdivZ0Z_7));
    Odrv4 I__5321 (
            .O(N__30135),
            .I(clkdivZ0Z_7));
    InMux I__5320 (
            .O(N__30118),
            .I(N__30114));
    InMux I__5319 (
            .O(N__30117),
            .I(N__30111));
    LocalMux I__5318 (
            .O(N__30114),
            .I(N__30108));
    LocalMux I__5317 (
            .O(N__30111),
            .I(N__30104));
    Span4Mux_h I__5316 (
            .O(N__30108),
            .I(N__30101));
    InMux I__5315 (
            .O(N__30107),
            .I(N__30098));
    Span4Mux_h I__5314 (
            .O(N__30104),
            .I(N__30095));
    Span4Mux_v I__5313 (
            .O(N__30101),
            .I(N__30090));
    LocalMux I__5312 (
            .O(N__30098),
            .I(N__30090));
    Odrv4 I__5311 (
            .O(N__30095),
            .I(r0_15));
    Odrv4 I__5310 (
            .O(N__30090),
            .I(r0_15));
    InMux I__5309 (
            .O(N__30085),
            .I(N__30074));
    InMux I__5308 (
            .O(N__30084),
            .I(N__30074));
    InMux I__5307 (
            .O(N__30083),
            .I(N__30069));
    InMux I__5306 (
            .O(N__30082),
            .I(N__30069));
    CascadeMux I__5305 (
            .O(N__30081),
            .I(N__30055));
    CascadeMux I__5304 (
            .O(N__30080),
            .I(N__30051));
    InMux I__5303 (
            .O(N__30079),
            .I(N__30033));
    LocalMux I__5302 (
            .O(N__30074),
            .I(N__30028));
    LocalMux I__5301 (
            .O(N__30069),
            .I(N__30028));
    InMux I__5300 (
            .O(N__30068),
            .I(N__30021));
    InMux I__5299 (
            .O(N__30067),
            .I(N__30021));
    InMux I__5298 (
            .O(N__30066),
            .I(N__30021));
    InMux I__5297 (
            .O(N__30065),
            .I(N__30012));
    InMux I__5296 (
            .O(N__30064),
            .I(N__30012));
    InMux I__5295 (
            .O(N__30063),
            .I(N__30012));
    InMux I__5294 (
            .O(N__30062),
            .I(N__30012));
    InMux I__5293 (
            .O(N__30061),
            .I(N__30005));
    InMux I__5292 (
            .O(N__30060),
            .I(N__30005));
    InMux I__5291 (
            .O(N__30059),
            .I(N__30005));
    InMux I__5290 (
            .O(N__30058),
            .I(N__29998));
    InMux I__5289 (
            .O(N__30055),
            .I(N__29998));
    InMux I__5288 (
            .O(N__30054),
            .I(N__29998));
    InMux I__5287 (
            .O(N__30051),
            .I(N__29991));
    InMux I__5286 (
            .O(N__30050),
            .I(N__29991));
    InMux I__5285 (
            .O(N__30049),
            .I(N__29991));
    CascadeMux I__5284 (
            .O(N__30048),
            .I(N__29982));
    InMux I__5283 (
            .O(N__30047),
            .I(N__29977));
    InMux I__5282 (
            .O(N__30046),
            .I(N__29977));
    InMux I__5281 (
            .O(N__30045),
            .I(N__29962));
    InMux I__5280 (
            .O(N__30044),
            .I(N__29962));
    InMux I__5279 (
            .O(N__30043),
            .I(N__29953));
    InMux I__5278 (
            .O(N__30042),
            .I(N__29953));
    InMux I__5277 (
            .O(N__30041),
            .I(N__29953));
    InMux I__5276 (
            .O(N__30040),
            .I(N__29953));
    InMux I__5275 (
            .O(N__30039),
            .I(N__29944));
    InMux I__5274 (
            .O(N__30038),
            .I(N__29944));
    InMux I__5273 (
            .O(N__30037),
            .I(N__29944));
    InMux I__5272 (
            .O(N__30036),
            .I(N__29944));
    LocalMux I__5271 (
            .O(N__30033),
            .I(N__29935));
    Span4Mux_v I__5270 (
            .O(N__30028),
            .I(N__29935));
    LocalMux I__5269 (
            .O(N__30021),
            .I(N__29935));
    LocalMux I__5268 (
            .O(N__30012),
            .I(N__29935));
    LocalMux I__5267 (
            .O(N__30005),
            .I(N__29924));
    LocalMux I__5266 (
            .O(N__29998),
            .I(N__29924));
    LocalMux I__5265 (
            .O(N__29991),
            .I(N__29921));
    InMux I__5264 (
            .O(N__29990),
            .I(N__29914));
    InMux I__5263 (
            .O(N__29989),
            .I(N__29914));
    InMux I__5262 (
            .O(N__29988),
            .I(N__29914));
    InMux I__5261 (
            .O(N__29987),
            .I(N__29911));
    InMux I__5260 (
            .O(N__29986),
            .I(N__29904));
    InMux I__5259 (
            .O(N__29985),
            .I(N__29904));
    InMux I__5258 (
            .O(N__29982),
            .I(N__29904));
    LocalMux I__5257 (
            .O(N__29977),
            .I(N__29900));
    InMux I__5256 (
            .O(N__29976),
            .I(N__29895));
    InMux I__5255 (
            .O(N__29975),
            .I(N__29895));
    InMux I__5254 (
            .O(N__29974),
            .I(N__29888));
    InMux I__5253 (
            .O(N__29973),
            .I(N__29888));
    InMux I__5252 (
            .O(N__29972),
            .I(N__29888));
    InMux I__5251 (
            .O(N__29971),
            .I(N__29881));
    InMux I__5250 (
            .O(N__29970),
            .I(N__29876));
    InMux I__5249 (
            .O(N__29969),
            .I(N__29876));
    InMux I__5248 (
            .O(N__29968),
            .I(N__29871));
    InMux I__5247 (
            .O(N__29967),
            .I(N__29871));
    LocalMux I__5246 (
            .O(N__29962),
            .I(N__29868));
    LocalMux I__5245 (
            .O(N__29953),
            .I(N__29865));
    LocalMux I__5244 (
            .O(N__29944),
            .I(N__29860));
    Span4Mux_h I__5243 (
            .O(N__29935),
            .I(N__29860));
    InMux I__5242 (
            .O(N__29934),
            .I(N__29856));
    InMux I__5241 (
            .O(N__29933),
            .I(N__29845));
    InMux I__5240 (
            .O(N__29932),
            .I(N__29845));
    InMux I__5239 (
            .O(N__29931),
            .I(N__29845));
    InMux I__5238 (
            .O(N__29930),
            .I(N__29845));
    InMux I__5237 (
            .O(N__29929),
            .I(N__29845));
    Sp12to4 I__5236 (
            .O(N__29924),
            .I(N__29839));
    Span4Mux_h I__5235 (
            .O(N__29921),
            .I(N__29834));
    LocalMux I__5234 (
            .O(N__29914),
            .I(N__29834));
    LocalMux I__5233 (
            .O(N__29911),
            .I(N__29831));
    LocalMux I__5232 (
            .O(N__29904),
            .I(N__29828));
    InMux I__5231 (
            .O(N__29903),
            .I(N__29825));
    Span4Mux_v I__5230 (
            .O(N__29900),
            .I(N__29822));
    LocalMux I__5229 (
            .O(N__29895),
            .I(N__29819));
    LocalMux I__5228 (
            .O(N__29888),
            .I(N__29816));
    InMux I__5227 (
            .O(N__29887),
            .I(N__29811));
    InMux I__5226 (
            .O(N__29886),
            .I(N__29811));
    InMux I__5225 (
            .O(N__29885),
            .I(N__29806));
    InMux I__5224 (
            .O(N__29884),
            .I(N__29806));
    LocalMux I__5223 (
            .O(N__29881),
            .I(N__29797));
    LocalMux I__5222 (
            .O(N__29876),
            .I(N__29797));
    LocalMux I__5221 (
            .O(N__29871),
            .I(N__29797));
    Span4Mux_v I__5220 (
            .O(N__29868),
            .I(N__29797));
    Span4Mux_v I__5219 (
            .O(N__29865),
            .I(N__29792));
    Span4Mux_h I__5218 (
            .O(N__29860),
            .I(N__29792));
    InMux I__5217 (
            .O(N__29859),
            .I(N__29789));
    LocalMux I__5216 (
            .O(N__29856),
            .I(N__29784));
    LocalMux I__5215 (
            .O(N__29845),
            .I(N__29784));
    InMux I__5214 (
            .O(N__29844),
            .I(N__29779));
    InMux I__5213 (
            .O(N__29843),
            .I(N__29779));
    InMux I__5212 (
            .O(N__29842),
            .I(N__29776));
    Span12Mux_h I__5211 (
            .O(N__29839),
            .I(N__29773));
    Span4Mux_h I__5210 (
            .O(N__29834),
            .I(N__29770));
    Span4Mux_h I__5209 (
            .O(N__29831),
            .I(N__29763));
    Span4Mux_h I__5208 (
            .O(N__29828),
            .I(N__29763));
    LocalMux I__5207 (
            .O(N__29825),
            .I(N__29763));
    Span4Mux_h I__5206 (
            .O(N__29822),
            .I(N__29756));
    Span4Mux_v I__5205 (
            .O(N__29819),
            .I(N__29756));
    Span4Mux_h I__5204 (
            .O(N__29816),
            .I(N__29756));
    LocalMux I__5203 (
            .O(N__29811),
            .I(N__29747));
    LocalMux I__5202 (
            .O(N__29806),
            .I(N__29747));
    Span4Mux_h I__5201 (
            .O(N__29797),
            .I(N__29747));
    Span4Mux_v I__5200 (
            .O(N__29792),
            .I(N__29747));
    LocalMux I__5199 (
            .O(N__29789),
            .I(clkdivZ0Z_6));
    Odrv12 I__5198 (
            .O(N__29784),
            .I(clkdivZ0Z_6));
    LocalMux I__5197 (
            .O(N__29779),
            .I(clkdivZ0Z_6));
    LocalMux I__5196 (
            .O(N__29776),
            .I(clkdivZ0Z_6));
    Odrv12 I__5195 (
            .O(N__29773),
            .I(clkdivZ0Z_6));
    Odrv4 I__5194 (
            .O(N__29770),
            .I(clkdivZ0Z_6));
    Odrv4 I__5193 (
            .O(N__29763),
            .I(clkdivZ0Z_6));
    Odrv4 I__5192 (
            .O(N__29756),
            .I(clkdivZ0Z_6));
    Odrv4 I__5191 (
            .O(N__29747),
            .I(clkdivZ0Z_6));
    CascadeMux I__5190 (
            .O(N__29728),
            .I(TXbuffer_18_3_ns_1_7_cascade_));
    InMux I__5189 (
            .O(N__29725),
            .I(N__29722));
    LocalMux I__5188 (
            .O(N__29722),
            .I(N__29718));
    InMux I__5187 (
            .O(N__29721),
            .I(N__29715));
    Span4Mux_v I__5186 (
            .O(N__29718),
            .I(N__29712));
    LocalMux I__5185 (
            .O(N__29715),
            .I(N__29709));
    Span4Mux_v I__5184 (
            .O(N__29712),
            .I(N__29705));
    Span4Mux_s2_h I__5183 (
            .O(N__29709),
            .I(N__29702));
    InMux I__5182 (
            .O(N__29708),
            .I(N__29699));
    Sp12to4 I__5181 (
            .O(N__29705),
            .I(N__29696));
    Span4Mux_h I__5180 (
            .O(N__29702),
            .I(N__29693));
    LocalMux I__5179 (
            .O(N__29699),
            .I(N__29690));
    Odrv12 I__5178 (
            .O(N__29696),
            .I(r4_15));
    Odrv4 I__5177 (
            .O(N__29693),
            .I(r4_15));
    Odrv4 I__5176 (
            .O(N__29690),
            .I(r4_15));
    InMux I__5175 (
            .O(N__29683),
            .I(N__29680));
    LocalMux I__5174 (
            .O(N__29680),
            .I(N__29677));
    Span4Mux_h I__5173 (
            .O(N__29677),
            .I(N__29671));
    InMux I__5172 (
            .O(N__29676),
            .I(N__29665));
    InMux I__5171 (
            .O(N__29675),
            .I(N__29662));
    CascadeMux I__5170 (
            .O(N__29674),
            .I(N__29658));
    Span4Mux_h I__5169 (
            .O(N__29671),
            .I(N__29655));
    InMux I__5168 (
            .O(N__29670),
            .I(N__29652));
    InMux I__5167 (
            .O(N__29669),
            .I(N__29649));
    InMux I__5166 (
            .O(N__29668),
            .I(N__29646));
    LocalMux I__5165 (
            .O(N__29665),
            .I(N__29643));
    LocalMux I__5164 (
            .O(N__29662),
            .I(N__29640));
    InMux I__5163 (
            .O(N__29661),
            .I(N__29637));
    InMux I__5162 (
            .O(N__29658),
            .I(N__29634));
    Span4Mux_h I__5161 (
            .O(N__29655),
            .I(N__29629));
    LocalMux I__5160 (
            .O(N__29652),
            .I(N__29629));
    LocalMux I__5159 (
            .O(N__29649),
            .I(N__29626));
    LocalMux I__5158 (
            .O(N__29646),
            .I(N__29623));
    Span12Mux_h I__5157 (
            .O(N__29643),
            .I(N__29619));
    Span12Mux_v I__5156 (
            .O(N__29640),
            .I(N__29616));
    LocalMux I__5155 (
            .O(N__29637),
            .I(N__29609));
    LocalMux I__5154 (
            .O(N__29634),
            .I(N__29609));
    Span4Mux_v I__5153 (
            .O(N__29629),
            .I(N__29609));
    Span4Mux_h I__5152 (
            .O(N__29626),
            .I(N__29606));
    Span4Mux_h I__5151 (
            .O(N__29623),
            .I(N__29603));
    InMux I__5150 (
            .O(N__29622),
            .I(N__29600));
    Odrv12 I__5149 (
            .O(N__29619),
            .I(clkdivZ0Z_5));
    Odrv12 I__5148 (
            .O(N__29616),
            .I(clkdivZ0Z_5));
    Odrv4 I__5147 (
            .O(N__29609),
            .I(clkdivZ0Z_5));
    Odrv4 I__5146 (
            .O(N__29606),
            .I(clkdivZ0Z_5));
    Odrv4 I__5145 (
            .O(N__29603),
            .I(clkdivZ0Z_5));
    LocalMux I__5144 (
            .O(N__29600),
            .I(clkdivZ0Z_5));
    CascadeMux I__5143 (
            .O(N__29587),
            .I(TXbuffer_RNO_5Z0Z_7_cascade_));
    InMux I__5142 (
            .O(N__29584),
            .I(N__29581));
    LocalMux I__5141 (
            .O(N__29581),
            .I(N__29578));
    Span4Mux_v I__5140 (
            .O(N__29578),
            .I(N__29575));
    Span4Mux_v I__5139 (
            .O(N__29575),
            .I(N__29572));
    Span4Mux_h I__5138 (
            .O(N__29572),
            .I(N__29569));
    Odrv4 I__5137 (
            .O(N__29569),
            .I(TXbuffer_RNO_6Z0Z_7));
    CascadeMux I__5136 (
            .O(N__29566),
            .I(\ALU.a_3_ns_1_1_cascade_ ));
    CascadeMux I__5135 (
            .O(N__29563),
            .I(N__29559));
    InMux I__5134 (
            .O(N__29562),
            .I(N__29556));
    InMux I__5133 (
            .O(N__29559),
            .I(N__29553));
    LocalMux I__5132 (
            .O(N__29556),
            .I(N__29550));
    LocalMux I__5131 (
            .O(N__29553),
            .I(N__29547));
    Span4Mux_v I__5130 (
            .O(N__29550),
            .I(N__29544));
    Odrv4 I__5129 (
            .O(N__29547),
            .I(\ALU.a3_b_2 ));
    Odrv4 I__5128 (
            .O(N__29544),
            .I(\ALU.a3_b_2 ));
    CascadeMux I__5127 (
            .O(N__29539),
            .I(\ALU.rshift_3_ns_1_7_cascade_ ));
    CascadeMux I__5126 (
            .O(N__29536),
            .I(\ALU.b_3_ns_1_7_cascade_ ));
    InMux I__5125 (
            .O(N__29533),
            .I(N__29530));
    LocalMux I__5124 (
            .O(N__29530),
            .I(N__29527));
    Span4Mux_h I__5123 (
            .O(N__29527),
            .I(N__29524));
    Span4Mux_h I__5122 (
            .O(N__29524),
            .I(N__29521));
    Odrv4 I__5121 (
            .O(N__29521),
            .I(\ALU.r4_RNI82OE1Z0Z_7 ));
    InMux I__5120 (
            .O(N__29518),
            .I(N__29509));
    InMux I__5119 (
            .O(N__29517),
            .I(N__29509));
    CascadeMux I__5118 (
            .O(N__29516),
            .I(N__29504));
    InMux I__5117 (
            .O(N__29515),
            .I(N__29499));
    InMux I__5116 (
            .O(N__29514),
            .I(N__29499));
    LocalMux I__5115 (
            .O(N__29509),
            .I(N__29496));
    InMux I__5114 (
            .O(N__29508),
            .I(N__29493));
    InMux I__5113 (
            .O(N__29507),
            .I(N__29490));
    InMux I__5112 (
            .O(N__29504),
            .I(N__29483));
    LocalMux I__5111 (
            .O(N__29499),
            .I(N__29476));
    Span4Mux_h I__5110 (
            .O(N__29496),
            .I(N__29476));
    LocalMux I__5109 (
            .O(N__29493),
            .I(N__29471));
    LocalMux I__5108 (
            .O(N__29490),
            .I(N__29471));
    InMux I__5107 (
            .O(N__29489),
            .I(N__29462));
    InMux I__5106 (
            .O(N__29488),
            .I(N__29462));
    InMux I__5105 (
            .O(N__29487),
            .I(N__29462));
    InMux I__5104 (
            .O(N__29486),
            .I(N__29462));
    LocalMux I__5103 (
            .O(N__29483),
            .I(N__29459));
    InMux I__5102 (
            .O(N__29482),
            .I(N__29454));
    InMux I__5101 (
            .O(N__29481),
            .I(N__29454));
    Span4Mux_h I__5100 (
            .O(N__29476),
            .I(N__29451));
    Odrv4 I__5099 (
            .O(N__29471),
            .I(b_0_repZ0Z2));
    LocalMux I__5098 (
            .O(N__29462),
            .I(b_0_repZ0Z2));
    Odrv12 I__5097 (
            .O(N__29459),
            .I(b_0_repZ0Z2));
    LocalMux I__5096 (
            .O(N__29454),
            .I(b_0_repZ0Z2));
    Odrv4 I__5095 (
            .O(N__29451),
            .I(b_0_repZ0Z2));
    InMux I__5094 (
            .O(N__29440),
            .I(N__29436));
    InMux I__5093 (
            .O(N__29439),
            .I(N__29433));
    LocalMux I__5092 (
            .O(N__29436),
            .I(N__29430));
    LocalMux I__5091 (
            .O(N__29433),
            .I(N__29426));
    Span4Mux_h I__5090 (
            .O(N__29430),
            .I(N__29423));
    InMux I__5089 (
            .O(N__29429),
            .I(N__29420));
    Span4Mux_h I__5088 (
            .O(N__29426),
            .I(N__29417));
    Span4Mux_v I__5087 (
            .O(N__29423),
            .I(N__29414));
    LocalMux I__5086 (
            .O(N__29420),
            .I(r7_1));
    Odrv4 I__5085 (
            .O(N__29417),
            .I(r7_1));
    Odrv4 I__5084 (
            .O(N__29414),
            .I(r7_1));
    InMux I__5083 (
            .O(N__29407),
            .I(N__29403));
    InMux I__5082 (
            .O(N__29406),
            .I(N__29400));
    LocalMux I__5081 (
            .O(N__29403),
            .I(N__29397));
    LocalMux I__5080 (
            .O(N__29400),
            .I(N__29393));
    Span4Mux_h I__5079 (
            .O(N__29397),
            .I(N__29390));
    InMux I__5078 (
            .O(N__29396),
            .I(N__29387));
    Span12Mux_v I__5077 (
            .O(N__29393),
            .I(N__29384));
    Span4Mux_v I__5076 (
            .O(N__29390),
            .I(N__29381));
    LocalMux I__5075 (
            .O(N__29387),
            .I(r6_1));
    Odrv12 I__5074 (
            .O(N__29384),
            .I(r6_1));
    Odrv4 I__5073 (
            .O(N__29381),
            .I(r6_1));
    InMux I__5072 (
            .O(N__29374),
            .I(N__29371));
    LocalMux I__5071 (
            .O(N__29371),
            .I(N__29368));
    Odrv12 I__5070 (
            .O(N__29368),
            .I(\ALU.r6_RNIC9P41Z0Z_1 ));
    InMux I__5069 (
            .O(N__29365),
            .I(N__29361));
    InMux I__5068 (
            .O(N__29364),
            .I(N__29356));
    LocalMux I__5067 (
            .O(N__29361),
            .I(N__29353));
    InMux I__5066 (
            .O(N__29360),
            .I(N__29350));
    InMux I__5065 (
            .O(N__29359),
            .I(N__29347));
    LocalMux I__5064 (
            .O(N__29356),
            .I(N__29344));
    Span4Mux_h I__5063 (
            .O(N__29353),
            .I(N__29339));
    LocalMux I__5062 (
            .O(N__29350),
            .I(N__29339));
    LocalMux I__5061 (
            .O(N__29347),
            .I(\ALU.r6_RNIE5FT1Z0Z_2 ));
    Odrv4 I__5060 (
            .O(N__29344),
            .I(\ALU.r6_RNIE5FT1Z0Z_2 ));
    Odrv4 I__5059 (
            .O(N__29339),
            .I(\ALU.r6_RNIE5FT1Z0Z_2 ));
    InMux I__5058 (
            .O(N__29332),
            .I(N__29326));
    InMux I__5057 (
            .O(N__29331),
            .I(N__29326));
    LocalMux I__5056 (
            .O(N__29326),
            .I(N__29323));
    Odrv4 I__5055 (
            .O(N__29323),
            .I(\ALU.madd_13 ));
    CascadeMux I__5054 (
            .O(N__29320),
            .I(N__29316));
    CascadeMux I__5053 (
            .O(N__29319),
            .I(N__29313));
    InMux I__5052 (
            .O(N__29316),
            .I(N__29310));
    InMux I__5051 (
            .O(N__29313),
            .I(N__29307));
    LocalMux I__5050 (
            .O(N__29310),
            .I(N__29304));
    LocalMux I__5049 (
            .O(N__29307),
            .I(\ALU.a2_b_0 ));
    Odrv12 I__5048 (
            .O(N__29304),
            .I(\ALU.a2_b_0 ));
    CascadeMux I__5047 (
            .O(N__29299),
            .I(N__29296));
    InMux I__5046 (
            .O(N__29296),
            .I(N__29293));
    LocalMux I__5045 (
            .O(N__29293),
            .I(\ALU.madd_3 ));
    InMux I__5044 (
            .O(N__29290),
            .I(N__29284));
    InMux I__5043 (
            .O(N__29289),
            .I(N__29284));
    LocalMux I__5042 (
            .O(N__29284),
            .I(N__29281));
    Odrv12 I__5041 (
            .O(N__29281),
            .I(\ALU.madd_4 ));
    CascadeMux I__5040 (
            .O(N__29278),
            .I(\ALU.madd_3_cascade_ ));
    InMux I__5039 (
            .O(N__29275),
            .I(N__29269));
    InMux I__5038 (
            .O(N__29274),
            .I(N__29269));
    LocalMux I__5037 (
            .O(N__29269),
            .I(\ALU.a0_b_3 ));
    InMux I__5036 (
            .O(N__29266),
            .I(N__29263));
    LocalMux I__5035 (
            .O(N__29263),
            .I(N__29259));
    InMux I__5034 (
            .O(N__29262),
            .I(N__29256));
    Span4Mux_s2_v I__5033 (
            .O(N__29259),
            .I(N__29251));
    LocalMux I__5032 (
            .O(N__29256),
            .I(N__29251));
    Span4Mux_v I__5031 (
            .O(N__29251),
            .I(N__29248));
    Odrv4 I__5030 (
            .O(N__29248),
            .I(\ALU.madd_66 ));
    CascadeMux I__5029 (
            .O(N__29245),
            .I(N__29241));
    CascadeMux I__5028 (
            .O(N__29244),
            .I(N__29238));
    InMux I__5027 (
            .O(N__29241),
            .I(N__29234));
    InMux I__5026 (
            .O(N__29238),
            .I(N__29231));
    InMux I__5025 (
            .O(N__29237),
            .I(N__29228));
    LocalMux I__5024 (
            .O(N__29234),
            .I(N__29221));
    LocalMux I__5023 (
            .O(N__29231),
            .I(N__29221));
    LocalMux I__5022 (
            .O(N__29228),
            .I(N__29216));
    CascadeMux I__5021 (
            .O(N__29227),
            .I(N__29212));
    CascadeMux I__5020 (
            .O(N__29226),
            .I(N__29209));
    Span4Mux_v I__5019 (
            .O(N__29221),
            .I(N__29203));
    InMux I__5018 (
            .O(N__29220),
            .I(N__29199));
    InMux I__5017 (
            .O(N__29219),
            .I(N__29196));
    Span4Mux_s3_v I__5016 (
            .O(N__29216),
            .I(N__29193));
    InMux I__5015 (
            .O(N__29215),
            .I(N__29190));
    InMux I__5014 (
            .O(N__29212),
            .I(N__29187));
    InMux I__5013 (
            .O(N__29209),
            .I(N__29184));
    CascadeMux I__5012 (
            .O(N__29208),
            .I(N__29180));
    InMux I__5011 (
            .O(N__29207),
            .I(N__29177));
    InMux I__5010 (
            .O(N__29206),
            .I(N__29174));
    Span4Mux_v I__5009 (
            .O(N__29203),
            .I(N__29171));
    InMux I__5008 (
            .O(N__29202),
            .I(N__29168));
    LocalMux I__5007 (
            .O(N__29199),
            .I(N__29161));
    LocalMux I__5006 (
            .O(N__29196),
            .I(N__29161));
    Span4Mux_h I__5005 (
            .O(N__29193),
            .I(N__29161));
    LocalMux I__5004 (
            .O(N__29190),
            .I(N__29157));
    LocalMux I__5003 (
            .O(N__29187),
            .I(N__29151));
    LocalMux I__5002 (
            .O(N__29184),
            .I(N__29151));
    InMux I__5001 (
            .O(N__29183),
            .I(N__29146));
    InMux I__5000 (
            .O(N__29180),
            .I(N__29146));
    LocalMux I__4999 (
            .O(N__29177),
            .I(N__29141));
    LocalMux I__4998 (
            .O(N__29174),
            .I(N__29141));
    Sp12to4 I__4997 (
            .O(N__29171),
            .I(N__29136));
    LocalMux I__4996 (
            .O(N__29168),
            .I(N__29136));
    Sp12to4 I__4995 (
            .O(N__29161),
            .I(N__29133));
    InMux I__4994 (
            .O(N__29160),
            .I(N__29130));
    Span4Mux_v I__4993 (
            .O(N__29157),
            .I(N__29127));
    InMux I__4992 (
            .O(N__29156),
            .I(N__29124));
    Span12Mux_s5_h I__4991 (
            .O(N__29151),
            .I(N__29119));
    LocalMux I__4990 (
            .O(N__29146),
            .I(N__29119));
    Span12Mux_v I__4989 (
            .O(N__29141),
            .I(N__29112));
    Span12Mux_s4_h I__4988 (
            .O(N__29136),
            .I(N__29112));
    Span12Mux_s8_v I__4987 (
            .O(N__29133),
            .I(N__29112));
    LocalMux I__4986 (
            .O(N__29130),
            .I(a_1_repZ0Z1));
    Odrv4 I__4985 (
            .O(N__29127),
            .I(a_1_repZ0Z1));
    LocalMux I__4984 (
            .O(N__29124),
            .I(a_1_repZ0Z1));
    Odrv12 I__4983 (
            .O(N__29119),
            .I(a_1_repZ0Z1));
    Odrv12 I__4982 (
            .O(N__29112),
            .I(a_1_repZ0Z1));
    InMux I__4981 (
            .O(N__29101),
            .I(N__29097));
    InMux I__4980 (
            .O(N__29100),
            .I(N__29091));
    LocalMux I__4979 (
            .O(N__29097),
            .I(N__29088));
    InMux I__4978 (
            .O(N__29096),
            .I(N__29081));
    InMux I__4977 (
            .O(N__29095),
            .I(N__29081));
    InMux I__4976 (
            .O(N__29094),
            .I(N__29081));
    LocalMux I__4975 (
            .O(N__29091),
            .I(N__29073));
    Span4Mux_s2_v I__4974 (
            .O(N__29088),
            .I(N__29068));
    LocalMux I__4973 (
            .O(N__29081),
            .I(N__29068));
    InMux I__4972 (
            .O(N__29080),
            .I(N__29065));
    InMux I__4971 (
            .O(N__29079),
            .I(N__29062));
    InMux I__4970 (
            .O(N__29078),
            .I(N__29059));
    InMux I__4969 (
            .O(N__29077),
            .I(N__29056));
    InMux I__4968 (
            .O(N__29076),
            .I(N__29053));
    Span4Mux_s2_v I__4967 (
            .O(N__29073),
            .I(N__29048));
    Span4Mux_h I__4966 (
            .O(N__29068),
            .I(N__29048));
    LocalMux I__4965 (
            .O(N__29065),
            .I(N__29045));
    LocalMux I__4964 (
            .O(N__29062),
            .I(N__29040));
    LocalMux I__4963 (
            .O(N__29059),
            .I(N__29040));
    LocalMux I__4962 (
            .O(N__29056),
            .I(N__29037));
    LocalMux I__4961 (
            .O(N__29053),
            .I(N__29034));
    Span4Mux_v I__4960 (
            .O(N__29048),
            .I(N__29031));
    Span4Mux_h I__4959 (
            .O(N__29045),
            .I(N__29026));
    Span4Mux_s3_v I__4958 (
            .O(N__29040),
            .I(N__29026));
    Sp12to4 I__4957 (
            .O(N__29037),
            .I(N__29021));
    Span12Mux_s7_v I__4956 (
            .O(N__29034),
            .I(N__29021));
    Odrv4 I__4955 (
            .O(N__29031),
            .I(\ALU.r6_RNIASIB2Z0Z_5 ));
    Odrv4 I__4954 (
            .O(N__29026),
            .I(\ALU.r6_RNIASIB2Z0Z_5 ));
    Odrv12 I__4953 (
            .O(N__29021),
            .I(\ALU.r6_RNIASIB2Z0Z_5 ));
    CascadeMux I__4952 (
            .O(N__29014),
            .I(N__29010));
    InMux I__4951 (
            .O(N__29013),
            .I(N__29006));
    InMux I__4950 (
            .O(N__29010),
            .I(N__29000));
    InMux I__4949 (
            .O(N__29009),
            .I(N__28994));
    LocalMux I__4948 (
            .O(N__29006),
            .I(N__28991));
    InMux I__4947 (
            .O(N__29005),
            .I(N__28988));
    InMux I__4946 (
            .O(N__29004),
            .I(N__28985));
    InMux I__4945 (
            .O(N__29003),
            .I(N__28982));
    LocalMux I__4944 (
            .O(N__29000),
            .I(N__28979));
    InMux I__4943 (
            .O(N__28999),
            .I(N__28971));
    InMux I__4942 (
            .O(N__28998),
            .I(N__28971));
    InMux I__4941 (
            .O(N__28997),
            .I(N__28971));
    LocalMux I__4940 (
            .O(N__28994),
            .I(N__28968));
    Span4Mux_h I__4939 (
            .O(N__28991),
            .I(N__28963));
    LocalMux I__4938 (
            .O(N__28988),
            .I(N__28963));
    LocalMux I__4937 (
            .O(N__28985),
            .I(N__28960));
    LocalMux I__4936 (
            .O(N__28982),
            .I(N__28957));
    Span4Mux_v I__4935 (
            .O(N__28979),
            .I(N__28954));
    InMux I__4934 (
            .O(N__28978),
            .I(N__28951));
    LocalMux I__4933 (
            .O(N__28971),
            .I(N__28946));
    Span4Mux_h I__4932 (
            .O(N__28968),
            .I(N__28946));
    Span4Mux_s1_v I__4931 (
            .O(N__28963),
            .I(N__28943));
    Span4Mux_v I__4930 (
            .O(N__28960),
            .I(N__28940));
    Span4Mux_v I__4929 (
            .O(N__28957),
            .I(N__28935));
    Span4Mux_v I__4928 (
            .O(N__28954),
            .I(N__28935));
    LocalMux I__4927 (
            .O(N__28951),
            .I(N__28930));
    Sp12to4 I__4926 (
            .O(N__28946),
            .I(N__28930));
    Span4Mux_v I__4925 (
            .O(N__28943),
            .I(N__28925));
    Span4Mux_h I__4924 (
            .O(N__28940),
            .I(N__28925));
    Odrv4 I__4923 (
            .O(N__28935),
            .I(\ALU.r4_RNI24Q22Z0Z_5 ));
    Odrv12 I__4922 (
            .O(N__28930),
            .I(\ALU.r4_RNI24Q22Z0Z_5 ));
    Odrv4 I__4921 (
            .O(N__28925),
            .I(\ALU.r4_RNI24Q22Z0Z_5 ));
    InMux I__4920 (
            .O(N__28918),
            .I(N__28909));
    InMux I__4919 (
            .O(N__28917),
            .I(N__28909));
    InMux I__4918 (
            .O(N__28916),
            .I(N__28909));
    LocalMux I__4917 (
            .O(N__28909),
            .I(\ALU.a0_b_4 ));
    InMux I__4916 (
            .O(N__28906),
            .I(N__28903));
    LocalMux I__4915 (
            .O(N__28903),
            .I(N__28900));
    Span4Mux_s3_v I__4914 (
            .O(N__28900),
            .I(N__28897));
    Odrv4 I__4913 (
            .O(N__28897),
            .I(\ALU.un2_addsub_axb_2 ));
    InMux I__4912 (
            .O(N__28894),
            .I(N__28887));
    InMux I__4911 (
            .O(N__28893),
            .I(N__28887));
    InMux I__4910 (
            .O(N__28892),
            .I(N__28884));
    LocalMux I__4909 (
            .O(N__28887),
            .I(N__28881));
    LocalMux I__4908 (
            .O(N__28884),
            .I(\ALU.madd_56 ));
    Odrv4 I__4907 (
            .O(N__28881),
            .I(\ALU.madd_56 ));
    InMux I__4906 (
            .O(N__28876),
            .I(N__28873));
    LocalMux I__4905 (
            .O(N__28873),
            .I(N__28870));
    Span4Mux_h I__4904 (
            .O(N__28870),
            .I(N__28865));
    InMux I__4903 (
            .O(N__28869),
            .I(N__28860));
    InMux I__4902 (
            .O(N__28868),
            .I(N__28860));
    Odrv4 I__4901 (
            .O(N__28865),
            .I(\ALU.madd_45 ));
    LocalMux I__4900 (
            .O(N__28860),
            .I(\ALU.madd_45 ));
    CascadeMux I__4899 (
            .O(N__28855),
            .I(N__28852));
    InMux I__4898 (
            .O(N__28852),
            .I(N__28849));
    LocalMux I__4897 (
            .O(N__28849),
            .I(N__28846));
    Span4Mux_h I__4896 (
            .O(N__28846),
            .I(N__28843));
    Odrv4 I__4895 (
            .O(N__28843),
            .I(\ALU.madd_cry_6_ma ));
    InMux I__4894 (
            .O(N__28840),
            .I(N__28835));
    CascadeMux I__4893 (
            .O(N__28839),
            .I(N__28832));
    InMux I__4892 (
            .O(N__28838),
            .I(N__28829));
    LocalMux I__4891 (
            .O(N__28835),
            .I(N__28826));
    InMux I__4890 (
            .O(N__28832),
            .I(N__28823));
    LocalMux I__4889 (
            .O(N__28829),
            .I(N__28820));
    Span4Mux_v I__4888 (
            .O(N__28826),
            .I(N__28817));
    LocalMux I__4887 (
            .O(N__28823),
            .I(N__28814));
    Span4Mux_s3_h I__4886 (
            .O(N__28820),
            .I(N__28811));
    Span4Mux_h I__4885 (
            .O(N__28817),
            .I(N__28808));
    Span4Mux_h I__4884 (
            .O(N__28814),
            .I(N__28805));
    Odrv4 I__4883 (
            .O(N__28811),
            .I(r3_0));
    Odrv4 I__4882 (
            .O(N__28808),
            .I(r3_0));
    Odrv4 I__4881 (
            .O(N__28805),
            .I(r3_0));
    InMux I__4880 (
            .O(N__28798),
            .I(N__28795));
    LocalMux I__4879 (
            .O(N__28795),
            .I(N__28792));
    Span4Mux_v I__4878 (
            .O(N__28792),
            .I(N__28785));
    InMux I__4877 (
            .O(N__28791),
            .I(N__28772));
    InMux I__4876 (
            .O(N__28790),
            .I(N__28772));
    InMux I__4875 (
            .O(N__28789),
            .I(N__28772));
    InMux I__4874 (
            .O(N__28788),
            .I(N__28772));
    Span4Mux_h I__4873 (
            .O(N__28785),
            .I(N__28769));
    InMux I__4872 (
            .O(N__28784),
            .I(N__28760));
    InMux I__4871 (
            .O(N__28783),
            .I(N__28760));
    InMux I__4870 (
            .O(N__28782),
            .I(N__28760));
    InMux I__4869 (
            .O(N__28781),
            .I(N__28760));
    LocalMux I__4868 (
            .O(N__28772),
            .I(a_0_repZ0Z2));
    Odrv4 I__4867 (
            .O(N__28769),
            .I(a_0_repZ0Z2));
    LocalMux I__4866 (
            .O(N__28760),
            .I(a_0_repZ0Z2));
    InMux I__4865 (
            .O(N__28753),
            .I(N__28750));
    LocalMux I__4864 (
            .O(N__28750),
            .I(N__28747));
    Span4Mux_s3_v I__4863 (
            .O(N__28747),
            .I(N__28744));
    Odrv4 I__4862 (
            .O(N__28744),
            .I(\ALU.r2_RNI18BOZ0Z_0 ));
    InMux I__4861 (
            .O(N__28741),
            .I(N__28737));
    InMux I__4860 (
            .O(N__28740),
            .I(N__28734));
    LocalMux I__4859 (
            .O(N__28737),
            .I(N__28731));
    LocalMux I__4858 (
            .O(N__28734),
            .I(N__28728));
    Sp12to4 I__4857 (
            .O(N__28731),
            .I(N__28725));
    Span4Mux_v I__4856 (
            .O(N__28728),
            .I(N__28721));
    Span12Mux_v I__4855 (
            .O(N__28725),
            .I(N__28718));
    InMux I__4854 (
            .O(N__28724),
            .I(N__28715));
    Span4Mux_h I__4853 (
            .O(N__28721),
            .I(N__28712));
    Odrv12 I__4852 (
            .O(N__28718),
            .I(r2_0));
    LocalMux I__4851 (
            .O(N__28715),
            .I(r2_0));
    Odrv4 I__4850 (
            .O(N__28712),
            .I(r2_0));
    InMux I__4849 (
            .O(N__28705),
            .I(N__28702));
    LocalMux I__4848 (
            .O(N__28702),
            .I(N__28697));
    InMux I__4847 (
            .O(N__28701),
            .I(N__28694));
    CascadeMux I__4846 (
            .O(N__28700),
            .I(N__28691));
    Span4Mux_h I__4845 (
            .O(N__28697),
            .I(N__28688));
    LocalMux I__4844 (
            .O(N__28694),
            .I(N__28685));
    InMux I__4843 (
            .O(N__28691),
            .I(N__28682));
    Span4Mux_h I__4842 (
            .O(N__28688),
            .I(N__28679));
    Span4Mux_h I__4841 (
            .O(N__28685),
            .I(N__28676));
    LocalMux I__4840 (
            .O(N__28682),
            .I(N__28673));
    Span4Mux_v I__4839 (
            .O(N__28679),
            .I(N__28670));
    Odrv4 I__4838 (
            .O(N__28676),
            .I(r3_1));
    Odrv4 I__4837 (
            .O(N__28673),
            .I(r3_1));
    Odrv4 I__4836 (
            .O(N__28670),
            .I(r3_1));
    InMux I__4835 (
            .O(N__28663),
            .I(N__28659));
    InMux I__4834 (
            .O(N__28662),
            .I(N__28656));
    LocalMux I__4833 (
            .O(N__28659),
            .I(N__28653));
    LocalMux I__4832 (
            .O(N__28656),
            .I(N__28649));
    Span12Mux_h I__4831 (
            .O(N__28653),
            .I(N__28646));
    InMux I__4830 (
            .O(N__28652),
            .I(N__28643));
    Odrv4 I__4829 (
            .O(N__28649),
            .I(r2_1));
    Odrv12 I__4828 (
            .O(N__28646),
            .I(r2_1));
    LocalMux I__4827 (
            .O(N__28643),
            .I(r2_1));
    CascadeMux I__4826 (
            .O(N__28636),
            .I(N__28633));
    InMux I__4825 (
            .O(N__28633),
            .I(N__28630));
    LocalMux I__4824 (
            .O(N__28630),
            .I(N__28627));
    Sp12to4 I__4823 (
            .O(N__28627),
            .I(N__28624));
    Odrv12 I__4822 (
            .O(N__28624),
            .I(\ALU.r2_RNI4H0SZ0Z_1 ));
    InMux I__4821 (
            .O(N__28621),
            .I(N__28618));
    LocalMux I__4820 (
            .O(N__28618),
            .I(N__28614));
    InMux I__4819 (
            .O(N__28617),
            .I(N__28611));
    Odrv4 I__4818 (
            .O(N__28614),
            .I(\ALU.madd_29_0 ));
    LocalMux I__4817 (
            .O(N__28611),
            .I(\ALU.madd_29_0 ));
    InMux I__4816 (
            .O(N__28606),
            .I(N__28603));
    LocalMux I__4815 (
            .O(N__28603),
            .I(N__28600));
    Odrv4 I__4814 (
            .O(N__28600),
            .I(\ALU.madd_18 ));
    InMux I__4813 (
            .O(N__28597),
            .I(N__28594));
    LocalMux I__4812 (
            .O(N__28594),
            .I(N__28590));
    InMux I__4811 (
            .O(N__28593),
            .I(N__28587));
    Odrv4 I__4810 (
            .O(N__28590),
            .I(\ALU.madd_34 ));
    LocalMux I__4809 (
            .O(N__28587),
            .I(\ALU.madd_34 ));
    CascadeMux I__4808 (
            .O(N__28582),
            .I(\ALU.madd_39_cascade_ ));
    InMux I__4807 (
            .O(N__28579),
            .I(N__28576));
    LocalMux I__4806 (
            .O(N__28576),
            .I(\ALU.madd_39 ));
    CascadeMux I__4805 (
            .O(N__28573),
            .I(\ALU.madd_23_cascade_ ));
    InMux I__4804 (
            .O(N__28570),
            .I(N__28567));
    LocalMux I__4803 (
            .O(N__28567),
            .I(N__28564));
    Span4Mux_v I__4802 (
            .O(N__28564),
            .I(N__28560));
    InMux I__4801 (
            .O(N__28563),
            .I(N__28557));
    Odrv4 I__4800 (
            .O(N__28560),
            .I(\ALU.madd_28 ));
    LocalMux I__4799 (
            .O(N__28557),
            .I(\ALU.madd_28 ));
    CascadeMux I__4798 (
            .O(N__28552),
            .I(N__28549));
    InMux I__4797 (
            .O(N__28549),
            .I(N__28546));
    LocalMux I__4796 (
            .O(N__28546),
            .I(N__28543));
    Span4Mux_v I__4795 (
            .O(N__28543),
            .I(N__28540));
    Odrv4 I__4794 (
            .O(N__28540),
            .I(\ALU.madd_axb_4_l_fx ));
    InMux I__4793 (
            .O(N__28537),
            .I(N__28528));
    InMux I__4792 (
            .O(N__28536),
            .I(N__28528));
    InMux I__4791 (
            .O(N__28535),
            .I(N__28528));
    LocalMux I__4790 (
            .O(N__28528),
            .I(\ALU.madd_8 ));
    InMux I__4789 (
            .O(N__28525),
            .I(N__28519));
    InMux I__4788 (
            .O(N__28524),
            .I(N__28519));
    LocalMux I__4787 (
            .O(N__28519),
            .I(N__28516));
    Span4Mux_h I__4786 (
            .O(N__28516),
            .I(N__28513));
    Odrv4 I__4785 (
            .O(N__28513),
            .I(\ALU.madd_19 ));
    InMux I__4784 (
            .O(N__28510),
            .I(N__28507));
    LocalMux I__4783 (
            .O(N__28507),
            .I(N__28504));
    Odrv4 I__4782 (
            .O(N__28504),
            .I(TXbuffer_RNO_1Z0Z_5));
    InMux I__4781 (
            .O(N__28501),
            .I(N__28498));
    LocalMux I__4780 (
            .O(N__28498),
            .I(N__28495));
    Odrv4 I__4779 (
            .O(N__28495),
            .I(TXbuffer_RNO_0Z0Z_5));
    InMux I__4778 (
            .O(N__28492),
            .I(N__28489));
    LocalMux I__4777 (
            .O(N__28489),
            .I(N__28486));
    Odrv4 I__4776 (
            .O(N__28486),
            .I(TXbuffer_18_15_ns_1_5));
    CascadeMux I__4775 (
            .O(N__28483),
            .I(\ALU.a2_b_1_cascade_ ));
    InMux I__4774 (
            .O(N__28480),
            .I(N__28477));
    LocalMux I__4773 (
            .O(N__28477),
            .I(\ALU.a1_b_2 ));
    InMux I__4772 (
            .O(N__28474),
            .I(N__28471));
    LocalMux I__4771 (
            .O(N__28471),
            .I(\ALU.a2_b_1 ));
    CascadeMux I__4770 (
            .O(N__28468),
            .I(\ALU.a1_b_2_cascade_ ));
    InMux I__4769 (
            .O(N__28465),
            .I(N__28462));
    LocalMux I__4768 (
            .O(N__28462),
            .I(\ALU.r0_12_prm_3_12_s0_sf ));
    InMux I__4767 (
            .O(N__28459),
            .I(N__28456));
    LocalMux I__4766 (
            .O(N__28456),
            .I(N__28453));
    Odrv12 I__4765 (
            .O(N__28453),
            .I(\ALU.mult_12 ));
    InMux I__4764 (
            .O(N__28450),
            .I(\ALU.r0_12_s0_12 ));
    CascadeMux I__4763 (
            .O(N__28447),
            .I(N__28443));
    InMux I__4762 (
            .O(N__28446),
            .I(N__28437));
    InMux I__4761 (
            .O(N__28443),
            .I(N__28434));
    InMux I__4760 (
            .O(N__28442),
            .I(N__28431));
    InMux I__4759 (
            .O(N__28441),
            .I(N__28428));
    InMux I__4758 (
            .O(N__28440),
            .I(N__28424));
    LocalMux I__4757 (
            .O(N__28437),
            .I(N__28420));
    LocalMux I__4756 (
            .O(N__28434),
            .I(N__28415));
    LocalMux I__4755 (
            .O(N__28431),
            .I(N__28415));
    LocalMux I__4754 (
            .O(N__28428),
            .I(N__28412));
    InMux I__4753 (
            .O(N__28427),
            .I(N__28409));
    LocalMux I__4752 (
            .O(N__28424),
            .I(N__28406));
    InMux I__4751 (
            .O(N__28423),
            .I(N__28403));
    Span4Mux_h I__4750 (
            .O(N__28420),
            .I(N__28397));
    Span4Mux_v I__4749 (
            .O(N__28415),
            .I(N__28397));
    Span4Mux_h I__4748 (
            .O(N__28412),
            .I(N__28392));
    LocalMux I__4747 (
            .O(N__28409),
            .I(N__28392));
    Span4Mux_v I__4746 (
            .O(N__28406),
            .I(N__28387));
    LocalMux I__4745 (
            .O(N__28403),
            .I(N__28387));
    InMux I__4744 (
            .O(N__28402),
            .I(N__28384));
    Odrv4 I__4743 (
            .O(N__28397),
            .I(\ALU.r0_12_12 ));
    Odrv4 I__4742 (
            .O(N__28392),
            .I(\ALU.r0_12_12 ));
    Odrv4 I__4741 (
            .O(N__28387),
            .I(\ALU.r0_12_12 ));
    LocalMux I__4740 (
            .O(N__28384),
            .I(\ALU.r0_12_12 ));
    InMux I__4739 (
            .O(N__28375),
            .I(N__28370));
    InMux I__4738 (
            .O(N__28374),
            .I(N__28367));
    InMux I__4737 (
            .O(N__28373),
            .I(N__28364));
    LocalMux I__4736 (
            .O(N__28370),
            .I(N__28361));
    LocalMux I__4735 (
            .O(N__28367),
            .I(N__28358));
    LocalMux I__4734 (
            .O(N__28364),
            .I(N__28355));
    Span4Mux_h I__4733 (
            .O(N__28361),
            .I(N__28352));
    Span4Mux_h I__4732 (
            .O(N__28358),
            .I(N__28349));
    Span4Mux_h I__4731 (
            .O(N__28355),
            .I(N__28346));
    Span4Mux_v I__4730 (
            .O(N__28352),
            .I(N__28343));
    Odrv4 I__4729 (
            .O(N__28349),
            .I(r0_12));
    Odrv4 I__4728 (
            .O(N__28346),
            .I(r0_12));
    Odrv4 I__4727 (
            .O(N__28343),
            .I(r0_12));
    CascadeMux I__4726 (
            .O(N__28336),
            .I(N__28333));
    InMux I__4725 (
            .O(N__28333),
            .I(N__28330));
    LocalMux I__4724 (
            .O(N__28330),
            .I(\ALU.r0_12_prm_3_14_s0_sf ));
    InMux I__4723 (
            .O(N__28327),
            .I(N__28324));
    LocalMux I__4722 (
            .O(N__28324),
            .I(N__28321));
    Span4Mux_v I__4721 (
            .O(N__28321),
            .I(N__28318));
    Odrv4 I__4720 (
            .O(N__28318),
            .I(\ALU.mult_14 ));
    InMux I__4719 (
            .O(N__28315),
            .I(\ALU.r0_12_s0_14 ));
    InMux I__4718 (
            .O(N__28312),
            .I(N__28305));
    InMux I__4717 (
            .O(N__28311),
            .I(N__28302));
    InMux I__4716 (
            .O(N__28310),
            .I(N__28299));
    InMux I__4715 (
            .O(N__28309),
            .I(N__28296));
    InMux I__4714 (
            .O(N__28308),
            .I(N__28290));
    LocalMux I__4713 (
            .O(N__28305),
            .I(N__28287));
    LocalMux I__4712 (
            .O(N__28302),
            .I(N__28284));
    LocalMux I__4711 (
            .O(N__28299),
            .I(N__28279));
    LocalMux I__4710 (
            .O(N__28296),
            .I(N__28279));
    InMux I__4709 (
            .O(N__28295),
            .I(N__28276));
    InMux I__4708 (
            .O(N__28294),
            .I(N__28273));
    InMux I__4707 (
            .O(N__28293),
            .I(N__28270));
    LocalMux I__4706 (
            .O(N__28290),
            .I(N__28267));
    Span4Mux_h I__4705 (
            .O(N__28287),
            .I(N__28264));
    Span4Mux_h I__4704 (
            .O(N__28284),
            .I(N__28259));
    Span4Mux_v I__4703 (
            .O(N__28279),
            .I(N__28259));
    LocalMux I__4702 (
            .O(N__28276),
            .I(\ALU.r0_12_14 ));
    LocalMux I__4701 (
            .O(N__28273),
            .I(\ALU.r0_12_14 ));
    LocalMux I__4700 (
            .O(N__28270),
            .I(\ALU.r0_12_14 ));
    Odrv4 I__4699 (
            .O(N__28267),
            .I(\ALU.r0_12_14 ));
    Odrv4 I__4698 (
            .O(N__28264),
            .I(\ALU.r0_12_14 ));
    Odrv4 I__4697 (
            .O(N__28259),
            .I(\ALU.r0_12_14 ));
    InMux I__4696 (
            .O(N__28246),
            .I(N__28242));
    InMux I__4695 (
            .O(N__28245),
            .I(N__28239));
    LocalMux I__4694 (
            .O(N__28242),
            .I(N__28235));
    LocalMux I__4693 (
            .O(N__28239),
            .I(N__28232));
    CascadeMux I__4692 (
            .O(N__28238),
            .I(N__28229));
    Span4Mux_h I__4691 (
            .O(N__28235),
            .I(N__28226));
    Span4Mux_h I__4690 (
            .O(N__28232),
            .I(N__28223));
    InMux I__4689 (
            .O(N__28229),
            .I(N__28220));
    Odrv4 I__4688 (
            .O(N__28226),
            .I(r1_14));
    Odrv4 I__4687 (
            .O(N__28223),
            .I(r1_14));
    LocalMux I__4686 (
            .O(N__28220),
            .I(r1_14));
    InMux I__4685 (
            .O(N__28213),
            .I(N__28210));
    LocalMux I__4684 (
            .O(N__28210),
            .I(\ALU.r0_12_prm_3_10_s0_sf ));
    InMux I__4683 (
            .O(N__28207),
            .I(N__28204));
    LocalMux I__4682 (
            .O(N__28204),
            .I(N__28201));
    Span4Mux_v I__4681 (
            .O(N__28201),
            .I(N__28198));
    Odrv4 I__4680 (
            .O(N__28198),
            .I(\ALU.mult_10 ));
    InMux I__4679 (
            .O(N__28195),
            .I(\ALU.r0_12_s0_10 ));
    InMux I__4678 (
            .O(N__28192),
            .I(N__28186));
    InMux I__4677 (
            .O(N__28191),
            .I(N__28183));
    InMux I__4676 (
            .O(N__28190),
            .I(N__28180));
    InMux I__4675 (
            .O(N__28189),
            .I(N__28177));
    LocalMux I__4674 (
            .O(N__28186),
            .I(N__28173));
    LocalMux I__4673 (
            .O(N__28183),
            .I(N__28170));
    LocalMux I__4672 (
            .O(N__28180),
            .I(N__28167));
    LocalMux I__4671 (
            .O(N__28177),
            .I(N__28164));
    InMux I__4670 (
            .O(N__28176),
            .I(N__28161));
    Span4Mux_h I__4669 (
            .O(N__28173),
            .I(N__28153));
    Span4Mux_h I__4668 (
            .O(N__28170),
            .I(N__28153));
    Span4Mux_v I__4667 (
            .O(N__28167),
            .I(N__28148));
    Span4Mux_v I__4666 (
            .O(N__28164),
            .I(N__28148));
    LocalMux I__4665 (
            .O(N__28161),
            .I(N__28145));
    InMux I__4664 (
            .O(N__28160),
            .I(N__28142));
    InMux I__4663 (
            .O(N__28159),
            .I(N__28139));
    InMux I__4662 (
            .O(N__28158),
            .I(N__28136));
    Odrv4 I__4661 (
            .O(N__28153),
            .I(\ALU.r0_12_10 ));
    Odrv4 I__4660 (
            .O(N__28148),
            .I(\ALU.r0_12_10 ));
    Odrv4 I__4659 (
            .O(N__28145),
            .I(\ALU.r0_12_10 ));
    LocalMux I__4658 (
            .O(N__28142),
            .I(\ALU.r0_12_10 ));
    LocalMux I__4657 (
            .O(N__28139),
            .I(\ALU.r0_12_10 ));
    LocalMux I__4656 (
            .O(N__28136),
            .I(\ALU.r0_12_10 ));
    InMux I__4655 (
            .O(N__28123),
            .I(N__28118));
    InMux I__4654 (
            .O(N__28122),
            .I(N__28115));
    InMux I__4653 (
            .O(N__28121),
            .I(N__28112));
    LocalMux I__4652 (
            .O(N__28118),
            .I(N__28109));
    LocalMux I__4651 (
            .O(N__28115),
            .I(N__28106));
    LocalMux I__4650 (
            .O(N__28112),
            .I(N__28103));
    Span4Mux_h I__4649 (
            .O(N__28109),
            .I(N__28100));
    Span12Mux_s6_h I__4648 (
            .O(N__28106),
            .I(N__28097));
    Odrv4 I__4647 (
            .O(N__28103),
            .I(r0_10));
    Odrv4 I__4646 (
            .O(N__28100),
            .I(r0_10));
    Odrv12 I__4645 (
            .O(N__28097),
            .I(r0_10));
    InMux I__4644 (
            .O(N__28090),
            .I(N__28083));
    InMux I__4643 (
            .O(N__28089),
            .I(N__28083));
    InMux I__4642 (
            .O(N__28088),
            .I(N__28080));
    LocalMux I__4641 (
            .O(N__28083),
            .I(N__28077));
    LocalMux I__4640 (
            .O(N__28080),
            .I(N__28074));
    Span4Mux_s3_h I__4639 (
            .O(N__28077),
            .I(N__28071));
    Span4Mux_v I__4638 (
            .O(N__28074),
            .I(N__28068));
    Span4Mux_h I__4637 (
            .O(N__28071),
            .I(N__28065));
    Odrv4 I__4636 (
            .O(N__28068),
            .I(r7_2));
    Odrv4 I__4635 (
            .O(N__28065),
            .I(r7_2));
    InMux I__4634 (
            .O(N__28060),
            .I(N__28056));
    InMux I__4633 (
            .O(N__28059),
            .I(N__28053));
    LocalMux I__4632 (
            .O(N__28056),
            .I(N__28050));
    LocalMux I__4631 (
            .O(N__28053),
            .I(N__28047));
    Span4Mux_v I__4630 (
            .O(N__28050),
            .I(N__28041));
    Span4Mux_v I__4629 (
            .O(N__28047),
            .I(N__28041));
    InMux I__4628 (
            .O(N__28046),
            .I(N__28038));
    Span4Mux_h I__4627 (
            .O(N__28041),
            .I(N__28035));
    LocalMux I__4626 (
            .O(N__28038),
            .I(N__28032));
    Odrv4 I__4625 (
            .O(N__28035),
            .I(r7_3));
    Odrv4 I__4624 (
            .O(N__28032),
            .I(r7_3));
    InMux I__4623 (
            .O(N__28027),
            .I(N__28024));
    LocalMux I__4622 (
            .O(N__28024),
            .I(N__28021));
    Span4Mux_v I__4621 (
            .O(N__28021),
            .I(N__28018));
    Span4Mux_h I__4620 (
            .O(N__28018),
            .I(N__28013));
    InMux I__4619 (
            .O(N__28017),
            .I(N__28008));
    InMux I__4618 (
            .O(N__28016),
            .I(N__28008));
    Span4Mux_v I__4617 (
            .O(N__28013),
            .I(N__28003));
    LocalMux I__4616 (
            .O(N__28008),
            .I(N__28003));
    Odrv4 I__4615 (
            .O(N__28003),
            .I(r7_4));
    CascadeMux I__4614 (
            .O(N__28000),
            .I(TXbuffer_18_10_ns_1_1_cascade_));
    InMux I__4613 (
            .O(N__27997),
            .I(N__27994));
    LocalMux I__4612 (
            .O(N__27994),
            .I(N__27991));
    Sp12to4 I__4611 (
            .O(N__27991),
            .I(N__27988));
    Span12Mux_v I__4610 (
            .O(N__27988),
            .I(N__27985));
    Odrv12 I__4609 (
            .O(N__27985),
            .I(TXbuffer_18_15_ns_1_1));
    CascadeMux I__4608 (
            .O(N__27982),
            .I(TXbuffer_RNO_0Z0Z_1_cascade_));
    InMux I__4607 (
            .O(N__27979),
            .I(N__27976));
    LocalMux I__4606 (
            .O(N__27976),
            .I(TXbuffer_RNO_1Z0Z_1));
    CascadeMux I__4605 (
            .O(N__27973),
            .I(N__27969));
    InMux I__4604 (
            .O(N__27972),
            .I(N__27966));
    InMux I__4603 (
            .O(N__27969),
            .I(N__27963));
    LocalMux I__4602 (
            .O(N__27966),
            .I(N__27959));
    LocalMux I__4601 (
            .O(N__27963),
            .I(N__27956));
    CascadeMux I__4600 (
            .O(N__27962),
            .I(N__27953));
    Span4Mux_h I__4599 (
            .O(N__27959),
            .I(N__27950));
    Span4Mux_h I__4598 (
            .O(N__27956),
            .I(N__27947));
    InMux I__4597 (
            .O(N__27953),
            .I(N__27944));
    Odrv4 I__4596 (
            .O(N__27950),
            .I(r1_10));
    Odrv4 I__4595 (
            .O(N__27947),
            .I(r1_10));
    LocalMux I__4594 (
            .O(N__27944),
            .I(r1_10));
    InMux I__4593 (
            .O(N__27937),
            .I(N__27933));
    InMux I__4592 (
            .O(N__27936),
            .I(N__27929));
    LocalMux I__4591 (
            .O(N__27933),
            .I(N__27926));
    InMux I__4590 (
            .O(N__27932),
            .I(N__27923));
    LocalMux I__4589 (
            .O(N__27929),
            .I(N__27920));
    Span4Mux_h I__4588 (
            .O(N__27926),
            .I(N__27917));
    LocalMux I__4587 (
            .O(N__27923),
            .I(N__27914));
    Span4Mux_v I__4586 (
            .O(N__27920),
            .I(N__27911));
    Span4Mux_v I__4585 (
            .O(N__27917),
            .I(N__27908));
    Span4Mux_h I__4584 (
            .O(N__27914),
            .I(N__27905));
    Odrv4 I__4583 (
            .O(N__27911),
            .I(r5_10));
    Odrv4 I__4582 (
            .O(N__27908),
            .I(r5_10));
    Odrv4 I__4581 (
            .O(N__27905),
            .I(r5_10));
    CascadeMux I__4580 (
            .O(N__27898),
            .I(TXbuffer_18_10_ns_1_2_cascade_));
    InMux I__4579 (
            .O(N__27895),
            .I(N__27892));
    LocalMux I__4578 (
            .O(N__27892),
            .I(N__27889));
    Span4Mux_v I__4577 (
            .O(N__27889),
            .I(N__27886));
    Odrv4 I__4576 (
            .O(N__27886),
            .I(TXbuffer_RNO_0Z0Z_2));
    InMux I__4575 (
            .O(N__27883),
            .I(N__27879));
    InMux I__4574 (
            .O(N__27882),
            .I(N__27875));
    LocalMux I__4573 (
            .O(N__27879),
            .I(N__27872));
    InMux I__4572 (
            .O(N__27878),
            .I(N__27869));
    LocalMux I__4571 (
            .O(N__27875),
            .I(N__27866));
    Span4Mux_h I__4570 (
            .O(N__27872),
            .I(N__27863));
    LocalMux I__4569 (
            .O(N__27869),
            .I(N__27860));
    Span4Mux_h I__4568 (
            .O(N__27866),
            .I(N__27853));
    Span4Mux_v I__4567 (
            .O(N__27863),
            .I(N__27853));
    Span4Mux_h I__4566 (
            .O(N__27860),
            .I(N__27853));
    Odrv4 I__4565 (
            .O(N__27853),
            .I(r7_6));
    InMux I__4564 (
            .O(N__27850),
            .I(N__27847));
    LocalMux I__4563 (
            .O(N__27847),
            .I(N__27844));
    Span4Mux_v I__4562 (
            .O(N__27844),
            .I(N__27839));
    InMux I__4561 (
            .O(N__27843),
            .I(N__27834));
    InMux I__4560 (
            .O(N__27842),
            .I(N__27834));
    Sp12to4 I__4559 (
            .O(N__27839),
            .I(N__27829));
    LocalMux I__4558 (
            .O(N__27834),
            .I(N__27829));
    Odrv12 I__4557 (
            .O(N__27829),
            .I(r7_7));
    InMux I__4556 (
            .O(N__27826),
            .I(N__27821));
    InMux I__4555 (
            .O(N__27825),
            .I(N__27816));
    InMux I__4554 (
            .O(N__27824),
            .I(N__27816));
    LocalMux I__4553 (
            .O(N__27821),
            .I(N__27813));
    LocalMux I__4552 (
            .O(N__27816),
            .I(N__27810));
    Span12Mux_s6_h I__4551 (
            .O(N__27813),
            .I(N__27807));
    Span4Mux_h I__4550 (
            .O(N__27810),
            .I(N__27804));
    Odrv12 I__4549 (
            .O(N__27807),
            .I(r7_8));
    Odrv4 I__4548 (
            .O(N__27804),
            .I(r7_8));
    CascadeMux I__4547 (
            .O(N__27799),
            .I(N__27796));
    InMux I__4546 (
            .O(N__27796),
            .I(N__27792));
    InMux I__4545 (
            .O(N__27795),
            .I(N__27789));
    LocalMux I__4544 (
            .O(N__27792),
            .I(N__27786));
    LocalMux I__4543 (
            .O(N__27789),
            .I(N__27782));
    Span4Mux_v I__4542 (
            .O(N__27786),
            .I(N__27779));
    InMux I__4541 (
            .O(N__27785),
            .I(N__27776));
    Span4Mux_h I__4540 (
            .O(N__27782),
            .I(N__27773));
    Span4Mux_s3_h I__4539 (
            .O(N__27779),
            .I(N__27770));
    LocalMux I__4538 (
            .O(N__27776),
            .I(r7_9));
    Odrv4 I__4537 (
            .O(N__27773),
            .I(r7_9));
    Odrv4 I__4536 (
            .O(N__27770),
            .I(r7_9));
    InMux I__4535 (
            .O(N__27763),
            .I(N__27760));
    LocalMux I__4534 (
            .O(N__27760),
            .I(\ALU.r4_RNIJJH11Z0Z_0 ));
    CascadeMux I__4533 (
            .O(N__27757),
            .I(\ALU.r0_RNIBROOZ0Z_0_cascade_ ));
    InMux I__4532 (
            .O(N__27754),
            .I(N__27745));
    InMux I__4531 (
            .O(N__27753),
            .I(N__27745));
    InMux I__4530 (
            .O(N__27752),
            .I(N__27742));
    InMux I__4529 (
            .O(N__27751),
            .I(N__27735));
    InMux I__4528 (
            .O(N__27750),
            .I(N__27735));
    LocalMux I__4527 (
            .O(N__27745),
            .I(N__27729));
    LocalMux I__4526 (
            .O(N__27742),
            .I(N__27729));
    InMux I__4525 (
            .O(N__27741),
            .I(N__27724));
    InMux I__4524 (
            .O(N__27740),
            .I(N__27724));
    LocalMux I__4523 (
            .O(N__27735),
            .I(N__27721));
    InMux I__4522 (
            .O(N__27734),
            .I(N__27717));
    Span4Mux_v I__4521 (
            .O(N__27729),
            .I(N__27710));
    LocalMux I__4520 (
            .O(N__27724),
            .I(N__27710));
    Span4Mux_h I__4519 (
            .O(N__27721),
            .I(N__27710));
    InMux I__4518 (
            .O(N__27720),
            .I(N__27707));
    LocalMux I__4517 (
            .O(N__27717),
            .I(a_fastZ0Z_1));
    Odrv4 I__4516 (
            .O(N__27710),
            .I(a_fastZ0Z_1));
    LocalMux I__4515 (
            .O(N__27707),
            .I(a_fastZ0Z_1));
    InMux I__4514 (
            .O(N__27700),
            .I(N__27697));
    LocalMux I__4513 (
            .O(N__27697),
            .I(N__27694));
    Span4Mux_s2_v I__4512 (
            .O(N__27694),
            .I(N__27691));
    Span4Mux_v I__4511 (
            .O(N__27691),
            .I(N__27688));
    Odrv4 I__4510 (
            .O(N__27688),
            .I(\ALU.a_7_ns_1_0 ));
    InMux I__4509 (
            .O(N__27685),
            .I(N__27682));
    LocalMux I__4508 (
            .O(N__27682),
            .I(N__27677));
    InMux I__4507 (
            .O(N__27681),
            .I(N__27672));
    InMux I__4506 (
            .O(N__27680),
            .I(N__27672));
    Span4Mux_h I__4505 (
            .O(N__27677),
            .I(N__27669));
    LocalMux I__4504 (
            .O(N__27672),
            .I(N__27666));
    Span4Mux_v I__4503 (
            .O(N__27669),
            .I(N__27661));
    Span4Mux_v I__4502 (
            .O(N__27666),
            .I(N__27661));
    Odrv4 I__4501 (
            .O(N__27661),
            .I(r4_0));
    CascadeMux I__4500 (
            .O(N__27658),
            .I(TXbuffer_18_3_ns_1_0_cascade_));
    InMux I__4499 (
            .O(N__27655),
            .I(N__27652));
    LocalMux I__4498 (
            .O(N__27652),
            .I(N__27649));
    Span4Mux_v I__4497 (
            .O(N__27649),
            .I(N__27646));
    Span4Mux_h I__4496 (
            .O(N__27646),
            .I(N__27643));
    Odrv4 I__4495 (
            .O(N__27643),
            .I(TXbuffer_RNO_5Z0Z_0));
    CascadeMux I__4494 (
            .O(N__27640),
            .I(TXbuffer_18_10_ns_1_0_cascade_));
    CascadeMux I__4493 (
            .O(N__27637),
            .I(N__27634));
    InMux I__4492 (
            .O(N__27634),
            .I(N__27631));
    LocalMux I__4491 (
            .O(N__27631),
            .I(N__27626));
    InMux I__4490 (
            .O(N__27630),
            .I(N__27621));
    InMux I__4489 (
            .O(N__27629),
            .I(N__27621));
    Span4Mux_v I__4488 (
            .O(N__27626),
            .I(N__27618));
    LocalMux I__4487 (
            .O(N__27621),
            .I(N__27615));
    Span4Mux_v I__4486 (
            .O(N__27618),
            .I(N__27610));
    Span4Mux_v I__4485 (
            .O(N__27615),
            .I(N__27610));
    Odrv4 I__4484 (
            .O(N__27610),
            .I(r5_0));
    InMux I__4483 (
            .O(N__27607),
            .I(N__27604));
    LocalMux I__4482 (
            .O(N__27604),
            .I(N__27601));
    Span4Mux_s2_h I__4481 (
            .O(N__27601),
            .I(N__27598));
    Span4Mux_h I__4480 (
            .O(N__27598),
            .I(N__27595));
    Sp12to4 I__4479 (
            .O(N__27595),
            .I(N__27592));
    Odrv12 I__4478 (
            .O(N__27592),
            .I(TXbuffer_RNO_0Z0Z_0));
    InMux I__4477 (
            .O(N__27589),
            .I(N__27585));
    CascadeMux I__4476 (
            .O(N__27588),
            .I(N__27582));
    LocalMux I__4475 (
            .O(N__27585),
            .I(N__27578));
    InMux I__4474 (
            .O(N__27582),
            .I(N__27575));
    InMux I__4473 (
            .O(N__27581),
            .I(N__27572));
    Span4Mux_v I__4472 (
            .O(N__27578),
            .I(N__27567));
    LocalMux I__4471 (
            .O(N__27575),
            .I(N__27567));
    LocalMux I__4470 (
            .O(N__27572),
            .I(N__27562));
    Span4Mux_h I__4469 (
            .O(N__27567),
            .I(N__27562));
    Odrv4 I__4468 (
            .O(N__27562),
            .I(r3_9));
    CascadeMux I__4467 (
            .O(N__27559),
            .I(N__27556));
    InMux I__4466 (
            .O(N__27556),
            .I(N__27553));
    LocalMux I__4465 (
            .O(N__27553),
            .I(TXbuffer_18_13_ns_1_1));
    CascadeMux I__4464 (
            .O(N__27550),
            .I(N__27547));
    InMux I__4463 (
            .O(N__27547),
            .I(N__27544));
    LocalMux I__4462 (
            .O(N__27544),
            .I(N__27541));
    Odrv12 I__4461 (
            .O(N__27541),
            .I(\ALU.madd_cry_9_ma ));
    InMux I__4460 (
            .O(N__27538),
            .I(\ALU.madd_cry_8 ));
    CascadeMux I__4459 (
            .O(N__27535),
            .I(N__27531));
    InMux I__4458 (
            .O(N__27534),
            .I(N__27528));
    InMux I__4457 (
            .O(N__27531),
            .I(N__27525));
    LocalMux I__4456 (
            .O(N__27528),
            .I(N__27522));
    LocalMux I__4455 (
            .O(N__27525),
            .I(N__27519));
    Span12Mux_h I__4454 (
            .O(N__27522),
            .I(N__27516));
    Span12Mux_v I__4453 (
            .O(N__27519),
            .I(N__27513));
    Odrv12 I__4452 (
            .O(N__27516),
            .I(\ALU.madd_axb_10 ));
    Odrv12 I__4451 (
            .O(N__27513),
            .I(\ALU.madd_axb_10 ));
    CascadeMux I__4450 (
            .O(N__27508),
            .I(N__27505));
    InMux I__4449 (
            .O(N__27505),
            .I(N__27502));
    LocalMux I__4448 (
            .O(N__27502),
            .I(N__27499));
    Span4Mux_v I__4447 (
            .O(N__27499),
            .I(N__27496));
    Span4Mux_h I__4446 (
            .O(N__27496),
            .I(N__27493));
    Odrv4 I__4445 (
            .O(N__27493),
            .I(\ALU.madd_cry_9_THRU_CO ));
    InMux I__4444 (
            .O(N__27490),
            .I(\ALU.madd_cry_9 ));
    InMux I__4443 (
            .O(N__27487),
            .I(N__27484));
    LocalMux I__4442 (
            .O(N__27484),
            .I(N__27481));
    Span4Mux_v I__4441 (
            .O(N__27481),
            .I(N__27477));
    InMux I__4440 (
            .O(N__27480),
            .I(N__27474));
    Span4Mux_h I__4439 (
            .O(N__27477),
            .I(N__27471));
    LocalMux I__4438 (
            .O(N__27474),
            .I(N__27468));
    Span4Mux_v I__4437 (
            .O(N__27471),
            .I(N__27465));
    Odrv4 I__4436 (
            .O(N__27468),
            .I(\ALU.g0_13 ));
    Odrv4 I__4435 (
            .O(N__27465),
            .I(\ALU.g0_13 ));
    CascadeMux I__4434 (
            .O(N__27460),
            .I(N__27457));
    InMux I__4433 (
            .O(N__27457),
            .I(N__27454));
    LocalMux I__4432 (
            .O(N__27454),
            .I(N__27451));
    Span4Mux_v I__4431 (
            .O(N__27451),
            .I(N__27448));
    Odrv4 I__4430 (
            .O(N__27448),
            .I(\ALU.madd_axb_11_l_fx ));
    InMux I__4429 (
            .O(N__27445),
            .I(\ALU.madd_cry_10 ));
    InMux I__4428 (
            .O(N__27442),
            .I(N__27439));
    LocalMux I__4427 (
            .O(N__27439),
            .I(N__27436));
    Span4Mux_v I__4426 (
            .O(N__27436),
            .I(N__27433));
    Odrv4 I__4425 (
            .O(N__27433),
            .I(\ALU.madd_cry_12_ma ));
    CascadeMux I__4424 (
            .O(N__27430),
            .I(N__27427));
    InMux I__4423 (
            .O(N__27427),
            .I(N__27424));
    LocalMux I__4422 (
            .O(N__27424),
            .I(N__27421));
    Span4Mux_v I__4421 (
            .O(N__27421),
            .I(N__27418));
    Span4Mux_h I__4420 (
            .O(N__27418),
            .I(N__27415));
    Odrv4 I__4419 (
            .O(N__27415),
            .I(\ALU.madd_axb_12_l_ofx ));
    InMux I__4418 (
            .O(N__27412),
            .I(N__27409));
    LocalMux I__4417 (
            .O(N__27409),
            .I(N__27406));
    Span4Mux_v I__4416 (
            .O(N__27406),
            .I(N__27403));
    Span4Mux_v I__4415 (
            .O(N__27403),
            .I(N__27400));
    Odrv4 I__4414 (
            .O(N__27400),
            .I(\ALU.mult_13 ));
    InMux I__4413 (
            .O(N__27397),
            .I(\ALU.madd_cry_11 ));
    InMux I__4412 (
            .O(N__27394),
            .I(N__27391));
    LocalMux I__4411 (
            .O(N__27391),
            .I(N__27388));
    Span4Mux_h I__4410 (
            .O(N__27388),
            .I(N__27385));
    Span4Mux_s3_h I__4409 (
            .O(N__27385),
            .I(N__27382));
    Odrv4 I__4408 (
            .O(N__27382),
            .I(\ALU.madd_axb_13_l_ofx ));
    CascadeMux I__4407 (
            .O(N__27379),
            .I(N__27376));
    InMux I__4406 (
            .O(N__27376),
            .I(N__27373));
    LocalMux I__4405 (
            .O(N__27373),
            .I(N__27370));
    Span4Mux_h I__4404 (
            .O(N__27370),
            .I(N__27367));
    Odrv4 I__4403 (
            .O(N__27367),
            .I(\ALU.madd_cry_13_ma ));
    InMux I__4402 (
            .O(N__27364),
            .I(\ALU.madd_cry_12 ));
    InMux I__4401 (
            .O(N__27361),
            .I(\ALU.madd_cry_13 ));
    CascadeMux I__4400 (
            .O(N__27358),
            .I(N__27355));
    InMux I__4399 (
            .O(N__27355),
            .I(N__27352));
    LocalMux I__4398 (
            .O(N__27352),
            .I(N__27349));
    Span12Mux_v I__4397 (
            .O(N__27349),
            .I(N__27346));
    Odrv12 I__4396 (
            .O(N__27346),
            .I(\ALU.madd_cry_13_THRU_CO ));
    InMux I__4395 (
            .O(N__27343),
            .I(N__27338));
    InMux I__4394 (
            .O(N__27342),
            .I(N__27333));
    InMux I__4393 (
            .O(N__27341),
            .I(N__27333));
    LocalMux I__4392 (
            .O(N__27338),
            .I(\ALU.a13_b_1 ));
    LocalMux I__4391 (
            .O(N__27333),
            .I(\ALU.a13_b_1 ));
    InMux I__4390 (
            .O(N__27328),
            .I(N__27325));
    LocalMux I__4389 (
            .O(N__27325),
            .I(N__27322));
    Span4Mux_v I__4388 (
            .O(N__27322),
            .I(N__27319));
    Odrv4 I__4387 (
            .O(N__27319),
            .I(\ALU.madd_373_0 ));
    CascadeMux I__4386 (
            .O(N__27316),
            .I(N__27313));
    InMux I__4385 (
            .O(N__27313),
            .I(N__27310));
    LocalMux I__4384 (
            .O(N__27310),
            .I(\ALU.madd_368_0 ));
    InMux I__4383 (
            .O(N__27307),
            .I(N__27303));
    InMux I__4382 (
            .O(N__27306),
            .I(N__27300));
    LocalMux I__4381 (
            .O(N__27303),
            .I(N__27297));
    LocalMux I__4380 (
            .O(N__27300),
            .I(N__27294));
    Span4Mux_v I__4379 (
            .O(N__27297),
            .I(N__27291));
    Span4Mux_v I__4378 (
            .O(N__27294),
            .I(N__27288));
    Span4Mux_h I__4377 (
            .O(N__27291),
            .I(N__27285));
    Odrv4 I__4376 (
            .O(N__27288),
            .I(\ALU.a9_b_5 ));
    Odrv4 I__4375 (
            .O(N__27285),
            .I(\ALU.a9_b_5 ));
    InMux I__4374 (
            .O(N__27280),
            .I(N__27274));
    InMux I__4373 (
            .O(N__27279),
            .I(N__27274));
    LocalMux I__4372 (
            .O(N__27274),
            .I(N__27271));
    Odrv12 I__4371 (
            .O(N__27271),
            .I(\ALU.madd_398_0 ));
    InMux I__4370 (
            .O(N__27268),
            .I(\ALU.madd_cry_0 ));
    InMux I__4369 (
            .O(N__27265),
            .I(\ALU.madd_cry_1 ));
    InMux I__4368 (
            .O(N__27262),
            .I(\ALU.madd_cry_2 ));
    InMux I__4367 (
            .O(N__27259),
            .I(\ALU.madd_cry_3 ));
    CascadeMux I__4366 (
            .O(N__27256),
            .I(N__27253));
    InMux I__4365 (
            .O(N__27253),
            .I(N__27250));
    LocalMux I__4364 (
            .O(N__27250),
            .I(N__27247));
    Odrv12 I__4363 (
            .O(N__27247),
            .I(\ALU.madd_axb_5_l_fx ));
    InMux I__4362 (
            .O(N__27244),
            .I(\ALU.madd_cry_4 ));
    InMux I__4361 (
            .O(N__27241),
            .I(N__27238));
    LocalMux I__4360 (
            .O(N__27238),
            .I(N__27235));
    Span4Mux_v I__4359 (
            .O(N__27235),
            .I(N__27232));
    Odrv4 I__4358 (
            .O(N__27232),
            .I(\ALU.madd_axb_6_l_ofx ));
    InMux I__4357 (
            .O(N__27229),
            .I(\ALU.madd_cry_5 ));
    InMux I__4356 (
            .O(N__27226),
            .I(\ALU.madd_cry_6 ));
    CascadeMux I__4355 (
            .O(N__27223),
            .I(N__27220));
    InMux I__4354 (
            .O(N__27220),
            .I(N__27216));
    InMux I__4353 (
            .O(N__27219),
            .I(N__27213));
    LocalMux I__4352 (
            .O(N__27216),
            .I(N__27210));
    LocalMux I__4351 (
            .O(N__27213),
            .I(N__27207));
    Span4Mux_v I__4350 (
            .O(N__27210),
            .I(N__27204));
    Span4Mux_v I__4349 (
            .O(N__27207),
            .I(N__27201));
    Odrv4 I__4348 (
            .O(N__27204),
            .I(\ALU.madd_165 ));
    Odrv4 I__4347 (
            .O(N__27201),
            .I(\ALU.madd_165 ));
    CascadeMux I__4346 (
            .O(N__27196),
            .I(N__27193));
    InMux I__4345 (
            .O(N__27193),
            .I(N__27190));
    LocalMux I__4344 (
            .O(N__27190),
            .I(N__27187));
    Span4Mux_v I__4343 (
            .O(N__27187),
            .I(N__27184));
    Odrv4 I__4342 (
            .O(N__27184),
            .I(\ALU.madd_axb_8_l_fx ));
    InMux I__4341 (
            .O(N__27181),
            .I(bfn_7_7_0_));
    InMux I__4340 (
            .O(N__27178),
            .I(N__27175));
    LocalMux I__4339 (
            .O(N__27175),
            .I(N__27172));
    Span4Mux_v I__4338 (
            .O(N__27172),
            .I(N__27169));
    Odrv4 I__4337 (
            .O(N__27169),
            .I(\ALU.madd_axb_9_l_ofx ));
    CascadeMux I__4336 (
            .O(N__27166),
            .I(\ALU.a5_b_1_cascade_ ));
    InMux I__4335 (
            .O(N__27163),
            .I(N__27160));
    LocalMux I__4334 (
            .O(N__27160),
            .I(N__27157));
    Odrv4 I__4333 (
            .O(N__27157),
            .I(\ALU.madd_50 ));
    InMux I__4332 (
            .O(N__27154),
            .I(N__27150));
    InMux I__4331 (
            .O(N__27153),
            .I(N__27147));
    LocalMux I__4330 (
            .O(N__27150),
            .I(\ALU.madd_55 ));
    LocalMux I__4329 (
            .O(N__27147),
            .I(\ALU.madd_55 ));
    CascadeMux I__4328 (
            .O(N__27142),
            .I(\ALU.madd_50_cascade_ ));
    InMux I__4327 (
            .O(N__27139),
            .I(N__27135));
    InMux I__4326 (
            .O(N__27138),
            .I(N__27132));
    LocalMux I__4325 (
            .O(N__27135),
            .I(\ALU.madd_73 ));
    LocalMux I__4324 (
            .O(N__27132),
            .I(\ALU.madd_73 ));
    CascadeMux I__4323 (
            .O(N__27127),
            .I(N__27124));
    InMux I__4322 (
            .O(N__27124),
            .I(N__27118));
    InMux I__4321 (
            .O(N__27123),
            .I(N__27118));
    LocalMux I__4320 (
            .O(N__27118),
            .I(\ALU.madd_83 ));
    InMux I__4319 (
            .O(N__27115),
            .I(N__27112));
    LocalMux I__4318 (
            .O(N__27112),
            .I(N__27109));
    Span4Mux_v I__4317 (
            .O(N__27109),
            .I(N__27106));
    Span4Mux_h I__4316 (
            .O(N__27106),
            .I(N__27103));
    Sp12to4 I__4315 (
            .O(N__27103),
            .I(N__27100));
    Odrv12 I__4314 (
            .O(N__27100),
            .I(TXbuffer_RNO_1Z0Z_2));
    InMux I__4313 (
            .O(N__27097),
            .I(N__27094));
    LocalMux I__4312 (
            .O(N__27094),
            .I(N__27091));
    Span4Mux_v I__4311 (
            .O(N__27091),
            .I(N__27088));
    Span4Mux_h I__4310 (
            .O(N__27088),
            .I(N__27085));
    Odrv4 I__4309 (
            .O(N__27085),
            .I(TXbuffer_18_15_ns_1_2));
    InMux I__4308 (
            .O(N__27082),
            .I(N__27079));
    LocalMux I__4307 (
            .O(N__27079),
            .I(N__27076));
    Sp12to4 I__4306 (
            .O(N__27076),
            .I(N__27071));
    InMux I__4305 (
            .O(N__27075),
            .I(N__27068));
    InMux I__4304 (
            .O(N__27074),
            .I(N__27065));
    Span12Mux_v I__4303 (
            .O(N__27071),
            .I(N__27062));
    LocalMux I__4302 (
            .O(N__27068),
            .I(clkdivZ0Z_1));
    LocalMux I__4301 (
            .O(N__27065),
            .I(clkdivZ0Z_1));
    Odrv12 I__4300 (
            .O(N__27062),
            .I(clkdivZ0Z_1));
    InMux I__4299 (
            .O(N__27055),
            .I(N__27052));
    LocalMux I__4298 (
            .O(N__27052),
            .I(N__27047));
    InMux I__4297 (
            .O(N__27051),
            .I(N__27044));
    InMux I__4296 (
            .O(N__27050),
            .I(N__27041));
    Span12Mux_v I__4295 (
            .O(N__27047),
            .I(N__27038));
    LocalMux I__4294 (
            .O(N__27044),
            .I(clkdivZ0Z_2));
    LocalMux I__4293 (
            .O(N__27041),
            .I(clkdivZ0Z_2));
    Odrv12 I__4292 (
            .O(N__27038),
            .I(clkdivZ0Z_2));
    CascadeMux I__4291 (
            .O(N__27031),
            .I(N__27028));
    InMux I__4290 (
            .O(N__27028),
            .I(N__27025));
    LocalMux I__4289 (
            .O(N__27025),
            .I(N__27022));
    Span4Mux_v I__4288 (
            .O(N__27022),
            .I(N__27019));
    Span4Mux_h I__4287 (
            .O(N__27019),
            .I(N__27016));
    IoSpan4Mux I__4286 (
            .O(N__27016),
            .I(N__27012));
    CascadeMux I__4285 (
            .O(N__27015),
            .I(N__27009));
    IoSpan4Mux I__4284 (
            .O(N__27012),
            .I(N__27005));
    InMux I__4283 (
            .O(N__27009),
            .I(N__27002));
    InMux I__4282 (
            .O(N__27008),
            .I(N__26999));
    Span4Mux_s1_h I__4281 (
            .O(N__27005),
            .I(N__26996));
    LocalMux I__4280 (
            .O(N__27002),
            .I(clkdivZ0Z_3));
    LocalMux I__4279 (
            .O(N__26999),
            .I(clkdivZ0Z_3));
    Odrv4 I__4278 (
            .O(N__26996),
            .I(clkdivZ0Z_3));
    InMux I__4277 (
            .O(N__26989),
            .I(N__26986));
    LocalMux I__4276 (
            .O(N__26986),
            .I(N__26983));
    Span4Mux_h I__4275 (
            .O(N__26983),
            .I(N__26980));
    Span4Mux_h I__4274 (
            .O(N__26980),
            .I(N__26977));
    Span4Mux_v I__4273 (
            .O(N__26977),
            .I(N__26972));
    InMux I__4272 (
            .O(N__26976),
            .I(N__26969));
    InMux I__4271 (
            .O(N__26975),
            .I(N__26966));
    Span4Mux_v I__4270 (
            .O(N__26972),
            .I(N__26963));
    LocalMux I__4269 (
            .O(N__26969),
            .I(clkdivZ0Z_0));
    LocalMux I__4268 (
            .O(N__26966),
            .I(clkdivZ0Z_0));
    Odrv4 I__4267 (
            .O(N__26963),
            .I(clkdivZ0Z_0));
    IoInMux I__4266 (
            .O(N__26956),
            .I(N__26953));
    LocalMux I__4265 (
            .O(N__26953),
            .I(N__26950));
    Span12Mux_s11_h I__4264 (
            .O(N__26950),
            .I(N__26947));
    Span12Mux_v I__4263 (
            .O(N__26947),
            .I(N__26944));
    Odrv12 I__4262 (
            .O(N__26944),
            .I(params5));
    CascadeMux I__4261 (
            .O(N__26941),
            .I(\ALU.madd_axb_3_cascade_ ));
    InMux I__4260 (
            .O(N__26938),
            .I(N__26932));
    InMux I__4259 (
            .O(N__26937),
            .I(N__26932));
    LocalMux I__4258 (
            .O(N__26932),
            .I(N__26929));
    Odrv12 I__4257 (
            .O(N__26929),
            .I(\ALU.madd_14 ));
    InMux I__4256 (
            .O(N__26926),
            .I(N__26923));
    LocalMux I__4255 (
            .O(N__26923),
            .I(N__26920));
    Odrv4 I__4254 (
            .O(N__26920),
            .I(\ALU.madd_cry_0_ma ));
    CascadeMux I__4253 (
            .O(N__26917),
            .I(N__26914));
    InMux I__4252 (
            .O(N__26914),
            .I(N__26911));
    LocalMux I__4251 (
            .O(N__26911),
            .I(N__26908));
    Odrv4 I__4250 (
            .O(N__26908),
            .I(\ALU.madd_axb_0_l_ofx ));
    CascadeMux I__4249 (
            .O(N__26905),
            .I(\ALU.madd_73_0_cascade_ ));
    InMux I__4248 (
            .O(N__26902),
            .I(N__26899));
    LocalMux I__4247 (
            .O(N__26899),
            .I(N__26896));
    Odrv4 I__4246 (
            .O(N__26896),
            .I(\ALU.a1_b_5 ));
    CascadeMux I__4245 (
            .O(N__26893),
            .I(N__26890));
    InMux I__4244 (
            .O(N__26890),
            .I(N__26886));
    InMux I__4243 (
            .O(N__26889),
            .I(N__26883));
    LocalMux I__4242 (
            .O(N__26886),
            .I(\ALU.a2_b_4 ));
    LocalMux I__4241 (
            .O(N__26883),
            .I(\ALU.a2_b_4 ));
    CascadeMux I__4240 (
            .O(N__26878),
            .I(\ALU.a1_b_5_cascade_ ));
    InMux I__4239 (
            .O(N__26875),
            .I(N__26871));
    InMux I__4238 (
            .O(N__26874),
            .I(N__26868));
    LocalMux I__4237 (
            .O(N__26871),
            .I(N__26865));
    LocalMux I__4236 (
            .O(N__26868),
            .I(b_fastZ0Z_1));
    Odrv4 I__4235 (
            .O(N__26865),
            .I(b_fastZ0Z_1));
    CascadeMux I__4234 (
            .O(N__26860),
            .I(N__26853));
    CascadeMux I__4233 (
            .O(N__26859),
            .I(N__26847));
    CascadeMux I__4232 (
            .O(N__26858),
            .I(N__26841));
    InMux I__4231 (
            .O(N__26857),
            .I(N__26834));
    InMux I__4230 (
            .O(N__26856),
            .I(N__26834));
    InMux I__4229 (
            .O(N__26853),
            .I(N__26834));
    InMux I__4228 (
            .O(N__26852),
            .I(N__26829));
    InMux I__4227 (
            .O(N__26851),
            .I(N__26824));
    InMux I__4226 (
            .O(N__26850),
            .I(N__26821));
    InMux I__4225 (
            .O(N__26847),
            .I(N__26816));
    InMux I__4224 (
            .O(N__26846),
            .I(N__26816));
    InMux I__4223 (
            .O(N__26845),
            .I(N__26809));
    InMux I__4222 (
            .O(N__26844),
            .I(N__26809));
    InMux I__4221 (
            .O(N__26841),
            .I(N__26809));
    LocalMux I__4220 (
            .O(N__26834),
            .I(N__26806));
    InMux I__4219 (
            .O(N__26833),
            .I(N__26803));
    InMux I__4218 (
            .O(N__26832),
            .I(N__26800));
    LocalMux I__4217 (
            .O(N__26829),
            .I(N__26794));
    InMux I__4216 (
            .O(N__26828),
            .I(N__26791));
    InMux I__4215 (
            .O(N__26827),
            .I(N__26788));
    LocalMux I__4214 (
            .O(N__26824),
            .I(N__26783));
    LocalMux I__4213 (
            .O(N__26821),
            .I(N__26783));
    LocalMux I__4212 (
            .O(N__26816),
            .I(N__26780));
    LocalMux I__4211 (
            .O(N__26809),
            .I(N__26775));
    Span4Mux_v I__4210 (
            .O(N__26806),
            .I(N__26775));
    LocalMux I__4209 (
            .O(N__26803),
            .I(N__26772));
    LocalMux I__4208 (
            .O(N__26800),
            .I(N__26769));
    InMux I__4207 (
            .O(N__26799),
            .I(N__26762));
    InMux I__4206 (
            .O(N__26798),
            .I(N__26762));
    InMux I__4205 (
            .O(N__26797),
            .I(N__26762));
    Sp12to4 I__4204 (
            .O(N__26794),
            .I(N__26757));
    LocalMux I__4203 (
            .O(N__26791),
            .I(N__26757));
    LocalMux I__4202 (
            .O(N__26788),
            .I(N__26752));
    Span4Mux_v I__4201 (
            .O(N__26783),
            .I(N__26752));
    Span4Mux_h I__4200 (
            .O(N__26780),
            .I(N__26747));
    Span4Mux_h I__4199 (
            .O(N__26775),
            .I(N__26747));
    Odrv4 I__4198 (
            .O(N__26772),
            .I(b_2_repZ0Z2));
    Odrv12 I__4197 (
            .O(N__26769),
            .I(b_2_repZ0Z2));
    LocalMux I__4196 (
            .O(N__26762),
            .I(b_2_repZ0Z2));
    Odrv12 I__4195 (
            .O(N__26757),
            .I(b_2_repZ0Z2));
    Odrv4 I__4194 (
            .O(N__26752),
            .I(b_2_repZ0Z2));
    Odrv4 I__4193 (
            .O(N__26747),
            .I(b_2_repZ0Z2));
    CascadeMux I__4192 (
            .O(N__26734),
            .I(\ALU.r4_RNIMTDQZ0Z_1_cascade_ ));
    InMux I__4191 (
            .O(N__26731),
            .I(N__26728));
    LocalMux I__4190 (
            .O(N__26728),
            .I(\ALU.b_7_ns_1_1 ));
    InMux I__4189 (
            .O(N__26725),
            .I(N__26719));
    InMux I__4188 (
            .O(N__26724),
            .I(N__26719));
    LocalMux I__4187 (
            .O(N__26719),
            .I(N__26715));
    InMux I__4186 (
            .O(N__26718),
            .I(N__26712));
    Odrv4 I__4185 (
            .O(N__26715),
            .I(\ALU.madd_46 ));
    LocalMux I__4184 (
            .O(N__26712),
            .I(\ALU.madd_46 ));
    CascadeMux I__4183 (
            .O(N__26707),
            .I(N__26704));
    InMux I__4182 (
            .O(N__26704),
            .I(N__26701));
    LocalMux I__4181 (
            .O(N__26701),
            .I(N__26698));
    Odrv4 I__4180 (
            .O(N__26698),
            .I(\ALU.a5_b_1 ));
    CascadeMux I__4179 (
            .O(N__26695),
            .I(\ALU.madd_18_cascade_ ));
    CascadeMux I__4178 (
            .O(N__26692),
            .I(\ALU.madd_43_cascade_ ));
    InMux I__4177 (
            .O(N__26689),
            .I(N__26683));
    InMux I__4176 (
            .O(N__26688),
            .I(N__26683));
    LocalMux I__4175 (
            .O(N__26683),
            .I(\ALU.a2_b_3 ));
    InMux I__4174 (
            .O(N__26680),
            .I(N__26676));
    InMux I__4173 (
            .O(N__26679),
            .I(N__26673));
    LocalMux I__4172 (
            .O(N__26676),
            .I(\ALU.madd_332 ));
    LocalMux I__4171 (
            .O(N__26673),
            .I(\ALU.madd_332 ));
    InMux I__4170 (
            .O(N__26668),
            .I(N__26665));
    LocalMux I__4169 (
            .O(N__26665),
            .I(\ALU.madd_94 ));
    InMux I__4168 (
            .O(N__26662),
            .I(N__26658));
    InMux I__4167 (
            .O(N__26661),
            .I(N__26655));
    LocalMux I__4166 (
            .O(N__26658),
            .I(\ALU.madd_33 ));
    LocalMux I__4165 (
            .O(N__26655),
            .I(\ALU.madd_33 ));
    InMux I__4164 (
            .O(N__26650),
            .I(N__26647));
    LocalMux I__4163 (
            .O(N__26647),
            .I(\ALU.madd_38 ));
    InMux I__4162 (
            .O(N__26644),
            .I(N__26640));
    InMux I__4161 (
            .O(N__26643),
            .I(N__26637));
    LocalMux I__4160 (
            .O(N__26640),
            .I(\ALU.a0_b_6 ));
    LocalMux I__4159 (
            .O(N__26637),
            .I(\ALU.a0_b_6 ));
    CascadeMux I__4158 (
            .O(N__26632),
            .I(N__26629));
    InMux I__4157 (
            .O(N__26629),
            .I(N__26625));
    InMux I__4156 (
            .O(N__26628),
            .I(N__26622));
    LocalMux I__4155 (
            .O(N__26625),
            .I(N__26619));
    LocalMux I__4154 (
            .O(N__26622),
            .I(\ALU.madd_51 ));
    Odrv4 I__4153 (
            .O(N__26619),
            .I(\ALU.madd_51 ));
    CascadeMux I__4152 (
            .O(N__26614),
            .I(\ALU.madd_51_cascade_ ));
    InMux I__4151 (
            .O(N__26611),
            .I(N__26607));
    InMux I__4150 (
            .O(N__26610),
            .I(N__26604));
    LocalMux I__4149 (
            .O(N__26607),
            .I(\ALU.madd_43 ));
    LocalMux I__4148 (
            .O(N__26604),
            .I(\ALU.madd_43 ));
    InMux I__4147 (
            .O(N__26599),
            .I(N__26593));
    InMux I__4146 (
            .O(N__26598),
            .I(N__26593));
    LocalMux I__4145 (
            .O(N__26593),
            .I(\ALU.madd_331 ));
    InMux I__4144 (
            .O(N__26590),
            .I(N__26584));
    InMux I__4143 (
            .O(N__26589),
            .I(N__26584));
    LocalMux I__4142 (
            .O(N__26584),
            .I(\ALU.a1_b_4 ));
    InMux I__4141 (
            .O(N__26581),
            .I(N__26578));
    LocalMux I__4140 (
            .O(N__26578),
            .I(\ALU.madd_87 ));
    InMux I__4139 (
            .O(N__26575),
            .I(N__26572));
    LocalMux I__4138 (
            .O(N__26572),
            .I(N__26569));
    Span4Mux_s1_v I__4137 (
            .O(N__26569),
            .I(N__26565));
    InMux I__4136 (
            .O(N__26568),
            .I(N__26562));
    Odrv4 I__4135 (
            .O(N__26565),
            .I(\ALU.madd_110 ));
    LocalMux I__4134 (
            .O(N__26562),
            .I(\ALU.madd_110 ));
    InMux I__4133 (
            .O(N__26557),
            .I(N__26553));
    InMux I__4132 (
            .O(N__26556),
            .I(N__26550));
    LocalMux I__4131 (
            .O(N__26553),
            .I(\ALU.madd_115 ));
    LocalMux I__4130 (
            .O(N__26550),
            .I(\ALU.madd_115 ));
    InMux I__4129 (
            .O(N__26545),
            .I(N__26539));
    InMux I__4128 (
            .O(N__26544),
            .I(N__26539));
    LocalMux I__4127 (
            .O(N__26539),
            .I(\ALU.madd_124 ));
    CascadeMux I__4126 (
            .O(N__26536),
            .I(\ALU.madd_124_cascade_ ));
    InMux I__4125 (
            .O(N__26533),
            .I(N__26528));
    InMux I__4124 (
            .O(N__26532),
            .I(N__26523));
    InMux I__4123 (
            .O(N__26531),
            .I(N__26523));
    LocalMux I__4122 (
            .O(N__26528),
            .I(N__26518));
    LocalMux I__4121 (
            .O(N__26523),
            .I(N__26518));
    Odrv12 I__4120 (
            .O(N__26518),
            .I(\ALU.madd_160 ));
    CascadeMux I__4119 (
            .O(N__26515),
            .I(N__26509));
    InMux I__4118 (
            .O(N__26514),
            .I(N__26505));
    InMux I__4117 (
            .O(N__26513),
            .I(N__26501));
    InMux I__4116 (
            .O(N__26512),
            .I(N__26498));
    InMux I__4115 (
            .O(N__26509),
            .I(N__26495));
    InMux I__4114 (
            .O(N__26508),
            .I(N__26492));
    LocalMux I__4113 (
            .O(N__26505),
            .I(N__26489));
    InMux I__4112 (
            .O(N__26504),
            .I(N__26486));
    LocalMux I__4111 (
            .O(N__26501),
            .I(N__26483));
    LocalMux I__4110 (
            .O(N__26498),
            .I(N__26480));
    LocalMux I__4109 (
            .O(N__26495),
            .I(N__26477));
    LocalMux I__4108 (
            .O(N__26492),
            .I(N__26474));
    Span12Mux_s7_v I__4107 (
            .O(N__26489),
            .I(N__26471));
    LocalMux I__4106 (
            .O(N__26486),
            .I(N__26466));
    Span4Mux_v I__4105 (
            .O(N__26483),
            .I(N__26466));
    Span12Mux_s7_v I__4104 (
            .O(N__26480),
            .I(N__26463));
    Span12Mux_s4_h I__4103 (
            .O(N__26477),
            .I(N__26458));
    Span12Mux_s1_v I__4102 (
            .O(N__26474),
            .I(N__26458));
    Odrv12 I__4101 (
            .O(N__26471),
            .I(\ALU.r6_RNIE0JB2Z0Z_6 ));
    Odrv4 I__4100 (
            .O(N__26466),
            .I(\ALU.r6_RNIE0JB2Z0Z_6 ));
    Odrv12 I__4099 (
            .O(N__26463),
            .I(\ALU.r6_RNIE0JB2Z0Z_6 ));
    Odrv12 I__4098 (
            .O(N__26458),
            .I(\ALU.r6_RNIE0JB2Z0Z_6 ));
    InMux I__4097 (
            .O(N__26449),
            .I(N__26444));
    InMux I__4096 (
            .O(N__26448),
            .I(N__26441));
    InMux I__4095 (
            .O(N__26447),
            .I(N__26438));
    LocalMux I__4094 (
            .O(N__26444),
            .I(N__26432));
    LocalMux I__4093 (
            .O(N__26441),
            .I(N__26429));
    LocalMux I__4092 (
            .O(N__26438),
            .I(N__26426));
    InMux I__4091 (
            .O(N__26437),
            .I(N__26423));
    InMux I__4090 (
            .O(N__26436),
            .I(N__26420));
    InMux I__4089 (
            .O(N__26435),
            .I(N__26417));
    Span4Mux_v I__4088 (
            .O(N__26432),
            .I(N__26414));
    Span4Mux_h I__4087 (
            .O(N__26429),
            .I(N__26411));
    Span4Mux_h I__4086 (
            .O(N__26426),
            .I(N__26406));
    LocalMux I__4085 (
            .O(N__26423),
            .I(N__26406));
    LocalMux I__4084 (
            .O(N__26420),
            .I(N__26403));
    LocalMux I__4083 (
            .O(N__26417),
            .I(N__26400));
    Span4Mux_h I__4082 (
            .O(N__26414),
            .I(N__26395));
    Span4Mux_v I__4081 (
            .O(N__26411),
            .I(N__26395));
    Span4Mux_v I__4080 (
            .O(N__26406),
            .I(N__26390));
    Span4Mux_v I__4079 (
            .O(N__26403),
            .I(N__26390));
    Odrv12 I__4078 (
            .O(N__26400),
            .I(\ALU.r4_RNI68Q22Z0Z_6 ));
    Odrv4 I__4077 (
            .O(N__26395),
            .I(\ALU.r4_RNI68Q22Z0Z_6 ));
    Odrv4 I__4076 (
            .O(N__26390),
            .I(\ALU.r4_RNI68Q22Z0Z_6 ));
    CascadeMux I__4075 (
            .O(N__26383),
            .I(N__26380));
    InMux I__4074 (
            .O(N__26380),
            .I(N__26377));
    LocalMux I__4073 (
            .O(N__26377),
            .I(\ALU.a3_b_1 ));
    CascadeMux I__4072 (
            .O(N__26374),
            .I(\ALU.a3_b_1_cascade_ ));
    CascadeMux I__4071 (
            .O(N__26371),
            .I(N__26368));
    InMux I__4070 (
            .O(N__26368),
            .I(N__26365));
    LocalMux I__4069 (
            .O(N__26365),
            .I(N__26362));
    Odrv12 I__4068 (
            .O(N__26362),
            .I(\ALU.r5_RNIK81F5Z0Z_13 ));
    InMux I__4067 (
            .O(N__26359),
            .I(N__26356));
    LocalMux I__4066 (
            .O(N__26356),
            .I(N__26353));
    Odrv4 I__4065 (
            .O(N__26353),
            .I(\ALU.r0_12_prm_5_13_s0_c_RNOZ0 ));
    CascadeMux I__4064 (
            .O(N__26350),
            .I(N__26347));
    InMux I__4063 (
            .O(N__26347),
            .I(N__26344));
    LocalMux I__4062 (
            .O(N__26344),
            .I(N__26341));
    Span4Mux_v I__4061 (
            .O(N__26341),
            .I(N__26338));
    Odrv4 I__4060 (
            .O(N__26338),
            .I(\ALU.r0_12_prm_6_13_s0_c_RNOZ0 ));
    CascadeMux I__4059 (
            .O(N__26335),
            .I(N__26332));
    InMux I__4058 (
            .O(N__26332),
            .I(N__26329));
    LocalMux I__4057 (
            .O(N__26329),
            .I(N__26326));
    Odrv4 I__4056 (
            .O(N__26326),
            .I(\ALU.r0_12_prm_7_13_s0_c_RNOZ0 ));
    CascadeMux I__4055 (
            .O(N__26323),
            .I(N__26320));
    InMux I__4054 (
            .O(N__26320),
            .I(N__26316));
    InMux I__4053 (
            .O(N__26319),
            .I(N__26313));
    LocalMux I__4052 (
            .O(N__26316),
            .I(N__26310));
    LocalMux I__4051 (
            .O(N__26313),
            .I(\ALU.madd_334 ));
    Odrv12 I__4050 (
            .O(N__26310),
            .I(\ALU.madd_334 ));
    InMux I__4049 (
            .O(N__26305),
            .I(N__26301));
    InMux I__4048 (
            .O(N__26304),
            .I(N__26298));
    LocalMux I__4047 (
            .O(N__26301),
            .I(N__26295));
    LocalMux I__4046 (
            .O(N__26298),
            .I(\ALU.madd_333 ));
    Odrv12 I__4045 (
            .O(N__26295),
            .I(\ALU.madd_333 ));
    InMux I__4044 (
            .O(N__26290),
            .I(N__26287));
    LocalMux I__4043 (
            .O(N__26287),
            .I(\ALU.r0_12_prm_3_13_s0_sf ));
    InMux I__4042 (
            .O(N__26284),
            .I(\ALU.r0_12_s0_13 ));
    InMux I__4041 (
            .O(N__26281),
            .I(N__26274));
    InMux I__4040 (
            .O(N__26280),
            .I(N__26271));
    InMux I__4039 (
            .O(N__26279),
            .I(N__26268));
    InMux I__4038 (
            .O(N__26278),
            .I(N__26265));
    InMux I__4037 (
            .O(N__26277),
            .I(N__26262));
    LocalMux I__4036 (
            .O(N__26274),
            .I(N__26258));
    LocalMux I__4035 (
            .O(N__26271),
            .I(N__26255));
    LocalMux I__4034 (
            .O(N__26268),
            .I(N__26252));
    LocalMux I__4033 (
            .O(N__26265),
            .I(N__26249));
    LocalMux I__4032 (
            .O(N__26262),
            .I(N__26246));
    InMux I__4031 (
            .O(N__26261),
            .I(N__26243));
    Span4Mux_h I__4030 (
            .O(N__26258),
            .I(N__26232));
    Span4Mux_v I__4029 (
            .O(N__26255),
            .I(N__26232));
    Span4Mux_h I__4028 (
            .O(N__26252),
            .I(N__26232));
    Span4Mux_v I__4027 (
            .O(N__26249),
            .I(N__26232));
    Span4Mux_h I__4026 (
            .O(N__26246),
            .I(N__26227));
    LocalMux I__4025 (
            .O(N__26243),
            .I(N__26227));
    InMux I__4024 (
            .O(N__26242),
            .I(N__26224));
    InMux I__4023 (
            .O(N__26241),
            .I(N__26221));
    Odrv4 I__4022 (
            .O(N__26232),
            .I(\ALU.r0_12_13 ));
    Odrv4 I__4021 (
            .O(N__26227),
            .I(\ALU.r0_12_13 ));
    LocalMux I__4020 (
            .O(N__26224),
            .I(\ALU.r0_12_13 ));
    LocalMux I__4019 (
            .O(N__26221),
            .I(\ALU.r0_12_13 ));
    InMux I__4018 (
            .O(N__26212),
            .I(N__26208));
    InMux I__4017 (
            .O(N__26211),
            .I(N__26205));
    LocalMux I__4016 (
            .O(N__26208),
            .I(N__26202));
    LocalMux I__4015 (
            .O(N__26205),
            .I(N__26199));
    Span4Mux_h I__4014 (
            .O(N__26202),
            .I(N__26193));
    Span4Mux_h I__4013 (
            .O(N__26199),
            .I(N__26193));
    InMux I__4012 (
            .O(N__26198),
            .I(N__26190));
    Odrv4 I__4011 (
            .O(N__26193),
            .I(r0_13));
    LocalMux I__4010 (
            .O(N__26190),
            .I(r0_13));
    InMux I__4009 (
            .O(N__26185),
            .I(N__26180));
    InMux I__4008 (
            .O(N__26184),
            .I(N__26177));
    InMux I__4007 (
            .O(N__26183),
            .I(N__26173));
    LocalMux I__4006 (
            .O(N__26180),
            .I(N__26169));
    LocalMux I__4005 (
            .O(N__26177),
            .I(N__26166));
    InMux I__4004 (
            .O(N__26176),
            .I(N__26163));
    LocalMux I__4003 (
            .O(N__26173),
            .I(N__26160));
    InMux I__4002 (
            .O(N__26172),
            .I(N__26157));
    Span4Mux_v I__4001 (
            .O(N__26169),
            .I(N__26149));
    Span4Mux_v I__4000 (
            .O(N__26166),
            .I(N__26149));
    LocalMux I__3999 (
            .O(N__26163),
            .I(N__26146));
    Span4Mux_h I__3998 (
            .O(N__26160),
            .I(N__26141));
    LocalMux I__3997 (
            .O(N__26157),
            .I(N__26141));
    InMux I__3996 (
            .O(N__26156),
            .I(N__26138));
    InMux I__3995 (
            .O(N__26155),
            .I(N__26135));
    InMux I__3994 (
            .O(N__26154),
            .I(N__26132));
    Odrv4 I__3993 (
            .O(N__26149),
            .I(\ALU.r0_12_11 ));
    Odrv4 I__3992 (
            .O(N__26146),
            .I(\ALU.r0_12_11 ));
    Odrv4 I__3991 (
            .O(N__26141),
            .I(\ALU.r0_12_11 ));
    LocalMux I__3990 (
            .O(N__26138),
            .I(\ALU.r0_12_11 ));
    LocalMux I__3989 (
            .O(N__26135),
            .I(\ALU.r0_12_11 ));
    LocalMux I__3988 (
            .O(N__26132),
            .I(\ALU.r0_12_11 ));
    InMux I__3987 (
            .O(N__26119),
            .I(N__26115));
    InMux I__3986 (
            .O(N__26118),
            .I(N__26112));
    LocalMux I__3985 (
            .O(N__26115),
            .I(N__26108));
    LocalMux I__3984 (
            .O(N__26112),
            .I(N__26105));
    InMux I__3983 (
            .O(N__26111),
            .I(N__26102));
    Span4Mux_v I__3982 (
            .O(N__26108),
            .I(N__26099));
    Span4Mux_v I__3981 (
            .O(N__26105),
            .I(N__26094));
    LocalMux I__3980 (
            .O(N__26102),
            .I(N__26094));
    Span4Mux_h I__3979 (
            .O(N__26099),
            .I(N__26091));
    Span4Mux_h I__3978 (
            .O(N__26094),
            .I(N__26088));
    Odrv4 I__3977 (
            .O(N__26091),
            .I(r5_11));
    Odrv4 I__3976 (
            .O(N__26088),
            .I(r5_11));
    InMux I__3975 (
            .O(N__26083),
            .I(N__26080));
    LocalMux I__3974 (
            .O(N__26080),
            .I(N__26075));
    InMux I__3973 (
            .O(N__26079),
            .I(N__26072));
    InMux I__3972 (
            .O(N__26078),
            .I(N__26069));
    Span4Mux_s1_h I__3971 (
            .O(N__26075),
            .I(N__26064));
    LocalMux I__3970 (
            .O(N__26072),
            .I(N__26064));
    LocalMux I__3969 (
            .O(N__26069),
            .I(N__26061));
    Span4Mux_h I__3968 (
            .O(N__26064),
            .I(N__26058));
    Span4Mux_h I__3967 (
            .O(N__26061),
            .I(N__26055));
    Odrv4 I__3966 (
            .O(N__26058),
            .I(r5_12));
    Odrv4 I__3965 (
            .O(N__26055),
            .I(r5_12));
    InMux I__3964 (
            .O(N__26050),
            .I(N__26046));
    InMux I__3963 (
            .O(N__26049),
            .I(N__26042));
    LocalMux I__3962 (
            .O(N__26046),
            .I(N__26039));
    InMux I__3961 (
            .O(N__26045),
            .I(N__26036));
    LocalMux I__3960 (
            .O(N__26042),
            .I(N__26029));
    Span4Mux_h I__3959 (
            .O(N__26039),
            .I(N__26029));
    LocalMux I__3958 (
            .O(N__26036),
            .I(N__26029));
    Odrv4 I__3957 (
            .O(N__26029),
            .I(r5_13));
    InMux I__3956 (
            .O(N__26026),
            .I(N__26022));
    InMux I__3955 (
            .O(N__26025),
            .I(N__26018));
    LocalMux I__3954 (
            .O(N__26022),
            .I(N__26015));
    InMux I__3953 (
            .O(N__26021),
            .I(N__26012));
    LocalMux I__3952 (
            .O(N__26018),
            .I(N__26009));
    Span4Mux_s3_h I__3951 (
            .O(N__26015),
            .I(N__26006));
    LocalMux I__3950 (
            .O(N__26012),
            .I(N__26003));
    Span4Mux_v I__3949 (
            .O(N__26009),
            .I(N__25998));
    Span4Mux_v I__3948 (
            .O(N__26006),
            .I(N__25998));
    Odrv4 I__3947 (
            .O(N__26003),
            .I(r5_14));
    Odrv4 I__3946 (
            .O(N__25998),
            .I(r5_14));
    CascadeMux I__3945 (
            .O(N__25993),
            .I(N__25990));
    InMux I__3944 (
            .O(N__25990),
            .I(N__25983));
    InMux I__3943 (
            .O(N__25989),
            .I(N__25980));
    InMux I__3942 (
            .O(N__25988),
            .I(N__25977));
    InMux I__3941 (
            .O(N__25987),
            .I(N__25973));
    CascadeMux I__3940 (
            .O(N__25986),
            .I(N__25969));
    LocalMux I__3939 (
            .O(N__25983),
            .I(N__25965));
    LocalMux I__3938 (
            .O(N__25980),
            .I(N__25962));
    LocalMux I__3937 (
            .O(N__25977),
            .I(N__25959));
    InMux I__3936 (
            .O(N__25976),
            .I(N__25956));
    LocalMux I__3935 (
            .O(N__25973),
            .I(N__25953));
    InMux I__3934 (
            .O(N__25972),
            .I(N__25950));
    InMux I__3933 (
            .O(N__25969),
            .I(N__25947));
    InMux I__3932 (
            .O(N__25968),
            .I(N__25944));
    Odrv4 I__3931 (
            .O(N__25965),
            .I(\ALU.r0_12_15 ));
    Odrv4 I__3930 (
            .O(N__25962),
            .I(\ALU.r0_12_15 ));
    Odrv4 I__3929 (
            .O(N__25959),
            .I(\ALU.r0_12_15 ));
    LocalMux I__3928 (
            .O(N__25956),
            .I(\ALU.r0_12_15 ));
    Odrv4 I__3927 (
            .O(N__25953),
            .I(\ALU.r0_12_15 ));
    LocalMux I__3926 (
            .O(N__25950),
            .I(\ALU.r0_12_15 ));
    LocalMux I__3925 (
            .O(N__25947),
            .I(\ALU.r0_12_15 ));
    LocalMux I__3924 (
            .O(N__25944),
            .I(\ALU.r0_12_15 ));
    InMux I__3923 (
            .O(N__25927),
            .I(N__25923));
    InMux I__3922 (
            .O(N__25926),
            .I(N__25919));
    LocalMux I__3921 (
            .O(N__25923),
            .I(N__25916));
    InMux I__3920 (
            .O(N__25922),
            .I(N__25913));
    LocalMux I__3919 (
            .O(N__25919),
            .I(N__25910));
    Span4Mux_h I__3918 (
            .O(N__25916),
            .I(N__25907));
    LocalMux I__3917 (
            .O(N__25913),
            .I(N__25904));
    Span12Mux_s5_h I__3916 (
            .O(N__25910),
            .I(N__25901));
    Span4Mux_v I__3915 (
            .O(N__25907),
            .I(N__25898));
    Odrv4 I__3914 (
            .O(N__25904),
            .I(r5_5));
    Odrv12 I__3913 (
            .O(N__25901),
            .I(r5_5));
    Odrv4 I__3912 (
            .O(N__25898),
            .I(r5_5));
    CascadeMux I__3911 (
            .O(N__25891),
            .I(\ALU.a_3_ns_1_14_cascade_ ));
    InMux I__3910 (
            .O(N__25888),
            .I(N__25884));
    InMux I__3909 (
            .O(N__25887),
            .I(N__25881));
    LocalMux I__3908 (
            .O(N__25884),
            .I(N__25877));
    LocalMux I__3907 (
            .O(N__25881),
            .I(N__25874));
    InMux I__3906 (
            .O(N__25880),
            .I(N__25871));
    Span4Mux_v I__3905 (
            .O(N__25877),
            .I(N__25866));
    Span4Mux_v I__3904 (
            .O(N__25874),
            .I(N__25866));
    LocalMux I__3903 (
            .O(N__25871),
            .I(r4_14));
    Odrv4 I__3902 (
            .O(N__25866),
            .I(r4_14));
    InMux I__3901 (
            .O(N__25861),
            .I(N__25858));
    LocalMux I__3900 (
            .O(N__25858),
            .I(N__25854));
    InMux I__3899 (
            .O(N__25857),
            .I(N__25851));
    Span4Mux_v I__3898 (
            .O(N__25854),
            .I(N__25848));
    LocalMux I__3897 (
            .O(N__25851),
            .I(N__25845));
    Span4Mux_h I__3896 (
            .O(N__25848),
            .I(N__25839));
    Span4Mux_h I__3895 (
            .O(N__25845),
            .I(N__25839));
    InMux I__3894 (
            .O(N__25844),
            .I(N__25836));
    Odrv4 I__3893 (
            .O(N__25839),
            .I(r2_14));
    LocalMux I__3892 (
            .O(N__25836),
            .I(r2_14));
    CascadeMux I__3891 (
            .O(N__25831),
            .I(N__25827));
    InMux I__3890 (
            .O(N__25830),
            .I(N__25824));
    InMux I__3889 (
            .O(N__25827),
            .I(N__25821));
    LocalMux I__3888 (
            .O(N__25824),
            .I(N__25817));
    LocalMux I__3887 (
            .O(N__25821),
            .I(N__25814));
    InMux I__3886 (
            .O(N__25820),
            .I(N__25811));
    Span4Mux_v I__3885 (
            .O(N__25817),
            .I(N__25808));
    Span4Mux_h I__3884 (
            .O(N__25814),
            .I(N__25805));
    LocalMux I__3883 (
            .O(N__25811),
            .I(r3_14));
    Odrv4 I__3882 (
            .O(N__25808),
            .I(r3_14));
    Odrv4 I__3881 (
            .O(N__25805),
            .I(r3_14));
    InMux I__3880 (
            .O(N__25798),
            .I(N__25793));
    InMux I__3879 (
            .O(N__25797),
            .I(N__25790));
    InMux I__3878 (
            .O(N__25796),
            .I(N__25787));
    LocalMux I__3877 (
            .O(N__25793),
            .I(N__25784));
    LocalMux I__3876 (
            .O(N__25790),
            .I(N__25781));
    LocalMux I__3875 (
            .O(N__25787),
            .I(N__25776));
    Span4Mux_s3_h I__3874 (
            .O(N__25784),
            .I(N__25776));
    Span4Mux_h I__3873 (
            .O(N__25781),
            .I(N__25773));
    Odrv4 I__3872 (
            .O(N__25776),
            .I(r7_14));
    Odrv4 I__3871 (
            .O(N__25773),
            .I(r7_14));
    CascadeMux I__3870 (
            .O(N__25768),
            .I(\ALU.a_6_ns_1_14_cascade_ ));
    InMux I__3869 (
            .O(N__25765),
            .I(N__25760));
    InMux I__3868 (
            .O(N__25764),
            .I(N__25757));
    InMux I__3867 (
            .O(N__25763),
            .I(N__25754));
    LocalMux I__3866 (
            .O(N__25760),
            .I(N__25751));
    LocalMux I__3865 (
            .O(N__25757),
            .I(N__25748));
    LocalMux I__3864 (
            .O(N__25754),
            .I(N__25745));
    Span4Mux_h I__3863 (
            .O(N__25751),
            .I(N__25742));
    Odrv4 I__3862 (
            .O(N__25748),
            .I(r6_14));
    Odrv4 I__3861 (
            .O(N__25745),
            .I(r6_14));
    Odrv4 I__3860 (
            .O(N__25742),
            .I(r6_14));
    CascadeMux I__3859 (
            .O(N__25735),
            .I(\ALU.r6_RNID4772Z0Z_14_cascade_ ));
    InMux I__3858 (
            .O(N__25732),
            .I(N__25729));
    LocalMux I__3857 (
            .O(N__25729),
            .I(N__25726));
    Odrv4 I__3856 (
            .O(N__25726),
            .I(\ALU.r5_RNI54M52Z0Z_14 ));
    CascadeMux I__3855 (
            .O(N__25723),
            .I(N__25720));
    InMux I__3854 (
            .O(N__25720),
            .I(N__25716));
    InMux I__3853 (
            .O(N__25719),
            .I(N__25713));
    LocalMux I__3852 (
            .O(N__25716),
            .I(N__25710));
    LocalMux I__3851 (
            .O(N__25713),
            .I(N__25707));
    Span4Mux_v I__3850 (
            .O(N__25710),
            .I(N__25701));
    Span4Mux_v I__3849 (
            .O(N__25707),
            .I(N__25701));
    InMux I__3848 (
            .O(N__25706),
            .I(N__25698));
    Odrv4 I__3847 (
            .O(N__25701),
            .I(r0_14));
    LocalMux I__3846 (
            .O(N__25698),
            .I(r0_14));
    CascadeMux I__3845 (
            .O(N__25693),
            .I(N__25688));
    CascadeMux I__3844 (
            .O(N__25692),
            .I(N__25685));
    InMux I__3843 (
            .O(N__25691),
            .I(N__25665));
    InMux I__3842 (
            .O(N__25688),
            .I(N__25665));
    InMux I__3841 (
            .O(N__25685),
            .I(N__25665));
    InMux I__3840 (
            .O(N__25684),
            .I(N__25665));
    InMux I__3839 (
            .O(N__25683),
            .I(N__25665));
    InMux I__3838 (
            .O(N__25682),
            .I(N__25665));
    InMux I__3837 (
            .O(N__25681),
            .I(N__25657));
    InMux I__3836 (
            .O(N__25680),
            .I(N__25657));
    InMux I__3835 (
            .O(N__25679),
            .I(N__25652));
    InMux I__3834 (
            .O(N__25678),
            .I(N__25652));
    LocalMux I__3833 (
            .O(N__25665),
            .I(N__25644));
    InMux I__3832 (
            .O(N__25664),
            .I(N__25637));
    InMux I__3831 (
            .O(N__25663),
            .I(N__25637));
    InMux I__3830 (
            .O(N__25662),
            .I(N__25637));
    LocalMux I__3829 (
            .O(N__25657),
            .I(N__25634));
    LocalMux I__3828 (
            .O(N__25652),
            .I(N__25631));
    InMux I__3827 (
            .O(N__25651),
            .I(N__25620));
    InMux I__3826 (
            .O(N__25650),
            .I(N__25620));
    InMux I__3825 (
            .O(N__25649),
            .I(N__25620));
    InMux I__3824 (
            .O(N__25648),
            .I(N__25620));
    InMux I__3823 (
            .O(N__25647),
            .I(N__25620));
    Span4Mux_h I__3822 (
            .O(N__25644),
            .I(N__25615));
    LocalMux I__3821 (
            .O(N__25637),
            .I(N__25615));
    Span4Mux_v I__3820 (
            .O(N__25634),
            .I(N__25610));
    Span4Mux_h I__3819 (
            .O(N__25631),
            .I(N__25610));
    LocalMux I__3818 (
            .O(N__25620),
            .I(aZ0Z_0));
    Odrv4 I__3817 (
            .O(N__25615),
            .I(aZ0Z_0));
    Odrv4 I__3816 (
            .O(N__25610),
            .I(aZ0Z_0));
    InMux I__3815 (
            .O(N__25603),
            .I(N__25591));
    InMux I__3814 (
            .O(N__25602),
            .I(N__25591));
    InMux I__3813 (
            .O(N__25601),
            .I(N__25586));
    InMux I__3812 (
            .O(N__25600),
            .I(N__25586));
    InMux I__3811 (
            .O(N__25599),
            .I(N__25581));
    InMux I__3810 (
            .O(N__25598),
            .I(N__25581));
    InMux I__3809 (
            .O(N__25597),
            .I(N__25572));
    CascadeMux I__3808 (
            .O(N__25596),
            .I(N__25566));
    LocalMux I__3807 (
            .O(N__25591),
            .I(N__25560));
    LocalMux I__3806 (
            .O(N__25586),
            .I(N__25557));
    LocalMux I__3805 (
            .O(N__25581),
            .I(N__25554));
    InMux I__3804 (
            .O(N__25580),
            .I(N__25541));
    InMux I__3803 (
            .O(N__25579),
            .I(N__25541));
    InMux I__3802 (
            .O(N__25578),
            .I(N__25541));
    InMux I__3801 (
            .O(N__25577),
            .I(N__25541));
    InMux I__3800 (
            .O(N__25576),
            .I(N__25541));
    InMux I__3799 (
            .O(N__25575),
            .I(N__25541));
    LocalMux I__3798 (
            .O(N__25572),
            .I(N__25538));
    InMux I__3797 (
            .O(N__25571),
            .I(N__25531));
    InMux I__3796 (
            .O(N__25570),
            .I(N__25531));
    InMux I__3795 (
            .O(N__25569),
            .I(N__25531));
    InMux I__3794 (
            .O(N__25566),
            .I(N__25522));
    InMux I__3793 (
            .O(N__25565),
            .I(N__25522));
    InMux I__3792 (
            .O(N__25564),
            .I(N__25522));
    InMux I__3791 (
            .O(N__25563),
            .I(N__25522));
    Span4Mux_v I__3790 (
            .O(N__25560),
            .I(N__25519));
    Span4Mux_h I__3789 (
            .O(N__25557),
            .I(N__25512));
    Span4Mux_v I__3788 (
            .O(N__25554),
            .I(N__25512));
    LocalMux I__3787 (
            .O(N__25541),
            .I(N__25512));
    Span4Mux_h I__3786 (
            .O(N__25538),
            .I(N__25509));
    LocalMux I__3785 (
            .O(N__25531),
            .I(N__25506));
    LocalMux I__3784 (
            .O(N__25522),
            .I(aZ0Z_2));
    Odrv4 I__3783 (
            .O(N__25519),
            .I(aZ0Z_2));
    Odrv4 I__3782 (
            .O(N__25512),
            .I(aZ0Z_2));
    Odrv4 I__3781 (
            .O(N__25509),
            .I(aZ0Z_2));
    Odrv4 I__3780 (
            .O(N__25506),
            .I(aZ0Z_2));
    CascadeMux I__3779 (
            .O(N__25495),
            .I(\ALU.a_3_ns_1_15_cascade_ ));
    InMux I__3778 (
            .O(N__25492),
            .I(N__25489));
    LocalMux I__3777 (
            .O(N__25489),
            .I(N__25486));
    Odrv12 I__3776 (
            .O(N__25486),
            .I(\ALU.r5_RNI98M52Z0Z_15 ));
    InMux I__3775 (
            .O(N__25483),
            .I(N__25480));
    LocalMux I__3774 (
            .O(N__25480),
            .I(N__25475));
    InMux I__3773 (
            .O(N__25479),
            .I(N__25472));
    InMux I__3772 (
            .O(N__25478),
            .I(N__25469));
    Span4Mux_v I__3771 (
            .O(N__25475),
            .I(N__25464));
    LocalMux I__3770 (
            .O(N__25472),
            .I(N__25464));
    LocalMux I__3769 (
            .O(N__25469),
            .I(N__25461));
    Span4Mux_h I__3768 (
            .O(N__25464),
            .I(N__25458));
    Odrv12 I__3767 (
            .O(N__25461),
            .I(r4_10));
    Odrv4 I__3766 (
            .O(N__25458),
            .I(r4_10));
    InMux I__3765 (
            .O(N__25453),
            .I(N__25449));
    InMux I__3764 (
            .O(N__25452),
            .I(N__25445));
    LocalMux I__3763 (
            .O(N__25449),
            .I(N__25442));
    InMux I__3762 (
            .O(N__25448),
            .I(N__25439));
    LocalMux I__3761 (
            .O(N__25445),
            .I(N__25436));
    Span4Mux_h I__3760 (
            .O(N__25442),
            .I(N__25431));
    LocalMux I__3759 (
            .O(N__25439),
            .I(N__25431));
    Odrv12 I__3758 (
            .O(N__25436),
            .I(r4_12));
    Odrv4 I__3757 (
            .O(N__25431),
            .I(r4_12));
    InMux I__3756 (
            .O(N__25426),
            .I(N__25423));
    LocalMux I__3755 (
            .O(N__25423),
            .I(N__25420));
    Span4Mux_h I__3754 (
            .O(N__25420),
            .I(N__25416));
    InMux I__3753 (
            .O(N__25419),
            .I(N__25413));
    Span4Mux_v I__3752 (
            .O(N__25416),
            .I(N__25407));
    LocalMux I__3751 (
            .O(N__25413),
            .I(N__25407));
    InMux I__3750 (
            .O(N__25412),
            .I(N__25404));
    Span4Mux_h I__3749 (
            .O(N__25407),
            .I(N__25401));
    LocalMux I__3748 (
            .O(N__25404),
            .I(N__25398));
    Odrv4 I__3747 (
            .O(N__25401),
            .I(r4_13));
    Odrv4 I__3746 (
            .O(N__25398),
            .I(r4_13));
    InMux I__3745 (
            .O(N__25393),
            .I(N__25388));
    InMux I__3744 (
            .O(N__25392),
            .I(N__25385));
    InMux I__3743 (
            .O(N__25391),
            .I(N__25382));
    LocalMux I__3742 (
            .O(N__25388),
            .I(N__25379));
    LocalMux I__3741 (
            .O(N__25385),
            .I(N__25376));
    LocalMux I__3740 (
            .O(N__25382),
            .I(N__25373));
    Span4Mux_h I__3739 (
            .O(N__25379),
            .I(N__25370));
    Span12Mux_v I__3738 (
            .O(N__25376),
            .I(N__25365));
    Span12Mux_s11_v I__3737 (
            .O(N__25373),
            .I(N__25365));
    Odrv4 I__3736 (
            .O(N__25370),
            .I(r4_5));
    Odrv12 I__3735 (
            .O(N__25365),
            .I(r4_5));
    InMux I__3734 (
            .O(N__25360),
            .I(N__25357));
    LocalMux I__3733 (
            .O(N__25357),
            .I(N__25353));
    InMux I__3732 (
            .O(N__25356),
            .I(N__25349));
    Span4Mux_h I__3731 (
            .O(N__25353),
            .I(N__25346));
    InMux I__3730 (
            .O(N__25352),
            .I(N__25343));
    LocalMux I__3729 (
            .O(N__25349),
            .I(N__25340));
    Span4Mux_v I__3728 (
            .O(N__25346),
            .I(N__25337));
    LocalMux I__3727 (
            .O(N__25343),
            .I(N__25334));
    Span4Mux_v I__3726 (
            .O(N__25340),
            .I(N__25329));
    Span4Mux_v I__3725 (
            .O(N__25337),
            .I(N__25329));
    Sp12to4 I__3724 (
            .O(N__25334),
            .I(N__25326));
    Odrv4 I__3723 (
            .O(N__25329),
            .I(r4_6));
    Odrv12 I__3722 (
            .O(N__25326),
            .I(r4_6));
    CascadeMux I__3721 (
            .O(N__25321),
            .I(\ALU.r6_RNI7L2O1Z0Z_4_cascade_ ));
    InMux I__3720 (
            .O(N__25318),
            .I(N__25314));
    InMux I__3719 (
            .O(N__25317),
            .I(N__25311));
    LocalMux I__3718 (
            .O(N__25314),
            .I(N__25308));
    LocalMux I__3717 (
            .O(N__25311),
            .I(N__25305));
    Span4Mux_h I__3716 (
            .O(N__25308),
            .I(N__25301));
    Span4Mux_h I__3715 (
            .O(N__25305),
            .I(N__25298));
    InMux I__3714 (
            .O(N__25304),
            .I(N__25295));
    Odrv4 I__3713 (
            .O(N__25301),
            .I(r2_12));
    Odrv4 I__3712 (
            .O(N__25298),
            .I(r2_12));
    LocalMux I__3711 (
            .O(N__25295),
            .I(r2_12));
    CascadeMux I__3710 (
            .O(N__25288),
            .I(N__25284));
    CascadeMux I__3709 (
            .O(N__25287),
            .I(N__25281));
    InMux I__3708 (
            .O(N__25284),
            .I(N__25276));
    InMux I__3707 (
            .O(N__25281),
            .I(N__25276));
    LocalMux I__3706 (
            .O(N__25276),
            .I(N__25272));
    InMux I__3705 (
            .O(N__25275),
            .I(N__25269));
    Odrv12 I__3704 (
            .O(N__25272),
            .I(r2_4));
    LocalMux I__3703 (
            .O(N__25269),
            .I(r2_4));
    CascadeMux I__3702 (
            .O(N__25264),
            .I(TXbuffer_18_6_ns_1_4_cascade_));
    InMux I__3701 (
            .O(N__25261),
            .I(N__25258));
    LocalMux I__3700 (
            .O(N__25258),
            .I(N__25254));
    InMux I__3699 (
            .O(N__25257),
            .I(N__25250));
    Span4Mux_h I__3698 (
            .O(N__25254),
            .I(N__25247));
    InMux I__3697 (
            .O(N__25253),
            .I(N__25244));
    LocalMux I__3696 (
            .O(N__25250),
            .I(N__25241));
    Span4Mux_h I__3695 (
            .O(N__25247),
            .I(N__25236));
    LocalMux I__3694 (
            .O(N__25244),
            .I(N__25236));
    Odrv4 I__3693 (
            .O(N__25241),
            .I(r6_12));
    Odrv4 I__3692 (
            .O(N__25236),
            .I(r6_12));
    InMux I__3691 (
            .O(N__25231),
            .I(N__25228));
    LocalMux I__3690 (
            .O(N__25228),
            .I(N__25225));
    Span4Mux_v I__3689 (
            .O(N__25225),
            .I(N__25222));
    Sp12to4 I__3688 (
            .O(N__25222),
            .I(N__25219));
    Odrv12 I__3687 (
            .O(N__25219),
            .I(TXbuffer_RNO_6Z0Z_4));
    CascadeMux I__3686 (
            .O(N__25216),
            .I(N__25213));
    InMux I__3685 (
            .O(N__25213),
            .I(N__25209));
    CascadeMux I__3684 (
            .O(N__25212),
            .I(N__25206));
    LocalMux I__3683 (
            .O(N__25209),
            .I(N__25203));
    InMux I__3682 (
            .O(N__25206),
            .I(N__25200));
    Span4Mux_v I__3681 (
            .O(N__25203),
            .I(N__25197));
    LocalMux I__3680 (
            .O(N__25200),
            .I(N__25193));
    Span4Mux_s2_h I__3679 (
            .O(N__25197),
            .I(N__25190));
    CascadeMux I__3678 (
            .O(N__25196),
            .I(N__25187));
    Span12Mux_v I__3677 (
            .O(N__25193),
            .I(N__25184));
    Span4Mux_h I__3676 (
            .O(N__25190),
            .I(N__25181));
    InMux I__3675 (
            .O(N__25187),
            .I(N__25178));
    Odrv12 I__3674 (
            .O(N__25184),
            .I(r1_11));
    Odrv4 I__3673 (
            .O(N__25181),
            .I(r1_11));
    LocalMux I__3672 (
            .O(N__25178),
            .I(r1_11));
    InMux I__3671 (
            .O(N__25171),
            .I(N__25167));
    InMux I__3670 (
            .O(N__25170),
            .I(N__25164));
    LocalMux I__3669 (
            .O(N__25167),
            .I(N__25160));
    LocalMux I__3668 (
            .O(N__25164),
            .I(N__25157));
    CascadeMux I__3667 (
            .O(N__25163),
            .I(N__25154));
    Span12Mux_s5_h I__3666 (
            .O(N__25160),
            .I(N__25151));
    Span4Mux_v I__3665 (
            .O(N__25157),
            .I(N__25148));
    InMux I__3664 (
            .O(N__25154),
            .I(N__25145));
    Odrv12 I__3663 (
            .O(N__25151),
            .I(r1_12));
    Odrv4 I__3662 (
            .O(N__25148),
            .I(r1_12));
    LocalMux I__3661 (
            .O(N__25145),
            .I(r1_12));
    InMux I__3660 (
            .O(N__25138),
            .I(N__25133));
    CascadeMux I__3659 (
            .O(N__25137),
            .I(N__25130));
    InMux I__3658 (
            .O(N__25136),
            .I(N__25127));
    LocalMux I__3657 (
            .O(N__25133),
            .I(N__25124));
    InMux I__3656 (
            .O(N__25130),
            .I(N__25121));
    LocalMux I__3655 (
            .O(N__25127),
            .I(N__25118));
    Span4Mux_v I__3654 (
            .O(N__25124),
            .I(N__25113));
    LocalMux I__3653 (
            .O(N__25121),
            .I(N__25113));
    Span4Mux_v I__3652 (
            .O(N__25118),
            .I(N__25110));
    Span4Mux_v I__3651 (
            .O(N__25113),
            .I(N__25107));
    Odrv4 I__3650 (
            .O(N__25110),
            .I(r1_13));
    Odrv4 I__3649 (
            .O(N__25107),
            .I(r1_13));
    InMux I__3648 (
            .O(N__25102),
            .I(N__25093));
    InMux I__3647 (
            .O(N__25101),
            .I(N__25080));
    InMux I__3646 (
            .O(N__25100),
            .I(N__25080));
    InMux I__3645 (
            .O(N__25099),
            .I(N__25080));
    InMux I__3644 (
            .O(N__25098),
            .I(N__25080));
    InMux I__3643 (
            .O(N__25097),
            .I(N__25080));
    InMux I__3642 (
            .O(N__25096),
            .I(N__25080));
    LocalMux I__3641 (
            .O(N__25093),
            .I(N__25068));
    LocalMux I__3640 (
            .O(N__25080),
            .I(N__25068));
    InMux I__3639 (
            .O(N__25079),
            .I(N__25061));
    InMux I__3638 (
            .O(N__25078),
            .I(N__25061));
    InMux I__3637 (
            .O(N__25077),
            .I(N__25052));
    InMux I__3636 (
            .O(N__25076),
            .I(N__25052));
    InMux I__3635 (
            .O(N__25075),
            .I(N__25052));
    InMux I__3634 (
            .O(N__25074),
            .I(N__25052));
    CascadeMux I__3633 (
            .O(N__25073),
            .I(N__25048));
    Span12Mux_v I__3632 (
            .O(N__25068),
            .I(N__25043));
    InMux I__3631 (
            .O(N__25067),
            .I(N__25040));
    InMux I__3630 (
            .O(N__25066),
            .I(N__25037));
    LocalMux I__3629 (
            .O(N__25061),
            .I(N__25032));
    LocalMux I__3628 (
            .O(N__25052),
            .I(N__25032));
    InMux I__3627 (
            .O(N__25051),
            .I(N__25023));
    InMux I__3626 (
            .O(N__25048),
            .I(N__25023));
    InMux I__3625 (
            .O(N__25047),
            .I(N__25023));
    InMux I__3624 (
            .O(N__25046),
            .I(N__25023));
    Odrv12 I__3623 (
            .O(N__25043),
            .I(bZ0Z_0));
    LocalMux I__3622 (
            .O(N__25040),
            .I(bZ0Z_0));
    LocalMux I__3621 (
            .O(N__25037),
            .I(bZ0Z_0));
    Odrv4 I__3620 (
            .O(N__25032),
            .I(bZ0Z_0));
    LocalMux I__3619 (
            .O(N__25023),
            .I(bZ0Z_0));
    InMux I__3618 (
            .O(N__25012),
            .I(N__25008));
    InMux I__3617 (
            .O(N__25011),
            .I(N__25005));
    LocalMux I__3616 (
            .O(N__25008),
            .I(N__24995));
    LocalMux I__3615 (
            .O(N__25005),
            .I(N__24992));
    InMux I__3614 (
            .O(N__25004),
            .I(N__24989));
    InMux I__3613 (
            .O(N__25003),
            .I(N__24984));
    InMux I__3612 (
            .O(N__25002),
            .I(N__24984));
    InMux I__3611 (
            .O(N__25001),
            .I(N__24975));
    InMux I__3610 (
            .O(N__25000),
            .I(N__24975));
    InMux I__3609 (
            .O(N__24999),
            .I(N__24975));
    InMux I__3608 (
            .O(N__24998),
            .I(N__24975));
    Span4Mux_v I__3607 (
            .O(N__24995),
            .I(N__24972));
    Odrv12 I__3606 (
            .O(N__24992),
            .I(a_0_repZ0Z1));
    LocalMux I__3605 (
            .O(N__24989),
            .I(a_0_repZ0Z1));
    LocalMux I__3604 (
            .O(N__24984),
            .I(a_0_repZ0Z1));
    LocalMux I__3603 (
            .O(N__24975),
            .I(a_0_repZ0Z1));
    Odrv4 I__3602 (
            .O(N__24972),
            .I(a_0_repZ0Z1));
    CascadeMux I__3601 (
            .O(N__24961),
            .I(\ALU.a_6_ns_1_4_cascade_ ));
    CascadeMux I__3600 (
            .O(N__24958),
            .I(N__24954));
    CascadeMux I__3599 (
            .O(N__24957),
            .I(N__24950));
    InMux I__3598 (
            .O(N__24954),
            .I(N__24947));
    InMux I__3597 (
            .O(N__24953),
            .I(N__24942));
    InMux I__3596 (
            .O(N__24950),
            .I(N__24942));
    LocalMux I__3595 (
            .O(N__24947),
            .I(N__24939));
    LocalMux I__3594 (
            .O(N__24942),
            .I(N__24936));
    Span4Mux_h I__3593 (
            .O(N__24939),
            .I(N__24933));
    Span4Mux_v I__3592 (
            .O(N__24936),
            .I(N__24930));
    Odrv4 I__3591 (
            .O(N__24933),
            .I(r3_4));
    Odrv4 I__3590 (
            .O(N__24930),
            .I(r3_4));
    InMux I__3589 (
            .O(N__24925),
            .I(N__24919));
    InMux I__3588 (
            .O(N__24924),
            .I(N__24916));
    InMux I__3587 (
            .O(N__24923),
            .I(N__24913));
    CascadeMux I__3586 (
            .O(N__24922),
            .I(N__24910));
    LocalMux I__3585 (
            .O(N__24919),
            .I(N__24902));
    LocalMux I__3584 (
            .O(N__24916),
            .I(N__24899));
    LocalMux I__3583 (
            .O(N__24913),
            .I(N__24896));
    InMux I__3582 (
            .O(N__24910),
            .I(N__24893));
    InMux I__3581 (
            .O(N__24909),
            .I(N__24882));
    InMux I__3580 (
            .O(N__24908),
            .I(N__24882));
    InMux I__3579 (
            .O(N__24907),
            .I(N__24882));
    InMux I__3578 (
            .O(N__24906),
            .I(N__24882));
    InMux I__3577 (
            .O(N__24905),
            .I(N__24882));
    Span4Mux_v I__3576 (
            .O(N__24902),
            .I(N__24879));
    Span4Mux_h I__3575 (
            .O(N__24899),
            .I(N__24874));
    Span4Mux_v I__3574 (
            .O(N__24896),
            .I(N__24874));
    LocalMux I__3573 (
            .O(N__24893),
            .I(b_0_repZ0Z1));
    LocalMux I__3572 (
            .O(N__24882),
            .I(b_0_repZ0Z1));
    Odrv4 I__3571 (
            .O(N__24879),
            .I(b_0_repZ0Z1));
    Odrv4 I__3570 (
            .O(N__24874),
            .I(b_0_repZ0Z1));
    CascadeMux I__3569 (
            .O(N__24865),
            .I(\ALU.b_6_ns_1_4_cascade_ ));
    InMux I__3568 (
            .O(N__24862),
            .I(N__24859));
    LocalMux I__3567 (
            .O(N__24859),
            .I(N__24856));
    Span4Mux_v I__3566 (
            .O(N__24856),
            .I(N__24853));
    Odrv4 I__3565 (
            .O(N__24853),
            .I(\ALU.r6_RNI7L2O1Z0Z_4 ));
    CascadeMux I__3564 (
            .O(N__24850),
            .I(TXbuffer_18_3_ns_1_3_cascade_));
    CascadeMux I__3563 (
            .O(N__24847),
            .I(TXbuffer_RNO_5Z0Z_3_cascade_));
    InMux I__3562 (
            .O(N__24844),
            .I(N__24841));
    LocalMux I__3561 (
            .O(N__24841),
            .I(N__24838));
    Span4Mux_v I__3560 (
            .O(N__24838),
            .I(N__24835));
    Span4Mux_v I__3559 (
            .O(N__24835),
            .I(N__24832));
    Sp12to4 I__3558 (
            .O(N__24832),
            .I(N__24829));
    Span12Mux_s5_h I__3557 (
            .O(N__24829),
            .I(N__24826));
    Odrv12 I__3556 (
            .O(N__24826),
            .I(TXbuffer_18_15_ns_1_3));
    InMux I__3555 (
            .O(N__24823),
            .I(N__24820));
    LocalMux I__3554 (
            .O(N__24820),
            .I(N__24817));
    Span4Mux_h I__3553 (
            .O(N__24817),
            .I(N__24812));
    InMux I__3552 (
            .O(N__24816),
            .I(N__24809));
    InMux I__3551 (
            .O(N__24815),
            .I(N__24806));
    Odrv4 I__3550 (
            .O(N__24812),
            .I(r2_11));
    LocalMux I__3549 (
            .O(N__24809),
            .I(r2_11));
    LocalMux I__3548 (
            .O(N__24806),
            .I(r2_11));
    InMux I__3547 (
            .O(N__24799),
            .I(N__24796));
    LocalMux I__3546 (
            .O(N__24796),
            .I(N__24791));
    InMux I__3545 (
            .O(N__24795),
            .I(N__24788));
    InMux I__3544 (
            .O(N__24794),
            .I(N__24785));
    Span4Mux_h I__3543 (
            .O(N__24791),
            .I(N__24780));
    LocalMux I__3542 (
            .O(N__24788),
            .I(N__24780));
    LocalMux I__3541 (
            .O(N__24785),
            .I(N__24777));
    Odrv4 I__3540 (
            .O(N__24780),
            .I(r2_3));
    Odrv12 I__3539 (
            .O(N__24777),
            .I(r2_3));
    InMux I__3538 (
            .O(N__24772),
            .I(N__24769));
    LocalMux I__3537 (
            .O(N__24769),
            .I(N__24764));
    InMux I__3536 (
            .O(N__24768),
            .I(N__24761));
    InMux I__3535 (
            .O(N__24767),
            .I(N__24758));
    Span4Mux_h I__3534 (
            .O(N__24764),
            .I(N__24751));
    LocalMux I__3533 (
            .O(N__24761),
            .I(N__24751));
    LocalMux I__3532 (
            .O(N__24758),
            .I(N__24751));
    Span4Mux_v I__3531 (
            .O(N__24751),
            .I(N__24748));
    Odrv4 I__3530 (
            .O(N__24748),
            .I(r6_11));
    CascadeMux I__3529 (
            .O(N__24745),
            .I(TXbuffer_18_6_ns_1_3_cascade_));
    InMux I__3528 (
            .O(N__24742),
            .I(N__24739));
    LocalMux I__3527 (
            .O(N__24739),
            .I(TXbuffer_RNO_6Z0Z_3));
    InMux I__3526 (
            .O(N__24736),
            .I(N__24731));
    InMux I__3525 (
            .O(N__24735),
            .I(N__24728));
    InMux I__3524 (
            .O(N__24734),
            .I(N__24725));
    LocalMux I__3523 (
            .O(N__24731),
            .I(N__24722));
    LocalMux I__3522 (
            .O(N__24728),
            .I(N__24717));
    LocalMux I__3521 (
            .O(N__24725),
            .I(N__24717));
    Odrv4 I__3520 (
            .O(N__24722),
            .I(r4_11));
    Odrv4 I__3519 (
            .O(N__24717),
            .I(r4_11));
    InMux I__3518 (
            .O(N__24712),
            .I(N__24707));
    InMux I__3517 (
            .O(N__24711),
            .I(N__24702));
    InMux I__3516 (
            .O(N__24710),
            .I(N__24696));
    LocalMux I__3515 (
            .O(N__24707),
            .I(N__24693));
    InMux I__3514 (
            .O(N__24706),
            .I(N__24688));
    InMux I__3513 (
            .O(N__24705),
            .I(N__24688));
    LocalMux I__3512 (
            .O(N__24702),
            .I(N__24685));
    InMux I__3511 (
            .O(N__24701),
            .I(N__24680));
    InMux I__3510 (
            .O(N__24700),
            .I(N__24680));
    InMux I__3509 (
            .O(N__24699),
            .I(N__24677));
    LocalMux I__3508 (
            .O(N__24696),
            .I(N__24674));
    Span4Mux_h I__3507 (
            .O(N__24693),
            .I(N__24671));
    LocalMux I__3506 (
            .O(N__24688),
            .I(N__24664));
    Span4Mux_h I__3505 (
            .O(N__24685),
            .I(N__24664));
    LocalMux I__3504 (
            .O(N__24680),
            .I(N__24664));
    LocalMux I__3503 (
            .O(N__24677),
            .I(b_1_repZ0Z1));
    Odrv4 I__3502 (
            .O(N__24674),
            .I(b_1_repZ0Z1));
    Odrv4 I__3501 (
            .O(N__24671),
            .I(b_1_repZ0Z1));
    Odrv4 I__3500 (
            .O(N__24664),
            .I(b_1_repZ0Z1));
    CascadeMux I__3499 (
            .O(N__24655),
            .I(N__24650));
    InMux I__3498 (
            .O(N__24654),
            .I(N__24646));
    CascadeMux I__3497 (
            .O(N__24653),
            .I(N__24643));
    InMux I__3496 (
            .O(N__24650),
            .I(N__24638));
    InMux I__3495 (
            .O(N__24649),
            .I(N__24635));
    LocalMux I__3494 (
            .O(N__24646),
            .I(N__24632));
    InMux I__3493 (
            .O(N__24643),
            .I(N__24627));
    InMux I__3492 (
            .O(N__24642),
            .I(N__24624));
    InMux I__3491 (
            .O(N__24641),
            .I(N__24620));
    LocalMux I__3490 (
            .O(N__24638),
            .I(N__24617));
    LocalMux I__3489 (
            .O(N__24635),
            .I(N__24614));
    Span4Mux_v I__3488 (
            .O(N__24632),
            .I(N__24611));
    InMux I__3487 (
            .O(N__24631),
            .I(N__24608));
    InMux I__3486 (
            .O(N__24630),
            .I(N__24605));
    LocalMux I__3485 (
            .O(N__24627),
            .I(N__24602));
    LocalMux I__3484 (
            .O(N__24624),
            .I(N__24599));
    InMux I__3483 (
            .O(N__24623),
            .I(N__24596));
    LocalMux I__3482 (
            .O(N__24620),
            .I(N__24593));
    Span4Mux_v I__3481 (
            .O(N__24617),
            .I(N__24582));
    Span4Mux_v I__3480 (
            .O(N__24614),
            .I(N__24582));
    Span4Mux_s2_h I__3479 (
            .O(N__24611),
            .I(N__24582));
    LocalMux I__3478 (
            .O(N__24608),
            .I(N__24582));
    LocalMux I__3477 (
            .O(N__24605),
            .I(N__24582));
    Span4Mux_h I__3476 (
            .O(N__24602),
            .I(N__24578));
    Sp12to4 I__3475 (
            .O(N__24599),
            .I(N__24573));
    LocalMux I__3474 (
            .O(N__24596),
            .I(N__24573));
    Span4Mux_v I__3473 (
            .O(N__24593),
            .I(N__24568));
    Span4Mux_v I__3472 (
            .O(N__24582),
            .I(N__24568));
    InMux I__3471 (
            .O(N__24581),
            .I(N__24565));
    Sp12to4 I__3470 (
            .O(N__24578),
            .I(N__24562));
    Span12Mux_s6_v I__3469 (
            .O(N__24573),
            .I(N__24559));
    Span4Mux_h I__3468 (
            .O(N__24568),
            .I(N__24556));
    LocalMux I__3467 (
            .O(N__24565),
            .I(b_1_repZ0Z2));
    Odrv12 I__3466 (
            .O(N__24562),
            .I(b_1_repZ0Z2));
    Odrv12 I__3465 (
            .O(N__24559),
            .I(b_1_repZ0Z2));
    Odrv4 I__3464 (
            .O(N__24556),
            .I(b_1_repZ0Z2));
    InMux I__3463 (
            .O(N__24547),
            .I(N__24544));
    LocalMux I__3462 (
            .O(N__24544),
            .I(N__24540));
    InMux I__3461 (
            .O(N__24543),
            .I(N__24536));
    Span4Mux_h I__3460 (
            .O(N__24540),
            .I(N__24533));
    InMux I__3459 (
            .O(N__24539),
            .I(N__24530));
    LocalMux I__3458 (
            .O(N__24536),
            .I(N__24527));
    Span4Mux_s2_h I__3457 (
            .O(N__24533),
            .I(N__24524));
    LocalMux I__3456 (
            .O(N__24530),
            .I(N__24521));
    Span4Mux_v I__3455 (
            .O(N__24527),
            .I(N__24518));
    Odrv4 I__3454 (
            .O(N__24524),
            .I(r0_11));
    Odrv12 I__3453 (
            .O(N__24521),
            .I(r0_11));
    Odrv4 I__3452 (
            .O(N__24518),
            .I(r0_11));
    InMux I__3451 (
            .O(N__24511),
            .I(N__24508));
    LocalMux I__3450 (
            .O(N__24508),
            .I(N__24505));
    Span4Mux_v I__3449 (
            .O(N__24505),
            .I(N__24502));
    Span4Mux_h I__3448 (
            .O(N__24502),
            .I(N__24499));
    Odrv4 I__3447 (
            .O(N__24499),
            .I(\ALU.madd_368 ));
    CascadeMux I__3446 (
            .O(N__24496),
            .I(N__24493));
    InMux I__3445 (
            .O(N__24493),
            .I(N__24490));
    LocalMux I__3444 (
            .O(N__24490),
            .I(\ALU.a12_b_2 ));
    CascadeMux I__3443 (
            .O(N__24487),
            .I(\ALU.a12_b_2_cascade_ ));
    InMux I__3442 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__3441 (
            .O(N__24481),
            .I(N__24478));
    Span4Mux_v I__3440 (
            .O(N__24478),
            .I(N__24475));
    Span4Mux_h I__3439 (
            .O(N__24475),
            .I(N__24472));
    Odrv4 I__3438 (
            .O(N__24472),
            .I(\ALU.madd_372 ));
    CascadeMux I__3437 (
            .O(N__24469),
            .I(N__24466));
    InMux I__3436 (
            .O(N__24466),
            .I(N__24463));
    LocalMux I__3435 (
            .O(N__24463),
            .I(N__24459));
    InMux I__3434 (
            .O(N__24462),
            .I(N__24456));
    Span4Mux_s3_v I__3433 (
            .O(N__24459),
            .I(N__24453));
    LocalMux I__3432 (
            .O(N__24456),
            .I(N__24450));
    Odrv4 I__3431 (
            .O(N__24453),
            .I(\ALU.g1_2 ));
    Odrv4 I__3430 (
            .O(N__24450),
            .I(\ALU.g1_2 ));
    InMux I__3429 (
            .O(N__24445),
            .I(N__24442));
    LocalMux I__3428 (
            .O(N__24442),
            .I(N__24439));
    Span4Mux_s2_h I__3427 (
            .O(N__24439),
            .I(N__24436));
    Odrv4 I__3426 (
            .O(N__24436),
            .I(\ALU.madd_311_0 ));
    CascadeMux I__3425 (
            .O(N__24433),
            .I(\ALU.a_3_cascade_ ));
    InMux I__3424 (
            .O(N__24430),
            .I(N__24427));
    LocalMux I__3423 (
            .O(N__24427),
            .I(N__24424));
    Span4Mux_h I__3422 (
            .O(N__24424),
            .I(N__24421));
    Odrv4 I__3421 (
            .O(N__24421),
            .I(\ALU.g1_1 ));
    CascadeMux I__3420 (
            .O(N__24418),
            .I(\ALU.b_4_cascade_ ));
    InMux I__3419 (
            .O(N__24415),
            .I(N__24412));
    LocalMux I__3418 (
            .O(N__24412),
            .I(N__24409));
    Odrv12 I__3417 (
            .O(N__24409),
            .I(\ALU.madd_214_0 ));
    CascadeMux I__3416 (
            .O(N__24406),
            .I(\ALU.b_2_cascade_ ));
    InMux I__3415 (
            .O(N__24403),
            .I(N__24400));
    LocalMux I__3414 (
            .O(N__24400),
            .I(N__24397));
    Odrv4 I__3413 (
            .O(N__24397),
            .I(\ALU.madd_134_0_tz_0 ));
    InMux I__3412 (
            .O(N__24394),
            .I(N__24388));
    InMux I__3411 (
            .O(N__24393),
            .I(N__24388));
    LocalMux I__3410 (
            .O(N__24388),
            .I(N__24385));
    Span4Mux_s2_h I__3409 (
            .O(N__24385),
            .I(N__24382));
    Span4Mux_h I__3408 (
            .O(N__24382),
            .I(N__24379));
    Odrv4 I__3407 (
            .O(N__24379),
            .I(\ALU.madd_172_0 ));
    InMux I__3406 (
            .O(N__24376),
            .I(N__24373));
    LocalMux I__3405 (
            .O(N__24373),
            .I(N__24370));
    Span4Mux_v I__3404 (
            .O(N__24370),
            .I(N__24367));
    Span4Mux_h I__3403 (
            .O(N__24367),
            .I(N__24364));
    Span4Mux_v I__3402 (
            .O(N__24364),
            .I(N__24361));
    Odrv4 I__3401 (
            .O(N__24361),
            .I(\ALU.r6_RNIA0841Z0Z_0 ));
    InMux I__3400 (
            .O(N__24358),
            .I(N__24355));
    LocalMux I__3399 (
            .O(N__24355),
            .I(\ALU.madd_92 ));
    InMux I__3398 (
            .O(N__24352),
            .I(N__24348));
    InMux I__3397 (
            .O(N__24351),
            .I(N__24345));
    LocalMux I__3396 (
            .O(N__24348),
            .I(N__24342));
    LocalMux I__3395 (
            .O(N__24345),
            .I(\ALU.madd_120 ));
    Odrv4 I__3394 (
            .O(N__24342),
            .I(\ALU.madd_120 ));
    InMux I__3393 (
            .O(N__24337),
            .I(N__24333));
    InMux I__3392 (
            .O(N__24336),
            .I(N__24330));
    LocalMux I__3391 (
            .O(N__24333),
            .I(N__24324));
    LocalMux I__3390 (
            .O(N__24330),
            .I(N__24324));
    InMux I__3389 (
            .O(N__24329),
            .I(N__24321));
    Span4Mux_h I__3388 (
            .O(N__24324),
            .I(N__24318));
    LocalMux I__3387 (
            .O(N__24321),
            .I(N__24315));
    Odrv4 I__3386 (
            .O(N__24318),
            .I(\ALU.r6_RNII9FT1Z0Z_3 ));
    Odrv4 I__3385 (
            .O(N__24315),
            .I(\ALU.r6_RNII9FT1Z0Z_3 ));
    CascadeMux I__3384 (
            .O(N__24310),
            .I(\ALU.b_3_cascade_ ));
    InMux I__3383 (
            .O(N__24307),
            .I(N__24304));
    LocalMux I__3382 (
            .O(N__24304),
            .I(N__24301));
    Span4Mux_v I__3381 (
            .O(N__24301),
            .I(N__24298));
    Span4Mux_h I__3380 (
            .O(N__24298),
            .I(N__24295));
    Odrv4 I__3379 (
            .O(N__24295),
            .I(\ALU.un2_addsub_axb_3 ));
    CascadeMux I__3378 (
            .O(N__24292),
            .I(\ALU.b_1_cascade_ ));
    InMux I__3377 (
            .O(N__24289),
            .I(N__24286));
    LocalMux I__3376 (
            .O(N__24286),
            .I(N__24283));
    Odrv4 I__3375 (
            .O(N__24283),
            .I(\ALU.a4_b_1 ));
    CascadeMux I__3374 (
            .O(N__24280),
            .I(\ALU.madd_38_cascade_ ));
    CascadeMux I__3373 (
            .O(N__24277),
            .I(\ALU.madd_87_cascade_ ));
    CascadeMux I__3372 (
            .O(N__24274),
            .I(\ALU.madd_92_cascade_ ));
    InMux I__3371 (
            .O(N__24271),
            .I(N__24268));
    LocalMux I__3370 (
            .O(N__24268),
            .I(\ALU.madd_78_0 ));
    InMux I__3369 (
            .O(N__24265),
            .I(N__24259));
    InMux I__3368 (
            .O(N__24264),
            .I(N__24259));
    LocalMux I__3367 (
            .O(N__24259),
            .I(N__24256));
    Odrv4 I__3366 (
            .O(N__24256),
            .I(\ALU.madd_68 ));
    CascadeMux I__3365 (
            .O(N__24253),
            .I(\ALU.madd_78_0_cascade_ ));
    InMux I__3364 (
            .O(N__24250),
            .I(N__24244));
    InMux I__3363 (
            .O(N__24249),
            .I(N__24244));
    LocalMux I__3362 (
            .O(N__24244),
            .I(\ALU.madd_60 ));
    CascadeMux I__3361 (
            .O(N__24241),
            .I(\ALU.madd_332_cascade_ ));
    InMux I__3360 (
            .O(N__24238),
            .I(N__24234));
    InMux I__3359 (
            .O(N__24237),
            .I(N__24231));
    LocalMux I__3358 (
            .O(N__24234),
            .I(\ALU.madd_68_0 ));
    LocalMux I__3357 (
            .O(N__24231),
            .I(\ALU.madd_68_0 ));
    InMux I__3356 (
            .O(N__24226),
            .I(N__24223));
    LocalMux I__3355 (
            .O(N__24223),
            .I(N__24220));
    Odrv4 I__3354 (
            .O(N__24220),
            .I(\ALU.madd_46_0 ));
    InMux I__3353 (
            .O(N__24217),
            .I(N__24213));
    InMux I__3352 (
            .O(N__24216),
            .I(N__24210));
    LocalMux I__3351 (
            .O(N__24213),
            .I(\ALU.madd_100 ));
    LocalMux I__3350 (
            .O(N__24210),
            .I(\ALU.madd_100 ));
    InMux I__3349 (
            .O(N__24205),
            .I(N__24201));
    InMux I__3348 (
            .O(N__24204),
            .I(N__24198));
    LocalMux I__3347 (
            .O(N__24201),
            .I(\ALU.madd_105 ));
    LocalMux I__3346 (
            .O(N__24198),
            .I(\ALU.madd_105 ));
    CascadeMux I__3345 (
            .O(N__24193),
            .I(\ALU.madd_46_0_cascade_ ));
    InMux I__3344 (
            .O(N__24190),
            .I(N__24187));
    LocalMux I__3343 (
            .O(N__24187),
            .I(\ALU.madd_82_0 ));
    InMux I__3342 (
            .O(N__24184),
            .I(N__24178));
    InMux I__3341 (
            .O(N__24183),
            .I(N__24178));
    LocalMux I__3340 (
            .O(N__24178),
            .I(\ALU.a5_b_3 ));
    InMux I__3339 (
            .O(N__24175),
            .I(N__24172));
    LocalMux I__3338 (
            .O(N__24172),
            .I(N__24169));
    Odrv4 I__3337 (
            .O(N__24169),
            .I(\ALU.g2_0_0_0 ));
    InMux I__3336 (
            .O(N__24166),
            .I(N__24162));
    CascadeMux I__3335 (
            .O(N__24165),
            .I(N__24159));
    LocalMux I__3334 (
            .O(N__24162),
            .I(N__24156));
    InMux I__3333 (
            .O(N__24159),
            .I(N__24153));
    Odrv4 I__3332 (
            .O(N__24156),
            .I(\ALU.a0_b_7 ));
    LocalMux I__3331 (
            .O(N__24153),
            .I(\ALU.a0_b_7 ));
    CascadeMux I__3330 (
            .O(N__24148),
            .I(N__24145));
    InMux I__3329 (
            .O(N__24145),
            .I(N__24142));
    LocalMux I__3328 (
            .O(N__24142),
            .I(\ALU.a5_b_0 ));
    CascadeMux I__3327 (
            .O(N__24139),
            .I(N__24135));
    InMux I__3326 (
            .O(N__24138),
            .I(N__24132));
    InMux I__3325 (
            .O(N__24135),
            .I(N__24129));
    LocalMux I__3324 (
            .O(N__24132),
            .I(N__24123));
    LocalMux I__3323 (
            .O(N__24129),
            .I(N__24123));
    CascadeMux I__3322 (
            .O(N__24128),
            .I(N__24120));
    Span4Mux_v I__3321 (
            .O(N__24123),
            .I(N__24117));
    InMux I__3320 (
            .O(N__24120),
            .I(N__24114));
    Span4Mux_v I__3319 (
            .O(N__24117),
            .I(N__24111));
    LocalMux I__3318 (
            .O(N__24114),
            .I(r3_5));
    Odrv4 I__3317 (
            .O(N__24111),
            .I(r3_5));
    InMux I__3316 (
            .O(N__24106),
            .I(N__24103));
    LocalMux I__3315 (
            .O(N__24103),
            .I(N__24098));
    CascadeMux I__3314 (
            .O(N__24102),
            .I(N__24095));
    InMux I__3313 (
            .O(N__24101),
            .I(N__24092));
    Span4Mux_h I__3312 (
            .O(N__24098),
            .I(N__24089));
    InMux I__3311 (
            .O(N__24095),
            .I(N__24086));
    LocalMux I__3310 (
            .O(N__24092),
            .I(r3_13));
    Odrv4 I__3309 (
            .O(N__24089),
            .I(r3_13));
    LocalMux I__3308 (
            .O(N__24086),
            .I(r3_13));
    InMux I__3307 (
            .O(N__24079),
            .I(N__24075));
    InMux I__3306 (
            .O(N__24078),
            .I(N__24072));
    LocalMux I__3305 (
            .O(N__24075),
            .I(N__24068));
    LocalMux I__3304 (
            .O(N__24072),
            .I(N__24065));
    InMux I__3303 (
            .O(N__24071),
            .I(N__24062));
    Span4Mux_v I__3302 (
            .O(N__24068),
            .I(N__24057));
    Span4Mux_v I__3301 (
            .O(N__24065),
            .I(N__24057));
    LocalMux I__3300 (
            .O(N__24062),
            .I(N__24054));
    Odrv4 I__3299 (
            .O(N__24057),
            .I(r6_13));
    Odrv4 I__3298 (
            .O(N__24054),
            .I(r6_13));
    CascadeMux I__3297 (
            .O(N__24049),
            .I(N__24046));
    InMux I__3296 (
            .O(N__24046),
            .I(N__24043));
    LocalMux I__3295 (
            .O(N__24043),
            .I(N__24040));
    Odrv4 I__3294 (
            .O(N__24040),
            .I(TXbuffer_18_6_ns_1_5));
    InMux I__3293 (
            .O(N__24037),
            .I(N__24033));
    InMux I__3292 (
            .O(N__24036),
            .I(N__24029));
    LocalMux I__3291 (
            .O(N__24033),
            .I(N__24026));
    InMux I__3290 (
            .O(N__24032),
            .I(N__24023));
    LocalMux I__3289 (
            .O(N__24029),
            .I(N__24020));
    Span4Mux_h I__3288 (
            .O(N__24026),
            .I(N__24017));
    LocalMux I__3287 (
            .O(N__24023),
            .I(N__24014));
    Span4Mux_v I__3286 (
            .O(N__24020),
            .I(N__24011));
    Span4Mux_v I__3285 (
            .O(N__24017),
            .I(N__24008));
    Span4Mux_v I__3284 (
            .O(N__24014),
            .I(N__24005));
    Odrv4 I__3283 (
            .O(N__24011),
            .I(r6_5));
    Odrv4 I__3282 (
            .O(N__24008),
            .I(r6_5));
    Odrv4 I__3281 (
            .O(N__24005),
            .I(r6_5));
    InMux I__3280 (
            .O(N__23998),
            .I(N__23995));
    LocalMux I__3279 (
            .O(N__23995),
            .I(TXbuffer_RNO_5Z0Z_5));
    CascadeMux I__3278 (
            .O(N__23992),
            .I(TXbuffer_RNO_6Z0Z_5_cascade_));
    InMux I__3277 (
            .O(N__23989),
            .I(N__23985));
    InMux I__3276 (
            .O(N__23988),
            .I(N__23982));
    LocalMux I__3275 (
            .O(N__23985),
            .I(N__23978));
    LocalMux I__3274 (
            .O(N__23982),
            .I(N__23975));
    InMux I__3273 (
            .O(N__23981),
            .I(N__23972));
    Odrv4 I__3272 (
            .O(N__23978),
            .I(r7_13));
    Odrv4 I__3271 (
            .O(N__23975),
            .I(r7_13));
    LocalMux I__3270 (
            .O(N__23972),
            .I(r7_13));
    CascadeMux I__3269 (
            .O(N__23965),
            .I(N__23961));
    InMux I__3268 (
            .O(N__23964),
            .I(N__23958));
    InMux I__3267 (
            .O(N__23961),
            .I(N__23954));
    LocalMux I__3266 (
            .O(N__23958),
            .I(N__23951));
    InMux I__3265 (
            .O(N__23957),
            .I(N__23948));
    LocalMux I__3264 (
            .O(N__23954),
            .I(N__23945));
    Span4Mux_h I__3263 (
            .O(N__23951),
            .I(N__23940));
    LocalMux I__3262 (
            .O(N__23948),
            .I(N__23940));
    Span4Mux_v I__3261 (
            .O(N__23945),
            .I(N__23935));
    Span4Mux_v I__3260 (
            .O(N__23940),
            .I(N__23935));
    Odrv4 I__3259 (
            .O(N__23935),
            .I(r7_5));
    InMux I__3258 (
            .O(N__23932),
            .I(N__23929));
    LocalMux I__3257 (
            .O(N__23929),
            .I(TXbuffer_18_13_ns_1_5));
    InMux I__3256 (
            .O(N__23926),
            .I(N__23923));
    LocalMux I__3255 (
            .O(N__23923),
            .I(TXbuffer_18_10_ns_1_5));
    CascadeMux I__3254 (
            .O(N__23920),
            .I(\ALU.a_3_ns_1_13_cascade_ ));
    InMux I__3253 (
            .O(N__23917),
            .I(N__23913));
    InMux I__3252 (
            .O(N__23916),
            .I(N__23910));
    LocalMux I__3251 (
            .O(N__23913),
            .I(N__23907));
    LocalMux I__3250 (
            .O(N__23910),
            .I(N__23903));
    Span4Mux_v I__3249 (
            .O(N__23907),
            .I(N__23900));
    InMux I__3248 (
            .O(N__23906),
            .I(N__23897));
    Span4Mux_h I__3247 (
            .O(N__23903),
            .I(N__23894));
    Odrv4 I__3246 (
            .O(N__23900),
            .I(r2_13));
    LocalMux I__3245 (
            .O(N__23897),
            .I(r2_13));
    Odrv4 I__3244 (
            .O(N__23894),
            .I(r2_13));
    CascadeMux I__3243 (
            .O(N__23887),
            .I(\ALU.a_6_ns_1_13_cascade_ ));
    CascadeMux I__3242 (
            .O(N__23884),
            .I(\ALU.r6_RNI90772Z0Z_13_cascade_ ));
    InMux I__3241 (
            .O(N__23881),
            .I(N__23878));
    LocalMux I__3240 (
            .O(N__23878),
            .I(\ALU.r5_RNI10M52Z0Z_13 ));
    CascadeMux I__3239 (
            .O(N__23875),
            .I(\ALU.r5_RNIPV8A9Z0Z_13_cascade_ ));
    InMux I__3238 (
            .O(N__23872),
            .I(N__23867));
    InMux I__3237 (
            .O(N__23871),
            .I(N__23864));
    CascadeMux I__3236 (
            .O(N__23870),
            .I(N__23861));
    LocalMux I__3235 (
            .O(N__23867),
            .I(N__23858));
    LocalMux I__3234 (
            .O(N__23864),
            .I(N__23855));
    InMux I__3233 (
            .O(N__23861),
            .I(N__23852));
    Span4Mux_h I__3232 (
            .O(N__23858),
            .I(N__23849));
    Span4Mux_h I__3231 (
            .O(N__23855),
            .I(N__23846));
    LocalMux I__3230 (
            .O(N__23852),
            .I(N__23843));
    Odrv4 I__3229 (
            .O(N__23849),
            .I(r3_12));
    Odrv4 I__3228 (
            .O(N__23846),
            .I(r3_12));
    Odrv12 I__3227 (
            .O(N__23843),
            .I(r3_12));
    CascadeMux I__3226 (
            .O(N__23836),
            .I(N__23833));
    InMux I__3225 (
            .O(N__23833),
            .I(N__23830));
    LocalMux I__3224 (
            .O(N__23830),
            .I(N__23827));
    Span4Mux_v I__3223 (
            .O(N__23827),
            .I(N__23824));
    Odrv4 I__3222 (
            .O(N__23824),
            .I(\ALU.r0_12_prm_7_15_s1_c_RNOZ0 ));
    CascadeMux I__3221 (
            .O(N__23821),
            .I(N__23818));
    InMux I__3220 (
            .O(N__23818),
            .I(N__23815));
    LocalMux I__3219 (
            .O(N__23815),
            .I(N__23812));
    Span4Mux_h I__3218 (
            .O(N__23812),
            .I(N__23809));
    Odrv4 I__3217 (
            .O(N__23809),
            .I(\ALU.r0_12_prm_6_15_s1_c_RNOZ0 ));
    CascadeMux I__3216 (
            .O(N__23806),
            .I(N__23803));
    InMux I__3215 (
            .O(N__23803),
            .I(N__23800));
    LocalMux I__3214 (
            .O(N__23800),
            .I(N__23797));
    Span4Mux_h I__3213 (
            .O(N__23797),
            .I(N__23794));
    Odrv4 I__3212 (
            .O(N__23794),
            .I(\ALU.r0_12_prm_4_15_s1_c_RNOZ0 ));
    InMux I__3211 (
            .O(N__23791),
            .I(N__23788));
    LocalMux I__3210 (
            .O(N__23788),
            .I(N__23785));
    Span4Mux_v I__3209 (
            .O(N__23785),
            .I(N__23782));
    Odrv4 I__3208 (
            .O(N__23782),
            .I(\ALU.madd_axb_14 ));
    InMux I__3207 (
            .O(N__23779),
            .I(\ALU.r0_12_s1_15 ));
    InMux I__3206 (
            .O(N__23776),
            .I(N__23771));
    InMux I__3205 (
            .O(N__23775),
            .I(N__23768));
    InMux I__3204 (
            .O(N__23774),
            .I(N__23765));
    LocalMux I__3203 (
            .O(N__23771),
            .I(N__23762));
    LocalMux I__3202 (
            .O(N__23768),
            .I(N__23757));
    LocalMux I__3201 (
            .O(N__23765),
            .I(N__23757));
    Span4Mux_v I__3200 (
            .O(N__23762),
            .I(N__23752));
    Span4Mux_v I__3199 (
            .O(N__23757),
            .I(N__23752));
    Odrv4 I__3198 (
            .O(N__23752),
            .I(r2_5));
    InMux I__3197 (
            .O(N__23749),
            .I(N__23746));
    LocalMux I__3196 (
            .O(N__23746),
            .I(N__23742));
    InMux I__3195 (
            .O(N__23745),
            .I(N__23738));
    Span4Mux_h I__3194 (
            .O(N__23742),
            .I(N__23735));
    InMux I__3193 (
            .O(N__23741),
            .I(N__23732));
    LocalMux I__3192 (
            .O(N__23738),
            .I(N__23729));
    Span4Mux_s3_v I__3191 (
            .O(N__23735),
            .I(N__23726));
    LocalMux I__3190 (
            .O(N__23732),
            .I(N__23723));
    Span4Mux_h I__3189 (
            .O(N__23729),
            .I(N__23720));
    Span4Mux_v I__3188 (
            .O(N__23726),
            .I(N__23715));
    Span4Mux_h I__3187 (
            .O(N__23723),
            .I(N__23715));
    Odrv4 I__3186 (
            .O(N__23720),
            .I(r2_6));
    Odrv4 I__3185 (
            .O(N__23715),
            .I(r2_6));
    CascadeMux I__3184 (
            .O(N__23710),
            .I(N__23707));
    InMux I__3183 (
            .O(N__23707),
            .I(N__23702));
    InMux I__3182 (
            .O(N__23706),
            .I(N__23699));
    InMux I__3181 (
            .O(N__23705),
            .I(N__23696));
    LocalMux I__3180 (
            .O(N__23702),
            .I(N__23693));
    LocalMux I__3179 (
            .O(N__23699),
            .I(N__23690));
    LocalMux I__3178 (
            .O(N__23696),
            .I(N__23687));
    Span4Mux_v I__3177 (
            .O(N__23693),
            .I(N__23684));
    Span4Mux_h I__3176 (
            .O(N__23690),
            .I(N__23679));
    Span4Mux_h I__3175 (
            .O(N__23687),
            .I(N__23679));
    Odrv4 I__3174 (
            .O(N__23684),
            .I(r2_9));
    Odrv4 I__3173 (
            .O(N__23679),
            .I(r2_9));
    CascadeMux I__3172 (
            .O(N__23674),
            .I(\ALU.a_3_ns_1_11_cascade_ ));
    InMux I__3171 (
            .O(N__23671),
            .I(N__23668));
    LocalMux I__3170 (
            .O(N__23668),
            .I(\ALU.r5_RNI3VN52Z0Z_11 ));
    CascadeMux I__3169 (
            .O(N__23665),
            .I(N__23662));
    InMux I__3168 (
            .O(N__23662),
            .I(N__23659));
    LocalMux I__3167 (
            .O(N__23659),
            .I(N__23654));
    InMux I__3166 (
            .O(N__23658),
            .I(N__23651));
    InMux I__3165 (
            .O(N__23657),
            .I(N__23648));
    Span4Mux_v I__3164 (
            .O(N__23654),
            .I(N__23645));
    LocalMux I__3163 (
            .O(N__23651),
            .I(N__23642));
    LocalMux I__3162 (
            .O(N__23648),
            .I(N__23639));
    Span4Mux_h I__3161 (
            .O(N__23645),
            .I(N__23636));
    Odrv4 I__3160 (
            .O(N__23642),
            .I(r3_3));
    Odrv12 I__3159 (
            .O(N__23639),
            .I(r3_3));
    Odrv4 I__3158 (
            .O(N__23636),
            .I(r3_3));
    CascadeMux I__3157 (
            .O(N__23629),
            .I(\ALU.a_6_ns_1_3_cascade_ ));
    CascadeMux I__3156 (
            .O(N__23626),
            .I(\ALU.a_3_ns_1_12_cascade_ ));
    InMux I__3155 (
            .O(N__23623),
            .I(N__23618));
    InMux I__3154 (
            .O(N__23622),
            .I(N__23615));
    InMux I__3153 (
            .O(N__23621),
            .I(N__23612));
    LocalMux I__3152 (
            .O(N__23618),
            .I(N__23609));
    LocalMux I__3151 (
            .O(N__23615),
            .I(N__23606));
    LocalMux I__3150 (
            .O(N__23612),
            .I(N__23603));
    Span4Mux_s3_h I__3149 (
            .O(N__23609),
            .I(N__23600));
    Span4Mux_s3_h I__3148 (
            .O(N__23606),
            .I(N__23595));
    Span4Mux_h I__3147 (
            .O(N__23603),
            .I(N__23595));
    Odrv4 I__3146 (
            .O(N__23600),
            .I(r7_12));
    Odrv4 I__3145 (
            .O(N__23595),
            .I(r7_12));
    CascadeMux I__3144 (
            .O(N__23590),
            .I(\ALU.a_6_ns_1_12_cascade_ ));
    CascadeMux I__3143 (
            .O(N__23587),
            .I(\ALU.r6_RNI5S672Z0Z_12_cascade_ ));
    InMux I__3142 (
            .O(N__23584),
            .I(N__23581));
    LocalMux I__3141 (
            .O(N__23581),
            .I(\ALU.r5_RNIS3672Z0Z_12 ));
    InMux I__3140 (
            .O(N__23578),
            .I(N__23575));
    LocalMux I__3139 (
            .O(N__23575),
            .I(N__23572));
    Span4Mux_h I__3138 (
            .O(N__23572),
            .I(N__23568));
    CascadeMux I__3137 (
            .O(N__23571),
            .I(N__23565));
    Span4Mux_v I__3136 (
            .O(N__23568),
            .I(N__23561));
    InMux I__3135 (
            .O(N__23565),
            .I(N__23558));
    InMux I__3134 (
            .O(N__23564),
            .I(N__23555));
    Odrv4 I__3133 (
            .O(N__23561),
            .I(r2_8));
    LocalMux I__3132 (
            .O(N__23558),
            .I(r2_8));
    LocalMux I__3131 (
            .O(N__23555),
            .I(r2_8));
    CascadeMux I__3130 (
            .O(N__23548),
            .I(N__23543));
    InMux I__3129 (
            .O(N__23547),
            .I(N__23540));
    InMux I__3128 (
            .O(N__23546),
            .I(N__23535));
    InMux I__3127 (
            .O(N__23543),
            .I(N__23535));
    LocalMux I__3126 (
            .O(N__23540),
            .I(N__23532));
    LocalMux I__3125 (
            .O(N__23535),
            .I(N__23529));
    Span4Mux_v I__3124 (
            .O(N__23532),
            .I(N__23526));
    Span4Mux_h I__3123 (
            .O(N__23529),
            .I(N__23523));
    Odrv4 I__3122 (
            .O(N__23526),
            .I(r3_8));
    Odrv4 I__3121 (
            .O(N__23523),
            .I(r3_8));
    CascadeMux I__3120 (
            .O(N__23518),
            .I(\ALU.b_6_ns_1_8_cascade_ ));
    InMux I__3119 (
            .O(N__23515),
            .I(N__23512));
    LocalMux I__3118 (
            .O(N__23512),
            .I(N__23509));
    Odrv12 I__3117 (
            .O(N__23509),
            .I(\ALU.r6_RNIN53O1Z0Z_8 ));
    CascadeMux I__3116 (
            .O(N__23506),
            .I(\ALU.a_6_ns_1_1_cascade_ ));
    CascadeMux I__3115 (
            .O(N__23503),
            .I(\ALU.a_3_ns_1_10_cascade_ ));
    CascadeMux I__3114 (
            .O(N__23500),
            .I(\ALU.r5_RNIVQN52Z0Z_10_cascade_ ));
    InMux I__3113 (
            .O(N__23497),
            .I(N__23493));
    InMux I__3112 (
            .O(N__23496),
            .I(N__23490));
    LocalMux I__3111 (
            .O(N__23493),
            .I(N__23487));
    LocalMux I__3110 (
            .O(N__23490),
            .I(N__23484));
    Sp12to4 I__3109 (
            .O(N__23487),
            .I(N__23480));
    Span4Mux_h I__3108 (
            .O(N__23484),
            .I(N__23477));
    InMux I__3107 (
            .O(N__23483),
            .I(N__23474));
    Odrv12 I__3106 (
            .O(N__23480),
            .I(r0_6));
    Odrv4 I__3105 (
            .O(N__23477),
            .I(r0_6));
    LocalMux I__3104 (
            .O(N__23474),
            .I(r0_6));
    CascadeMux I__3103 (
            .O(N__23467),
            .I(\ALU.a_6_ns_1_5_cascade_ ));
    CascadeMux I__3102 (
            .O(N__23464),
            .I(N__23460));
    InMux I__3101 (
            .O(N__23463),
            .I(N__23457));
    InMux I__3100 (
            .O(N__23460),
            .I(N__23454));
    LocalMux I__3099 (
            .O(N__23457),
            .I(N__23450));
    LocalMux I__3098 (
            .O(N__23454),
            .I(N__23447));
    CascadeMux I__3097 (
            .O(N__23453),
            .I(N__23444));
    Span4Mux_v I__3096 (
            .O(N__23450),
            .I(N__23441));
    Span4Mux_v I__3095 (
            .O(N__23447),
            .I(N__23438));
    InMux I__3094 (
            .O(N__23444),
            .I(N__23435));
    Span4Mux_v I__3093 (
            .O(N__23441),
            .I(N__23432));
    Span4Mux_v I__3092 (
            .O(N__23438),
            .I(N__23429));
    LocalMux I__3091 (
            .O(N__23435),
            .I(r3_6));
    Odrv4 I__3090 (
            .O(N__23432),
            .I(r3_6));
    Odrv4 I__3089 (
            .O(N__23429),
            .I(r3_6));
    CascadeMux I__3088 (
            .O(N__23422),
            .I(\ALU.a_6_ns_1_6_cascade_ ));
    InMux I__3087 (
            .O(N__23419),
            .I(N__23416));
    LocalMux I__3086 (
            .O(N__23416),
            .I(\ALU.a_6_ns_1_9 ));
    CascadeMux I__3085 (
            .O(N__23413),
            .I(\ALU.a_6_ns_1_8_cascade_ ));
    InMux I__3084 (
            .O(N__23410),
            .I(N__23407));
    LocalMux I__3083 (
            .O(N__23407),
            .I(N__23401));
    InMux I__3082 (
            .O(N__23406),
            .I(N__23394));
    InMux I__3081 (
            .O(N__23405),
            .I(N__23394));
    InMux I__3080 (
            .O(N__23404),
            .I(N__23394));
    Span4Mux_h I__3079 (
            .O(N__23401),
            .I(N__23389));
    LocalMux I__3078 (
            .O(N__23394),
            .I(N__23389));
    Odrv4 I__3077 (
            .O(N__23389),
            .I(\ALU.r6_RNIKG3D2Z0Z_8 ));
    InMux I__3076 (
            .O(N__23386),
            .I(N__23383));
    LocalMux I__3075 (
            .O(N__23383),
            .I(N__23380));
    Span4Mux_v I__3074 (
            .O(N__23380),
            .I(N__23375));
    InMux I__3073 (
            .O(N__23379),
            .I(N__23370));
    InMux I__3072 (
            .O(N__23378),
            .I(N__23370));
    Span4Mux_h I__3071 (
            .O(N__23375),
            .I(N__23367));
    LocalMux I__3070 (
            .O(N__23370),
            .I(r2_2));
    Odrv4 I__3069 (
            .O(N__23367),
            .I(r2_2));
    CascadeMux I__3068 (
            .O(N__23362),
            .I(N__23358));
    CascadeMux I__3067 (
            .O(N__23361),
            .I(N__23354));
    InMux I__3066 (
            .O(N__23358),
            .I(N__23351));
    InMux I__3065 (
            .O(N__23357),
            .I(N__23346));
    InMux I__3064 (
            .O(N__23354),
            .I(N__23346));
    LocalMux I__3063 (
            .O(N__23351),
            .I(N__23343));
    LocalMux I__3062 (
            .O(N__23346),
            .I(N__23340));
    Span4Mux_h I__3061 (
            .O(N__23343),
            .I(N__23337));
    Odrv4 I__3060 (
            .O(N__23340),
            .I(r3_2));
    Odrv4 I__3059 (
            .O(N__23337),
            .I(r3_2));
    CascadeMux I__3058 (
            .O(N__23332),
            .I(\ALU.b_6_ns_1_2_cascade_ ));
    CascadeMux I__3057 (
            .O(N__23329),
            .I(\ALU.b_6_ns_1_3_cascade_ ));
    InMux I__3056 (
            .O(N__23326),
            .I(N__23322));
    InMux I__3055 (
            .O(N__23325),
            .I(N__23319));
    LocalMux I__3054 (
            .O(N__23322),
            .I(N__23315));
    LocalMux I__3053 (
            .O(N__23319),
            .I(N__23312));
    InMux I__3052 (
            .O(N__23318),
            .I(N__23309));
    Span4Mux_s3_h I__3051 (
            .O(N__23315),
            .I(N__23306));
    Span4Mux_v I__3050 (
            .O(N__23312),
            .I(N__23303));
    LocalMux I__3049 (
            .O(N__23309),
            .I(N__23300));
    Odrv4 I__3048 (
            .O(N__23306),
            .I(r7_0));
    Odrv4 I__3047 (
            .O(N__23303),
            .I(r7_0));
    Odrv12 I__3046 (
            .O(N__23300),
            .I(r7_0));
    CascadeMux I__3045 (
            .O(N__23293),
            .I(\ALU.b_6_ns_1_0_cascade_ ));
    InMux I__3044 (
            .O(N__23290),
            .I(N__23287));
    LocalMux I__3043 (
            .O(N__23287),
            .I(N__23284));
    Span4Mux_h I__3042 (
            .O(N__23284),
            .I(N__23279));
    InMux I__3041 (
            .O(N__23283),
            .I(N__23274));
    InMux I__3040 (
            .O(N__23282),
            .I(N__23274));
    Span4Mux_v I__3039 (
            .O(N__23279),
            .I(N__23271));
    LocalMux I__3038 (
            .O(N__23274),
            .I(r6_0));
    Odrv4 I__3037 (
            .O(N__23271),
            .I(r6_0));
    CascadeMux I__3036 (
            .O(N__23266),
            .I(\ALU.a_3_ns_1_6_cascade_ ));
    InMux I__3035 (
            .O(N__23263),
            .I(N__23257));
    InMux I__3034 (
            .O(N__23262),
            .I(N__23257));
    LocalMux I__3033 (
            .O(N__23257),
            .I(N__23253));
    InMux I__3032 (
            .O(N__23256),
            .I(N__23250));
    Span4Mux_h I__3031 (
            .O(N__23253),
            .I(N__23247));
    LocalMux I__3030 (
            .O(N__23250),
            .I(N__23244));
    Odrv4 I__3029 (
            .O(N__23247),
            .I(\ALU.a8_b_4 ));
    Odrv12 I__3028 (
            .O(N__23244),
            .I(\ALU.a8_b_4 ));
    CascadeMux I__3027 (
            .O(N__23239),
            .I(\ALU.g0_7_x1_cascade_ ));
    InMux I__3026 (
            .O(N__23236),
            .I(N__23233));
    LocalMux I__3025 (
            .O(N__23233),
            .I(\ALU.madd_76_1 ));
    CascadeMux I__3024 (
            .O(N__23230),
            .I(N__23225));
    InMux I__3023 (
            .O(N__23229),
            .I(N__23221));
    InMux I__3022 (
            .O(N__23228),
            .I(N__23218));
    InMux I__3021 (
            .O(N__23225),
            .I(N__23215));
    InMux I__3020 (
            .O(N__23224),
            .I(N__23212));
    LocalMux I__3019 (
            .O(N__23221),
            .I(N__23207));
    LocalMux I__3018 (
            .O(N__23218),
            .I(N__23207));
    LocalMux I__3017 (
            .O(N__23215),
            .I(N__23202));
    LocalMux I__3016 (
            .O(N__23212),
            .I(N__23202));
    Odrv4 I__3015 (
            .O(N__23207),
            .I(\ALU.r6_RNIPK3D2Z0Z_9 ));
    Odrv4 I__3014 (
            .O(N__23202),
            .I(\ALU.r6_RNIPK3D2Z0Z_9 ));
    CascadeMux I__3013 (
            .O(N__23197),
            .I(N__23193));
    CascadeMux I__3012 (
            .O(N__23196),
            .I(N__23190));
    InMux I__3011 (
            .O(N__23193),
            .I(N__23185));
    InMux I__3010 (
            .O(N__23190),
            .I(N__23185));
    LocalMux I__3009 (
            .O(N__23185),
            .I(N__23182));
    Span4Mux_s1_h I__3008 (
            .O(N__23182),
            .I(N__23179));
    Odrv4 I__3007 (
            .O(N__23179),
            .I(\ALU.a9_b_4 ));
    CascadeMux I__3006 (
            .O(N__23176),
            .I(\ALU.a_8_cascade_ ));
    InMux I__3005 (
            .O(N__23173),
            .I(N__23170));
    LocalMux I__3004 (
            .O(N__23170),
            .I(N__23167));
    Odrv4 I__3003 (
            .O(N__23167),
            .I(\ALU.madd_224_0 ));
    CascadeMux I__3002 (
            .O(N__23164),
            .I(N__23160));
    InMux I__3001 (
            .O(N__23163),
            .I(N__23155));
    InMux I__3000 (
            .O(N__23160),
            .I(N__23155));
    LocalMux I__2999 (
            .O(N__23155),
            .I(N__23152));
    Span4Mux_v I__2998 (
            .O(N__23152),
            .I(N__23149));
    Odrv4 I__2997 (
            .O(N__23149),
            .I(\ALU.madd_224 ));
    InMux I__2996 (
            .O(N__23146),
            .I(N__23143));
    LocalMux I__2995 (
            .O(N__23143),
            .I(\ALU.madd_121 ));
    InMux I__2994 (
            .O(N__23140),
            .I(N__23137));
    LocalMux I__2993 (
            .O(N__23137),
            .I(N__23134));
    Odrv12 I__2992 (
            .O(N__23134),
            .I(\ALU.b_3_ns_1_8 ));
    CascadeMux I__2991 (
            .O(N__23131),
            .I(\ALU.a_9_cascade_ ));
    InMux I__2990 (
            .O(N__23128),
            .I(N__23125));
    LocalMux I__2989 (
            .O(N__23125),
            .I(N__23122));
    Span4Mux_h I__2988 (
            .O(N__23122),
            .I(N__23119));
    Odrv4 I__2987 (
            .O(N__23119),
            .I(\ALU.N_675_1 ));
    CascadeMux I__2986 (
            .O(N__23116),
            .I(\ALU.bZ0Z_0_cascade_ ));
    InMux I__2985 (
            .O(N__23113),
            .I(N__23110));
    LocalMux I__2984 (
            .O(N__23110),
            .I(\ALU.madd_130_0_0 ));
    InMux I__2983 (
            .O(N__23107),
            .I(N__23103));
    InMux I__2982 (
            .O(N__23106),
            .I(N__23097));
    LocalMux I__2981 (
            .O(N__23103),
            .I(N__23094));
    InMux I__2980 (
            .O(N__23102),
            .I(N__23091));
    InMux I__2979 (
            .O(N__23101),
            .I(N__23088));
    InMux I__2978 (
            .O(N__23100),
            .I(N__23085));
    LocalMux I__2977 (
            .O(N__23097),
            .I(N__23082));
    Span4Mux_v I__2976 (
            .O(N__23094),
            .I(N__23077));
    LocalMux I__2975 (
            .O(N__23091),
            .I(N__23077));
    LocalMux I__2974 (
            .O(N__23088),
            .I(N__23074));
    LocalMux I__2973 (
            .O(N__23085),
            .I(N__23071));
    Span4Mux_s3_h I__2972 (
            .O(N__23082),
            .I(N__23068));
    Span4Mux_h I__2971 (
            .O(N__23077),
            .I(N__23063));
    Span4Mux_v I__2970 (
            .O(N__23074),
            .I(N__23063));
    Span4Mux_v I__2969 (
            .O(N__23071),
            .I(N__23060));
    Odrv4 I__2968 (
            .O(N__23068),
            .I(\ALU.r6_RNIGC3D2Z0Z_7 ));
    Odrv4 I__2967 (
            .O(N__23063),
            .I(\ALU.r6_RNIGC3D2Z0Z_7 ));
    Odrv4 I__2966 (
            .O(N__23060),
            .I(\ALU.r6_RNIGC3D2Z0Z_7 ));
    CascadeMux I__2965 (
            .O(N__23053),
            .I(\ALU.a_7_cascade_ ));
    CascadeMux I__2964 (
            .O(N__23050),
            .I(N__23046));
    CascadeMux I__2963 (
            .O(N__23049),
            .I(N__23043));
    InMux I__2962 (
            .O(N__23046),
            .I(N__23038));
    InMux I__2961 (
            .O(N__23043),
            .I(N__23038));
    LocalMux I__2960 (
            .O(N__23038),
            .I(N__23034));
    InMux I__2959 (
            .O(N__23037),
            .I(N__23031));
    Span4Mux_s2_h I__2958 (
            .O(N__23034),
            .I(N__23026));
    LocalMux I__2957 (
            .O(N__23031),
            .I(N__23026));
    Span4Mux_v I__2956 (
            .O(N__23026),
            .I(N__23023));
    Odrv4 I__2955 (
            .O(N__23023),
            .I(\ALU.madd_76 ));
    CascadeMux I__2954 (
            .O(N__23020),
            .I(N__23017));
    InMux I__2953 (
            .O(N__23017),
            .I(N__23014));
    LocalMux I__2952 (
            .O(N__23014),
            .I(\ALU.madd_213_0_tz ));
    InMux I__2951 (
            .O(N__23011),
            .I(N__23008));
    LocalMux I__2950 (
            .O(N__23008),
            .I(N__23005));
    Span4Mux_v I__2949 (
            .O(N__23005),
            .I(N__23002));
    Odrv4 I__2948 (
            .O(N__23002),
            .I(\ALU.madd_209_0 ));
    InMux I__2947 (
            .O(N__22999),
            .I(N__22996));
    LocalMux I__2946 (
            .O(N__22996),
            .I(\ALU.madd_223_0_tz ));
    InMux I__2945 (
            .O(N__22993),
            .I(N__22990));
    LocalMux I__2944 (
            .O(N__22990),
            .I(N__22987));
    Span4Mux_s1_v I__2943 (
            .O(N__22987),
            .I(N__22984));
    Odrv4 I__2942 (
            .O(N__22984),
            .I(\ALU.madd_105_0 ));
    InMux I__2941 (
            .O(N__22981),
            .I(N__22978));
    LocalMux I__2940 (
            .O(N__22978),
            .I(\ALU.r4_RNIU5NK1Z0Z_8 ));
    CascadeMux I__2939 (
            .O(N__22975),
            .I(\ALU.un9_addsub_axb_1_cascade_ ));
    InMux I__2938 (
            .O(N__22972),
            .I(N__22969));
    LocalMux I__2937 (
            .O(N__22969),
            .I(\ALU.a7_b_3 ));
    CascadeMux I__2936 (
            .O(N__22966),
            .I(\ALU.a_1_cascade_ ));
    InMux I__2935 (
            .O(N__22963),
            .I(N__22960));
    LocalMux I__2934 (
            .O(N__22960),
            .I(N__22957));
    Odrv4 I__2933 (
            .O(N__22957),
            .I(\ALU.madd_228_0_tz ));
    InMux I__2932 (
            .O(N__22954),
            .I(N__22951));
    LocalMux I__2931 (
            .O(N__22951),
            .I(\ALU.g3 ));
    InMux I__2930 (
            .O(N__22948),
            .I(N__22945));
    LocalMux I__2929 (
            .O(N__22945),
            .I(\ALU.madd_72_0_tz ));
    CascadeMux I__2928 (
            .O(N__22942),
            .I(\ALU.madd_40_cascade_ ));
    CascadeMux I__2927 (
            .O(N__22939),
            .I(N__22936));
    InMux I__2926 (
            .O(N__22936),
            .I(N__22930));
    InMux I__2925 (
            .O(N__22935),
            .I(N__22930));
    LocalMux I__2924 (
            .O(N__22930),
            .I(\ALU.madd_72 ));
    InMux I__2923 (
            .O(N__22927),
            .I(N__22924));
    LocalMux I__2922 (
            .O(N__22924),
            .I(N__22919));
    InMux I__2921 (
            .O(N__22923),
            .I(N__22914));
    InMux I__2920 (
            .O(N__22922),
            .I(N__22914));
    Odrv12 I__2919 (
            .O(N__22919),
            .I(\ALU.madd_95 ));
    LocalMux I__2918 (
            .O(N__22914),
            .I(\ALU.madd_95 ));
    CascadeMux I__2917 (
            .O(N__22909),
            .I(\ALU.madd_72_cascade_ ));
    InMux I__2916 (
            .O(N__22906),
            .I(N__22901));
    InMux I__2915 (
            .O(N__22905),
            .I(N__22896));
    InMux I__2914 (
            .O(N__22904),
            .I(N__22896));
    LocalMux I__2913 (
            .O(N__22901),
            .I(\ALU.madd_77 ));
    LocalMux I__2912 (
            .O(N__22896),
            .I(\ALU.madd_77 ));
    CascadeMux I__2911 (
            .O(N__22891),
            .I(\ALU.b_8_cascade_ ));
    InMux I__2910 (
            .O(N__22888),
            .I(N__22885));
    LocalMux I__2909 (
            .O(N__22885),
            .I(N__22882));
    Span4Mux_s2_v I__2908 (
            .O(N__22882),
            .I(N__22879));
    Odrv4 I__2907 (
            .O(N__22879),
            .I(\ALU.madd_82 ));
    CascadeMux I__2906 (
            .O(N__22876),
            .I(\ALU.madd_127_cascade_ ));
    InMux I__2905 (
            .O(N__22873),
            .I(N__22868));
    InMux I__2904 (
            .O(N__22872),
            .I(N__22865));
    InMux I__2903 (
            .O(N__22871),
            .I(N__22862));
    LocalMux I__2902 (
            .O(N__22868),
            .I(N__22857));
    LocalMux I__2901 (
            .O(N__22865),
            .I(N__22857));
    LocalMux I__2900 (
            .O(N__22862),
            .I(N__22854));
    Span4Mux_v I__2899 (
            .O(N__22857),
            .I(N__22851));
    Odrv4 I__2898 (
            .O(N__22854),
            .I(\ALU.madd_223 ));
    Odrv4 I__2897 (
            .O(N__22851),
            .I(\ALU.madd_223 ));
    CascadeMux I__2896 (
            .O(N__22846),
            .I(\ALU.a4_b_4_cascade_ ));
    InMux I__2895 (
            .O(N__22843),
            .I(N__22838));
    InMux I__2894 (
            .O(N__22842),
            .I(N__22833));
    InMux I__2893 (
            .O(N__22841),
            .I(N__22833));
    LocalMux I__2892 (
            .O(N__22838),
            .I(N__22830));
    LocalMux I__2891 (
            .O(N__22833),
            .I(N__22827));
    Odrv4 I__2890 (
            .O(N__22830),
            .I(\ALU.madd_104 ));
    Odrv12 I__2889 (
            .O(N__22827),
            .I(\ALU.madd_104 ));
    CascadeMux I__2888 (
            .O(N__22822),
            .I(\ALU.madd_68_cascade_ ));
    CascadeMux I__2887 (
            .O(N__22819),
            .I(\ALU.madd_82_0_cascade_ ));
    InMux I__2886 (
            .O(N__22816),
            .I(N__22807));
    InMux I__2885 (
            .O(N__22815),
            .I(N__22807));
    InMux I__2884 (
            .O(N__22814),
            .I(N__22807));
    LocalMux I__2883 (
            .O(N__22807),
            .I(N__22804));
    Odrv4 I__2882 (
            .O(N__22804),
            .I(\ALU.madd_119 ));
    CascadeMux I__2881 (
            .O(N__22801),
            .I(\ALU.a_6_cascade_ ));
    InMux I__2880 (
            .O(N__22798),
            .I(N__22795));
    LocalMux I__2879 (
            .O(N__22795),
            .I(\ALU.r0_12_prm_6_11_s0_c_RNOZ0 ));
    CascadeMux I__2878 (
            .O(N__22792),
            .I(N__22789));
    InMux I__2877 (
            .O(N__22789),
            .I(N__22786));
    LocalMux I__2876 (
            .O(N__22786),
            .I(\ALU.r0_12_prm_7_11_s0_c_RNOZ0 ));
    CascadeMux I__2875 (
            .O(N__22783),
            .I(N__22780));
    InMux I__2874 (
            .O(N__22780),
            .I(N__22777));
    LocalMux I__2873 (
            .O(N__22777),
            .I(N__22774));
    Span4Mux_v I__2872 (
            .O(N__22774),
            .I(N__22771));
    Odrv4 I__2871 (
            .O(N__22771),
            .I(\ALU.r0_12_prm_6_11_s1_c_RNOZ0 ));
    CascadeMux I__2870 (
            .O(N__22768),
            .I(N__22765));
    InMux I__2869 (
            .O(N__22765),
            .I(N__22762));
    LocalMux I__2868 (
            .O(N__22762),
            .I(N__22759));
    Odrv4 I__2867 (
            .O(N__22759),
            .I(TXbuffer_18_3_ns_1_5));
    CascadeMux I__2866 (
            .O(N__22756),
            .I(TXbuffer_18_10_ns_1_6_cascade_));
    InMux I__2865 (
            .O(N__22753),
            .I(N__22750));
    LocalMux I__2864 (
            .O(N__22750),
            .I(N__22747));
    Sp12to4 I__2863 (
            .O(N__22747),
            .I(N__22744));
    Odrv12 I__2862 (
            .O(N__22744),
            .I(TXbuffer_RNO_1Z0Z_6));
    CascadeMux I__2861 (
            .O(N__22741),
            .I(TXbuffer_RNO_0Z0Z_6_cascade_));
    InMux I__2860 (
            .O(N__22738),
            .I(N__22735));
    LocalMux I__2859 (
            .O(N__22735),
            .I(N__22732));
    Odrv12 I__2858 (
            .O(N__22732),
            .I(TXbuffer_18_6_ns_1_6));
    CascadeMux I__2857 (
            .O(N__22729),
            .I(TXbuffer_RNO_6Z0Z_6_cascade_));
    InMux I__2856 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__2855 (
            .O(N__22723),
            .I(TXbuffer_18_15_ns_1_6));
    CascadeMux I__2854 (
            .O(N__22720),
            .I(TXbuffer_18_3_ns_1_6_cascade_));
    InMux I__2853 (
            .O(N__22717),
            .I(N__22714));
    LocalMux I__2852 (
            .O(N__22714),
            .I(TXbuffer_RNO_5Z0Z_6));
    CascadeMux I__2851 (
            .O(N__22711),
            .I(N__22708));
    InMux I__2850 (
            .O(N__22708),
            .I(N__22705));
    LocalMux I__2849 (
            .O(N__22705),
            .I(N__22702));
    Span4Mux_v I__2848 (
            .O(N__22702),
            .I(N__22699));
    Odrv4 I__2847 (
            .O(N__22699),
            .I(\ALU.r0_12_prm_4_11_s1_c_RNOZ0 ));
    InMux I__2846 (
            .O(N__22696),
            .I(N__22693));
    LocalMux I__2845 (
            .O(N__22693),
            .I(\ALU.r5_RNIAFVE5Z0Z_11 ));
    InMux I__2844 (
            .O(N__22690),
            .I(N__22687));
    LocalMux I__2843 (
            .O(N__22687),
            .I(\ALU.r0_12_prm_5_11_s0_c_RNOZ0 ));
    InMux I__2842 (
            .O(N__22684),
            .I(N__22681));
    LocalMux I__2841 (
            .O(N__22681),
            .I(N__22676));
    InMux I__2840 (
            .O(N__22680),
            .I(N__22673));
    InMux I__2839 (
            .O(N__22679),
            .I(N__22670));
    Span4Mux_v I__2838 (
            .O(N__22676),
            .I(N__22667));
    LocalMux I__2837 (
            .O(N__22673),
            .I(N__22662));
    LocalMux I__2836 (
            .O(N__22670),
            .I(N__22662));
    Span4Mux_h I__2835 (
            .O(N__22667),
            .I(N__22659));
    Span4Mux_v I__2834 (
            .O(N__22662),
            .I(N__22656));
    Odrv4 I__2833 (
            .O(N__22659),
            .I(r7_10));
    Odrv4 I__2832 (
            .O(N__22656),
            .I(r7_10));
    CascadeMux I__2831 (
            .O(N__22651),
            .I(N__22646));
    InMux I__2830 (
            .O(N__22650),
            .I(N__22643));
    InMux I__2829 (
            .O(N__22649),
            .I(N__22640));
    InMux I__2828 (
            .O(N__22646),
            .I(N__22637));
    LocalMux I__2827 (
            .O(N__22643),
            .I(N__22632));
    LocalMux I__2826 (
            .O(N__22640),
            .I(N__22632));
    LocalMux I__2825 (
            .O(N__22637),
            .I(N__22629));
    Span4Mux_v I__2824 (
            .O(N__22632),
            .I(N__22626));
    Odrv12 I__2823 (
            .O(N__22629),
            .I(r7_11));
    Odrv4 I__2822 (
            .O(N__22626),
            .I(r7_11));
    InMux I__2821 (
            .O(N__22621),
            .I(N__22614));
    InMux I__2820 (
            .O(N__22620),
            .I(N__22614));
    InMux I__2819 (
            .O(N__22619),
            .I(N__22611));
    LocalMux I__2818 (
            .O(N__22614),
            .I(r7_15));
    LocalMux I__2817 (
            .O(N__22611),
            .I(r7_15));
    CascadeMux I__2816 (
            .O(N__22606),
            .I(TXbuffer_18_3_ns_1_2_cascade_));
    InMux I__2815 (
            .O(N__22603),
            .I(N__22600));
    LocalMux I__2814 (
            .O(N__22600),
            .I(N__22597));
    Span4Mux_v I__2813 (
            .O(N__22597),
            .I(N__22594));
    Span4Mux_v I__2812 (
            .O(N__22594),
            .I(N__22591));
    Odrv4 I__2811 (
            .O(N__22591),
            .I(TXbuffer_RNO_5Z0Z_2));
    CascadeMux I__2810 (
            .O(N__22588),
            .I(N__22585));
    InMux I__2809 (
            .O(N__22585),
            .I(N__22582));
    LocalMux I__2808 (
            .O(N__22582),
            .I(N__22579));
    Sp12to4 I__2807 (
            .O(N__22579),
            .I(N__22576));
    Odrv12 I__2806 (
            .O(N__22576),
            .I(TXbuffer_18_3_ns_1_4));
    InMux I__2805 (
            .O(N__22573),
            .I(N__22569));
    InMux I__2804 (
            .O(N__22572),
            .I(N__22565));
    LocalMux I__2803 (
            .O(N__22569),
            .I(N__22562));
    InMux I__2802 (
            .O(N__22568),
            .I(N__22559));
    LocalMux I__2801 (
            .O(N__22565),
            .I(N__22556));
    Span4Mux_s3_h I__2800 (
            .O(N__22562),
            .I(N__22551));
    LocalMux I__2799 (
            .O(N__22559),
            .I(N__22551));
    Span4Mux_v I__2798 (
            .O(N__22556),
            .I(N__22548));
    Span4Mux_h I__2797 (
            .O(N__22551),
            .I(N__22545));
    Span4Mux_h I__2796 (
            .O(N__22548),
            .I(N__22542));
    Span4Mux_s3_h I__2795 (
            .O(N__22545),
            .I(N__22539));
    Odrv4 I__2794 (
            .O(N__22542),
            .I(r6_10));
    Odrv4 I__2793 (
            .O(N__22539),
            .I(r6_10));
    InMux I__2792 (
            .O(N__22534),
            .I(N__22531));
    LocalMux I__2791 (
            .O(N__22531),
            .I(N__22526));
    InMux I__2790 (
            .O(N__22530),
            .I(N__22521));
    InMux I__2789 (
            .O(N__22529),
            .I(N__22521));
    Span4Mux_h I__2788 (
            .O(N__22526),
            .I(N__22516));
    LocalMux I__2787 (
            .O(N__22521),
            .I(N__22516));
    Odrv4 I__2786 (
            .O(N__22516),
            .I(r6_15));
    CascadeMux I__2785 (
            .O(N__22513),
            .I(N__22508));
    InMux I__2784 (
            .O(N__22512),
            .I(N__22503));
    InMux I__2783 (
            .O(N__22511),
            .I(N__22503));
    InMux I__2782 (
            .O(N__22508),
            .I(N__22500));
    LocalMux I__2781 (
            .O(N__22503),
            .I(N__22497));
    LocalMux I__2780 (
            .O(N__22500),
            .I(N__22494));
    Span4Mux_s2_h I__2779 (
            .O(N__22497),
            .I(N__22489));
    Span4Mux_v I__2778 (
            .O(N__22494),
            .I(N__22489));
    Odrv4 I__2777 (
            .O(N__22489),
            .I(r3_15));
    CascadeMux I__2776 (
            .O(N__22486),
            .I(N__22483));
    InMux I__2775 (
            .O(N__22483),
            .I(N__22478));
    CascadeMux I__2774 (
            .O(N__22482),
            .I(N__22475));
    CascadeMux I__2773 (
            .O(N__22481),
            .I(N__22472));
    LocalMux I__2772 (
            .O(N__22478),
            .I(N__22469));
    InMux I__2771 (
            .O(N__22475),
            .I(N__22466));
    InMux I__2770 (
            .O(N__22472),
            .I(N__22463));
    Odrv4 I__2769 (
            .O(N__22469),
            .I(r3_7));
    LocalMux I__2768 (
            .O(N__22466),
            .I(r3_7));
    LocalMux I__2767 (
            .O(N__22463),
            .I(r3_7));
    CascadeMux I__2766 (
            .O(N__22456),
            .I(TXbuffer_18_13_ns_1_6_cascade_));
    CascadeMux I__2765 (
            .O(N__22453),
            .I(\ALU.a_6_ns_1_7_cascade_ ));
    CascadeMux I__2764 (
            .O(N__22450),
            .I(\ALU.b_6_ns_1_7_cascade_ ));
    InMux I__2763 (
            .O(N__22447),
            .I(N__22444));
    LocalMux I__2762 (
            .O(N__22444),
            .I(N__22441));
    Span4Mux_v I__2761 (
            .O(N__22441),
            .I(N__22438));
    Odrv4 I__2760 (
            .O(N__22438),
            .I(\ALU.r6_RNIJ13O1Z0Z_7 ));
    InMux I__2759 (
            .O(N__22435),
            .I(N__22432));
    LocalMux I__2758 (
            .O(N__22432),
            .I(N__22428));
    InMux I__2757 (
            .O(N__22431),
            .I(N__22425));
    Span4Mux_h I__2756 (
            .O(N__22428),
            .I(N__22419));
    LocalMux I__2755 (
            .O(N__22425),
            .I(N__22419));
    InMux I__2754 (
            .O(N__22424),
            .I(N__22416));
    Odrv4 I__2753 (
            .O(N__22419),
            .I(r2_15));
    LocalMux I__2752 (
            .O(N__22416),
            .I(r2_15));
    CascadeMux I__2751 (
            .O(N__22411),
            .I(N__22408));
    InMux I__2750 (
            .O(N__22408),
            .I(N__22403));
    InMux I__2749 (
            .O(N__22407),
            .I(N__22398));
    InMux I__2748 (
            .O(N__22406),
            .I(N__22398));
    LocalMux I__2747 (
            .O(N__22403),
            .I(r2_7));
    LocalMux I__2746 (
            .O(N__22398),
            .I(r2_7));
    CascadeMux I__2745 (
            .O(N__22393),
            .I(TXbuffer_18_6_ns_1_7_cascade_));
    InMux I__2744 (
            .O(N__22390),
            .I(N__22386));
    CascadeMux I__2743 (
            .O(N__22389),
            .I(N__22382));
    LocalMux I__2742 (
            .O(N__22386),
            .I(N__22379));
    InMux I__2741 (
            .O(N__22385),
            .I(N__22376));
    InMux I__2740 (
            .O(N__22382),
            .I(N__22373));
    Span4Mux_s3_h I__2739 (
            .O(N__22379),
            .I(N__22366));
    LocalMux I__2738 (
            .O(N__22376),
            .I(N__22366));
    LocalMux I__2737 (
            .O(N__22373),
            .I(N__22366));
    Odrv4 I__2736 (
            .O(N__22366),
            .I(r3_10));
    CascadeMux I__2735 (
            .O(N__22363),
            .I(N__22358));
    InMux I__2734 (
            .O(N__22362),
            .I(N__22355));
    InMux I__2733 (
            .O(N__22361),
            .I(N__22352));
    InMux I__2732 (
            .O(N__22358),
            .I(N__22349));
    LocalMux I__2731 (
            .O(N__22355),
            .I(N__22346));
    LocalMux I__2730 (
            .O(N__22352),
            .I(N__22343));
    LocalMux I__2729 (
            .O(N__22349),
            .I(N__22340));
    Odrv4 I__2728 (
            .O(N__22346),
            .I(r3_11));
    Odrv4 I__2727 (
            .O(N__22343),
            .I(r3_11));
    Odrv4 I__2726 (
            .O(N__22340),
            .I(r3_11));
    InMux I__2725 (
            .O(N__22333),
            .I(N__22330));
    LocalMux I__2724 (
            .O(N__22330),
            .I(N__22327));
    Span4Mux_s3_h I__2723 (
            .O(N__22327),
            .I(N__22324));
    Span4Mux_v I__2722 (
            .O(N__22324),
            .I(N__22320));
    InMux I__2721 (
            .O(N__22323),
            .I(N__22317));
    Span4Mux_v I__2720 (
            .O(N__22320),
            .I(N__22313));
    LocalMux I__2719 (
            .O(N__22317),
            .I(N__22310));
    InMux I__2718 (
            .O(N__22316),
            .I(N__22307));
    Odrv4 I__2717 (
            .O(N__22313),
            .I(r0_5));
    Odrv4 I__2716 (
            .O(N__22310),
            .I(r0_5));
    LocalMux I__2715 (
            .O(N__22307),
            .I(r0_5));
    CascadeMux I__2714 (
            .O(N__22300),
            .I(\ALU.a_3_ns_1_5_cascade_ ));
    InMux I__2713 (
            .O(N__22297),
            .I(N__22294));
    LocalMux I__2712 (
            .O(N__22294),
            .I(N__22291));
    Span4Mux_s2_h I__2711 (
            .O(N__22291),
            .I(N__22286));
    InMux I__2710 (
            .O(N__22290),
            .I(N__22283));
    InMux I__2709 (
            .O(N__22289),
            .I(N__22280));
    Odrv4 I__2708 (
            .O(N__22286),
            .I(r2_10));
    LocalMux I__2707 (
            .O(N__22283),
            .I(r2_10));
    LocalMux I__2706 (
            .O(N__22280),
            .I(r2_10));
    CascadeMux I__2705 (
            .O(N__22273),
            .I(\ALU.a_6_ns_1_10_cascade_ ));
    CascadeMux I__2704 (
            .O(N__22270),
            .I(\ALU.a_6_ns_1_11_cascade_ ));
    CascadeMux I__2703 (
            .O(N__22267),
            .I(\ALU.r6_RNIT7372Z0Z_11_cascade_ ));
    CascadeMux I__2702 (
            .O(N__22264),
            .I(\ALU.b_5_cascade_ ));
    CascadeMux I__2701 (
            .O(N__22261),
            .I(TXbuffer_18_3_ns_1_1_cascade_));
    CascadeMux I__2700 (
            .O(N__22258),
            .I(TXbuffer_RNO_5Z0Z_1_cascade_));
    InMux I__2699 (
            .O(N__22255),
            .I(N__22250));
    InMux I__2698 (
            .O(N__22254),
            .I(N__22245));
    InMux I__2697 (
            .O(N__22253),
            .I(N__22245));
    LocalMux I__2696 (
            .O(N__22250),
            .I(r6_9));
    LocalMux I__2695 (
            .O(N__22245),
            .I(r6_9));
    CascadeMux I__2694 (
            .O(N__22240),
            .I(TXbuffer_18_6_ns_1_1_cascade_));
    InMux I__2693 (
            .O(N__22237),
            .I(N__22234));
    LocalMux I__2692 (
            .O(N__22234),
            .I(TXbuffer_RNO_6Z0Z_1));
    InMux I__2691 (
            .O(N__22231),
            .I(N__22228));
    LocalMux I__2690 (
            .O(N__22228),
            .I(N__22221));
    InMux I__2689 (
            .O(N__22227),
            .I(N__22212));
    InMux I__2688 (
            .O(N__22226),
            .I(N__22212));
    InMux I__2687 (
            .O(N__22225),
            .I(N__22212));
    InMux I__2686 (
            .O(N__22224),
            .I(N__22212));
    Odrv4 I__2685 (
            .O(N__22221),
            .I(\ALU.madd_213 ));
    LocalMux I__2684 (
            .O(N__22212),
            .I(\ALU.madd_213 ));
    InMux I__2683 (
            .O(N__22207),
            .I(N__22202));
    InMux I__2682 (
            .O(N__22206),
            .I(N__22197));
    InMux I__2681 (
            .O(N__22205),
            .I(N__22197));
    LocalMux I__2680 (
            .O(N__22202),
            .I(N__22194));
    LocalMux I__2679 (
            .O(N__22197),
            .I(\ALU.a9_b_3 ));
    Odrv4 I__2678 (
            .O(N__22194),
            .I(\ALU.a9_b_3 ));
    InMux I__2677 (
            .O(N__22189),
            .I(N__22186));
    LocalMux I__2676 (
            .O(N__22186),
            .I(N__22183));
    Span4Mux_s1_h I__2675 (
            .O(N__22183),
            .I(N__22180));
    Span4Mux_v I__2674 (
            .O(N__22180),
            .I(N__22177));
    Odrv4 I__2673 (
            .O(N__22177),
            .I(\ALU.madd_167_0 ));
    CascadeMux I__2672 (
            .O(N__22174),
            .I(\ALU.b_6_ns_1_5_cascade_ ));
    CascadeMux I__2671 (
            .O(N__22171),
            .I(\ALU.b_3_ns_1_5_cascade_ ));
    InMux I__2670 (
            .O(N__22168),
            .I(N__22165));
    LocalMux I__2669 (
            .O(N__22165),
            .I(\ALU.r6_RNIBP2O1Z0Z_5 ));
    CascadeMux I__2668 (
            .O(N__22162),
            .I(\ALU.r4_RNI0QNE1Z0Z_5_cascade_ ));
    InMux I__2667 (
            .O(N__22159),
            .I(N__22154));
    InMux I__2666 (
            .O(N__22158),
            .I(N__22149));
    InMux I__2665 (
            .O(N__22157),
            .I(N__22149));
    LocalMux I__2664 (
            .O(N__22154),
            .I(N__22146));
    LocalMux I__2663 (
            .O(N__22149),
            .I(N__22143));
    Span4Mux_v I__2662 (
            .O(N__22146),
            .I(N__22138));
    Span4Mux_v I__2661 (
            .O(N__22143),
            .I(N__22138));
    Odrv4 I__2660 (
            .O(N__22138),
            .I(\ALU.a0_b_14 ));
    InMux I__2659 (
            .O(N__22135),
            .I(N__22132));
    LocalMux I__2658 (
            .O(N__22132),
            .I(\ALU.g2_0 ));
    InMux I__2657 (
            .O(N__22129),
            .I(N__22126));
    LocalMux I__2656 (
            .O(N__22126),
            .I(\ALU.g0_2_N_4L5 ));
    InMux I__2655 (
            .O(N__22123),
            .I(N__22117));
    InMux I__2654 (
            .O(N__22122),
            .I(N__22117));
    LocalMux I__2653 (
            .O(N__22117),
            .I(N__22114));
    Span4Mux_h I__2652 (
            .O(N__22114),
            .I(N__22110));
    InMux I__2651 (
            .O(N__22113),
            .I(N__22107));
    Odrv4 I__2650 (
            .O(N__22110),
            .I(\ALU.madd_134_0_tz ));
    LocalMux I__2649 (
            .O(N__22107),
            .I(\ALU.madd_134_0_tz ));
    InMux I__2648 (
            .O(N__22102),
            .I(N__22099));
    LocalMux I__2647 (
            .O(N__22099),
            .I(\ALU.madd_130_0 ));
    InMux I__2646 (
            .O(N__22096),
            .I(N__22093));
    LocalMux I__2645 (
            .O(N__22093),
            .I(N__22088));
    InMux I__2644 (
            .O(N__22092),
            .I(N__22083));
    InMux I__2643 (
            .O(N__22091),
            .I(N__22083));
    Span4Mux_s1_v I__2642 (
            .O(N__22088),
            .I(N__22080));
    LocalMux I__2641 (
            .O(N__22083),
            .I(N__22077));
    Span4Mux_h I__2640 (
            .O(N__22080),
            .I(N__22074));
    Span4Mux_s1_v I__2639 (
            .O(N__22077),
            .I(N__22071));
    Odrv4 I__2638 (
            .O(N__22074),
            .I(\ALU.madd_130 ));
    Odrv4 I__2637 (
            .O(N__22071),
            .I(\ALU.madd_130 ));
    CascadeMux I__2636 (
            .O(N__22066),
            .I(N__22063));
    InMux I__2635 (
            .O(N__22063),
            .I(N__22060));
    LocalMux I__2634 (
            .O(N__22060),
            .I(N__22057));
    Span4Mux_s1_h I__2633 (
            .O(N__22057),
            .I(N__22054));
    Odrv4 I__2632 (
            .O(N__22054),
            .I(\ALU.madd_171_sx ));
    InMux I__2631 (
            .O(N__22051),
            .I(N__22048));
    LocalMux I__2630 (
            .O(N__22048),
            .I(\ALU.a5_b_8 ));
    CascadeMux I__2629 (
            .O(N__22045),
            .I(N__22042));
    InMux I__2628 (
            .O(N__22042),
            .I(N__22036));
    InMux I__2627 (
            .O(N__22041),
            .I(N__22036));
    LocalMux I__2626 (
            .O(N__22036),
            .I(\ALU.a6_b_7 ));
    InMux I__2625 (
            .O(N__22033),
            .I(N__22029));
    InMux I__2624 (
            .O(N__22032),
            .I(N__22026));
    LocalMux I__2623 (
            .O(N__22029),
            .I(N__22021));
    LocalMux I__2622 (
            .O(N__22026),
            .I(N__22021));
    Odrv4 I__2621 (
            .O(N__22021),
            .I(\ALU.madd_321 ));
    CascadeMux I__2620 (
            .O(N__22018),
            .I(\ALU.b_6_ns_1_6_cascade_ ));
    CascadeMux I__2619 (
            .O(N__22015),
            .I(\ALU.r6_RNIIH042Z0Z_6_cascade_ ));
    CascadeMux I__2618 (
            .O(N__22012),
            .I(\ALU.b_6_cascade_ ));
    InMux I__2617 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__2616 (
            .O(N__22006),
            .I(N__22003));
    Odrv4 I__2615 (
            .O(N__22003),
            .I(\ALU.g0_2_N_3L3 ));
    CascadeMux I__2614 (
            .O(N__22000),
            .I(N__21996));
    InMux I__2613 (
            .O(N__21999),
            .I(N__21986));
    InMux I__2612 (
            .O(N__21996),
            .I(N__21986));
    CascadeMux I__2611 (
            .O(N__21995),
            .I(N__21981));
    CascadeMux I__2610 (
            .O(N__21994),
            .I(N__21976));
    InMux I__2609 (
            .O(N__21993),
            .I(N__21971));
    InMux I__2608 (
            .O(N__21992),
            .I(N__21971));
    CascadeMux I__2607 (
            .O(N__21991),
            .I(N__21965));
    LocalMux I__2606 (
            .O(N__21986),
            .I(N__21960));
    InMux I__2605 (
            .O(N__21985),
            .I(N__21947));
    InMux I__2604 (
            .O(N__21984),
            .I(N__21947));
    InMux I__2603 (
            .O(N__21981),
            .I(N__21947));
    InMux I__2602 (
            .O(N__21980),
            .I(N__21947));
    InMux I__2601 (
            .O(N__21979),
            .I(N__21947));
    InMux I__2600 (
            .O(N__21976),
            .I(N__21947));
    LocalMux I__2599 (
            .O(N__21971),
            .I(N__21944));
    InMux I__2598 (
            .O(N__21970),
            .I(N__21936));
    InMux I__2597 (
            .O(N__21969),
            .I(N__21936));
    InMux I__2596 (
            .O(N__21968),
            .I(N__21936));
    InMux I__2595 (
            .O(N__21965),
            .I(N__21929));
    InMux I__2594 (
            .O(N__21964),
            .I(N__21929));
    InMux I__2593 (
            .O(N__21963),
            .I(N__21926));
    Span4Mux_v I__2592 (
            .O(N__21960),
            .I(N__21921));
    LocalMux I__2591 (
            .O(N__21947),
            .I(N__21921));
    Span4Mux_v I__2590 (
            .O(N__21944),
            .I(N__21918));
    InMux I__2589 (
            .O(N__21943),
            .I(N__21915));
    LocalMux I__2588 (
            .O(N__21936),
            .I(N__21912));
    InMux I__2587 (
            .O(N__21935),
            .I(N__21907));
    InMux I__2586 (
            .O(N__21934),
            .I(N__21907));
    LocalMux I__2585 (
            .O(N__21929),
            .I(bZ0Z_2));
    LocalMux I__2584 (
            .O(N__21926),
            .I(bZ0Z_2));
    Odrv4 I__2583 (
            .O(N__21921),
            .I(bZ0Z_2));
    Odrv4 I__2582 (
            .O(N__21918),
            .I(bZ0Z_2));
    LocalMux I__2581 (
            .O(N__21915),
            .I(bZ0Z_2));
    Odrv4 I__2580 (
            .O(N__21912),
            .I(bZ0Z_2));
    LocalMux I__2579 (
            .O(N__21907),
            .I(bZ0Z_2));
    CascadeMux I__2578 (
            .O(N__21892),
            .I(\ALU.b_3_ns_1_6_cascade_ ));
    InMux I__2577 (
            .O(N__21889),
            .I(N__21886));
    LocalMux I__2576 (
            .O(N__21886),
            .I(\ALU.r4_RNIAP7R1Z0Z_6 ));
    InMux I__2575 (
            .O(N__21883),
            .I(N__21880));
    LocalMux I__2574 (
            .O(N__21880),
            .I(N__21877));
    Odrv4 I__2573 (
            .O(N__21877),
            .I(\ALU.madd_144_0_tz ));
    InMux I__2572 (
            .O(N__21874),
            .I(N__21868));
    InMux I__2571 (
            .O(N__21873),
            .I(N__21865));
    InMux I__2570 (
            .O(N__21872),
            .I(N__21860));
    InMux I__2569 (
            .O(N__21871),
            .I(N__21860));
    LocalMux I__2568 (
            .O(N__21868),
            .I(N__21857));
    LocalMux I__2567 (
            .O(N__21865),
            .I(\ALU.a4_b_5 ));
    LocalMux I__2566 (
            .O(N__21860),
            .I(\ALU.a4_b_5 ));
    Odrv4 I__2565 (
            .O(N__21857),
            .I(\ALU.a4_b_5 ));
    InMux I__2564 (
            .O(N__21850),
            .I(N__21847));
    LocalMux I__2563 (
            .O(N__21847),
            .I(N__21844));
    Span4Mux_s0_v I__2562 (
            .O(N__21844),
            .I(N__21841));
    Odrv4 I__2561 (
            .O(N__21841),
            .I(\ALU.g0_6_1 ));
    InMux I__2560 (
            .O(N__21838),
            .I(N__21835));
    LocalMux I__2559 (
            .O(N__21835),
            .I(N__21831));
    InMux I__2558 (
            .O(N__21834),
            .I(N__21828));
    Span4Mux_v I__2557 (
            .O(N__21831),
            .I(N__21825));
    LocalMux I__2556 (
            .O(N__21828),
            .I(N__21822));
    Odrv4 I__2555 (
            .O(N__21825),
            .I(\ALU.r6_RNIUC0U1Z0Z_10 ));
    Odrv4 I__2554 (
            .O(N__21822),
            .I(\ALU.r6_RNIUC0U1Z0Z_10 ));
    InMux I__2553 (
            .O(N__21817),
            .I(N__21814));
    LocalMux I__2552 (
            .O(N__21814),
            .I(N__21811));
    Span4Mux_v I__2551 (
            .O(N__21811),
            .I(N__21807));
    InMux I__2550 (
            .O(N__21810),
            .I(N__21804));
    Odrv4 I__2549 (
            .O(N__21807),
            .I(\ALU.r5_RNIMCFS1Z0Z_10 ));
    LocalMux I__2548 (
            .O(N__21804),
            .I(\ALU.r5_RNIMCFS1Z0Z_10 ));
    InMux I__2547 (
            .O(N__21799),
            .I(N__21796));
    LocalMux I__2546 (
            .O(N__21796),
            .I(\ALU.a0_b_10 ));
    CascadeMux I__2545 (
            .O(N__21793),
            .I(\ALU.a5_b_8_cascade_ ));
    InMux I__2544 (
            .O(N__21790),
            .I(N__21787));
    LocalMux I__2543 (
            .O(N__21787),
            .I(N__21783));
    InMux I__2542 (
            .O(N__21786),
            .I(N__21780));
    Span4Mux_v I__2541 (
            .O(N__21783),
            .I(N__21777));
    LocalMux I__2540 (
            .O(N__21780),
            .I(N__21774));
    Span4Mux_v I__2539 (
            .O(N__21777),
            .I(N__21771));
    Span4Mux_s3_h I__2538 (
            .O(N__21774),
            .I(N__21768));
    Odrv4 I__2537 (
            .O(N__21771),
            .I(\ALU.madd_325 ));
    Odrv4 I__2536 (
            .O(N__21768),
            .I(\ALU.madd_325 ));
    CascadeMux I__2535 (
            .O(N__21763),
            .I(\ALU.b_7_cascade_ ));
    CascadeMux I__2534 (
            .O(N__21760),
            .I(N__21756));
    InMux I__2533 (
            .O(N__21759),
            .I(N__21753));
    InMux I__2532 (
            .O(N__21756),
            .I(N__21750));
    LocalMux I__2531 (
            .O(N__21753),
            .I(\ALU.a5_b_7 ));
    LocalMux I__2530 (
            .O(N__21750),
            .I(\ALU.a5_b_7 ));
    CascadeMux I__2529 (
            .O(N__21745),
            .I(\ALU.a5_b_5_cascade_ ));
    InMux I__2528 (
            .O(N__21742),
            .I(N__21736));
    InMux I__2527 (
            .O(N__21741),
            .I(N__21736));
    LocalMux I__2526 (
            .O(N__21736),
            .I(N__21731));
    InMux I__2525 (
            .O(N__21735),
            .I(N__21726));
    InMux I__2524 (
            .O(N__21734),
            .I(N__21726));
    Span4Mux_s2_v I__2523 (
            .O(N__21731),
            .I(N__21721));
    LocalMux I__2522 (
            .O(N__21726),
            .I(N__21721));
    Odrv4 I__2521 (
            .O(N__21721),
            .I(\ALU.madd_176 ));
    CascadeMux I__2520 (
            .O(N__21718),
            .I(\ALU.madd_43_0_cascade_ ));
    InMux I__2519 (
            .O(N__21715),
            .I(N__21712));
    LocalMux I__2518 (
            .O(N__21712),
            .I(\ALU.madd_77_0_tz ));
    InMux I__2517 (
            .O(N__21709),
            .I(N__21705));
    InMux I__2516 (
            .O(N__21708),
            .I(N__21702));
    LocalMux I__2515 (
            .O(N__21705),
            .I(N__21699));
    LocalMux I__2514 (
            .O(N__21702),
            .I(N__21696));
    Odrv4 I__2513 (
            .O(N__21699),
            .I(\ALU.madd_278 ));
    Odrv4 I__2512 (
            .O(N__21696),
            .I(\ALU.madd_278 ));
    InMux I__2511 (
            .O(N__21691),
            .I(N__21688));
    LocalMux I__2510 (
            .O(N__21688),
            .I(N__21684));
    InMux I__2509 (
            .O(N__21687),
            .I(N__21681));
    Span4Mux_s3_h I__2508 (
            .O(N__21684),
            .I(N__21678));
    LocalMux I__2507 (
            .O(N__21681),
            .I(\ALU.madd_273 ));
    Odrv4 I__2506 (
            .O(N__21678),
            .I(\ALU.madd_273 ));
    CascadeMux I__2505 (
            .O(N__21673),
            .I(N__21669));
    InMux I__2504 (
            .O(N__21672),
            .I(N__21665));
    InMux I__2503 (
            .O(N__21669),
            .I(N__21662));
    InMux I__2502 (
            .O(N__21668),
            .I(N__21659));
    LocalMux I__2501 (
            .O(N__21665),
            .I(N__21656));
    LocalMux I__2500 (
            .O(N__21662),
            .I(N__21653));
    LocalMux I__2499 (
            .O(N__21659),
            .I(N__21650));
    Span4Mux_v I__2498 (
            .O(N__21656),
            .I(N__21647));
    Span4Mux_s3_h I__2497 (
            .O(N__21653),
            .I(N__21642));
    Span4Mux_s3_h I__2496 (
            .O(N__21650),
            .I(N__21642));
    Span4Mux_h I__2495 (
            .O(N__21647),
            .I(N__21639));
    Span4Mux_v I__2494 (
            .O(N__21642),
            .I(N__21636));
    Odrv4 I__2493 (
            .O(N__21639),
            .I(\ALU.madd_345 ));
    Odrv4 I__2492 (
            .O(N__21636),
            .I(\ALU.madd_345 ));
    InMux I__2491 (
            .O(N__21631),
            .I(N__21628));
    LocalMux I__2490 (
            .O(N__21628),
            .I(\ALU.madd_159_N_3L3 ));
    InMux I__2489 (
            .O(N__21625),
            .I(N__21622));
    LocalMux I__2488 (
            .O(N__21622),
            .I(\ALU.madd_61 ));
    CascadeMux I__2487 (
            .O(N__21619),
            .I(N__21616));
    InMux I__2486 (
            .O(N__21616),
            .I(N__21613));
    LocalMux I__2485 (
            .O(N__21613),
            .I(\ALU.madd_140_0 ));
    CascadeMux I__2484 (
            .O(N__21610),
            .I(\ALU.madd_140_0_cascade_ ));
    InMux I__2483 (
            .O(N__21607),
            .I(N__21604));
    LocalMux I__2482 (
            .O(N__21604),
            .I(\ALU.madd_155_1 ));
    InMux I__2481 (
            .O(N__21601),
            .I(N__21597));
    CascadeMux I__2480 (
            .O(N__21600),
            .I(N__21594));
    LocalMux I__2479 (
            .O(N__21597),
            .I(N__21591));
    InMux I__2478 (
            .O(N__21594),
            .I(N__21588));
    Odrv12 I__2477 (
            .O(N__21591),
            .I(\ALU.a_i_11 ));
    LocalMux I__2476 (
            .O(N__21588),
            .I(\ALU.a_i_11 ));
    InMux I__2475 (
            .O(N__21583),
            .I(N__21580));
    LocalMux I__2474 (
            .O(N__21580),
            .I(\ALU.r0_12_prm_3_11_s0_sf ));
    InMux I__2473 (
            .O(N__21577),
            .I(\ALU.r0_12_s0_11 ));
    InMux I__2472 (
            .O(N__21574),
            .I(N__21571));
    LocalMux I__2471 (
            .O(N__21571),
            .I(N__21568));
    Span4Mux_h I__2470 (
            .O(N__21568),
            .I(N__21565));
    Odrv4 I__2469 (
            .O(N__21565),
            .I(\ALU.r0_12_s0_11_THRU_CO ));
    CascadeMux I__2468 (
            .O(N__21562),
            .I(\ALU.g1_7_cascade_ ));
    InMux I__2467 (
            .O(N__21559),
            .I(N__21556));
    LocalMux I__2466 (
            .O(N__21556),
            .I(\ALU.a4_b_0_0_5 ));
    CascadeMux I__2465 (
            .O(N__21553),
            .I(\ALU.N_663_0_cascade_ ));
    InMux I__2464 (
            .O(N__21550),
            .I(N__21543));
    InMux I__2463 (
            .O(N__21549),
            .I(N__21543));
    InMux I__2462 (
            .O(N__21548),
            .I(N__21540));
    LocalMux I__2461 (
            .O(N__21543),
            .I(\ALU.madd_109 ));
    LocalMux I__2460 (
            .O(N__21540),
            .I(\ALU.madd_109 ));
    InMux I__2459 (
            .O(N__21535),
            .I(N__21532));
    LocalMux I__2458 (
            .O(N__21532),
            .I(N__21529));
    Odrv4 I__2457 (
            .O(N__21529),
            .I(\ALU.N_683_0_0_0 ));
    CascadeMux I__2456 (
            .O(N__21526),
            .I(TXbuffer_18_6_ns_1_0_cascade_));
    InMux I__2455 (
            .O(N__21523),
            .I(N__21520));
    LocalMux I__2454 (
            .O(N__21520),
            .I(N__21517));
    Span4Mux_s2_h I__2453 (
            .O(N__21517),
            .I(N__21514));
    Odrv4 I__2452 (
            .O(N__21514),
            .I(TXbuffer_RNO_6Z0Z_0));
    InMux I__2451 (
            .O(N__21511),
            .I(N__21508));
    LocalMux I__2450 (
            .O(N__21508),
            .I(N__21505));
    Span4Mux_v I__2449 (
            .O(N__21505),
            .I(N__21502));
    Odrv4 I__2448 (
            .O(N__21502),
            .I(TXbuffer_18_13_ns_1_7));
    InMux I__2447 (
            .O(N__21499),
            .I(N__21495));
    InMux I__2446 (
            .O(N__21498),
            .I(N__21492));
    LocalMux I__2445 (
            .O(N__21495),
            .I(N__21489));
    LocalMux I__2444 (
            .O(N__21492),
            .I(N__21486));
    Span4Mux_h I__2443 (
            .O(N__21489),
            .I(N__21483));
    Odrv4 I__2442 (
            .O(N__21486),
            .I(\ALU.r5_RNIE0AK8_0Z0Z_11 ));
    Odrv4 I__2441 (
            .O(N__21483),
            .I(\ALU.r5_RNIE0AK8_0Z0Z_11 ));
    CascadeMux I__2440 (
            .O(N__21478),
            .I(N__21475));
    InMux I__2439 (
            .O(N__21475),
            .I(N__21472));
    LocalMux I__2438 (
            .O(N__21472),
            .I(N__21468));
    InMux I__2437 (
            .O(N__21471),
            .I(N__21465));
    Span4Mux_v I__2436 (
            .O(N__21468),
            .I(N__21462));
    LocalMux I__2435 (
            .O(N__21465),
            .I(\ALU.r5_RNIE0AK8_1Z0Z_11 ));
    Odrv4 I__2434 (
            .O(N__21462),
            .I(\ALU.r5_RNIE0AK8_1Z0Z_11 ));
    CascadeMux I__2433 (
            .O(N__21457),
            .I(\ALU.b_6_ns_1_12_cascade_ ));
    InMux I__2432 (
            .O(N__21454),
            .I(N__21451));
    LocalMux I__2431 (
            .O(N__21451),
            .I(N__21448));
    Odrv12 I__2430 (
            .O(N__21448),
            .I(\ALU.r6_RNI85GA2Z0Z_12 ));
    InMux I__2429 (
            .O(N__21445),
            .I(N__21442));
    LocalMux I__2428 (
            .O(N__21442),
            .I(N__21439));
    Span4Mux_v I__2427 (
            .O(N__21439),
            .I(N__21435));
    InMux I__2426 (
            .O(N__21438),
            .I(N__21432));
    Odrv4 I__2425 (
            .O(N__21435),
            .I(\ALU.r5_RNI05V82Z0Z_12 ));
    LocalMux I__2424 (
            .O(N__21432),
            .I(\ALU.r5_RNI05V82Z0Z_12 ));
    CascadeMux I__2423 (
            .O(N__21427),
            .I(\ALU.r6_RNI85GA2Z0Z_12_cascade_ ));
    CascadeMux I__2422 (
            .O(N__21424),
            .I(\ALU.b_3_ns_1_13_cascade_ ));
    InMux I__2421 (
            .O(N__21421),
            .I(N__21418));
    LocalMux I__2420 (
            .O(N__21418),
            .I(\ALU.r5_RNI49V82Z0Z_13 ));
    CascadeMux I__2419 (
            .O(N__21415),
            .I(\ALU.a_6_ns_1_15_cascade_ ));
    InMux I__2418 (
            .O(N__21412),
            .I(N__21409));
    LocalMux I__2417 (
            .O(N__21409),
            .I(\ALU.r6_RNIH8772Z0Z_15 ));
    InMux I__2416 (
            .O(N__21406),
            .I(N__21403));
    LocalMux I__2415 (
            .O(N__21403),
            .I(N__21400));
    Span4Mux_s3_h I__2414 (
            .O(N__21400),
            .I(N__21397));
    Odrv4 I__2413 (
            .O(N__21397),
            .I(\ALU.r6_RNINRNUZ0Z_15 ));
    CascadeMux I__2412 (
            .O(N__21394),
            .I(N__21391));
    InMux I__2411 (
            .O(N__21391),
            .I(N__21388));
    LocalMux I__2410 (
            .O(N__21388),
            .I(\ALU.r0_12_prm_1_11_s1_c_RNOZ0 ));
    InMux I__2409 (
            .O(N__21385),
            .I(\ALU.r0_12_s1_11 ));
    CascadeMux I__2408 (
            .O(N__21382),
            .I(\ALU.b_3_ns_1_12_cascade_ ));
    InMux I__2407 (
            .O(N__21379),
            .I(N__21376));
    LocalMux I__2406 (
            .O(N__21376),
            .I(\ALU.r5_RNIH9VTZ0Z_14 ));
    CascadeMux I__2405 (
            .O(N__21373),
            .I(\ALU.r1_RNI8DSRZ0Z_14_cascade_ ));
    InMux I__2404 (
            .O(N__21370),
            .I(N__21367));
    LocalMux I__2403 (
            .O(N__21367),
            .I(\ALU.r2_RNIDP6TZ0Z_14 ));
    CascadeMux I__2402 (
            .O(N__21364),
            .I(\ALU.b_7_ns_1_14_cascade_ ));
    InMux I__2401 (
            .O(N__21361),
            .I(N__21358));
    LocalMux I__2400 (
            .O(N__21358),
            .I(\ALU.r6_RNILPNUZ0Z_14 ));
    CascadeMux I__2399 (
            .O(N__21355),
            .I(\ALU.b_14_cascade_ ));
    CascadeMux I__2398 (
            .O(N__21352),
            .I(N__21349));
    InMux I__2397 (
            .O(N__21349),
            .I(N__21346));
    LocalMux I__2396 (
            .O(N__21346),
            .I(N__21343));
    Odrv4 I__2395 (
            .O(N__21343),
            .I(\ALU.r0_12_prm_7_11_s1_c_RNOZ0 ));
    CascadeMux I__2394 (
            .O(N__21340),
            .I(N__21337));
    InMux I__2393 (
            .O(N__21337),
            .I(N__21334));
    LocalMux I__2392 (
            .O(N__21334),
            .I(N__21331));
    Odrv4 I__2391 (
            .O(N__21331),
            .I(\ALU.r0_12_prm_5_11_s1_c_RNOZ0 ));
    CascadeMux I__2390 (
            .O(N__21328),
            .I(\ALU.b_6_ns_1_11_cascade_ ));
    InMux I__2389 (
            .O(N__21325),
            .I(N__21322));
    LocalMux I__2388 (
            .O(N__21322),
            .I(N__21319));
    Odrv4 I__2387 (
            .O(N__21319),
            .I(\ALU.r6_RNI2H0U1Z0Z_11 ));
    CascadeMux I__2386 (
            .O(N__21316),
            .I(\ALU.b_6_ns_1_9_cascade_ ));
    InMux I__2385 (
            .O(N__21313),
            .I(N__21310));
    LocalMux I__2384 (
            .O(N__21310),
            .I(N__21307));
    Span4Mux_v I__2383 (
            .O(N__21307),
            .I(N__21303));
    InMux I__2382 (
            .O(N__21306),
            .I(N__21300));
    Odrv4 I__2381 (
            .O(N__21303),
            .I(\ALU.r6_RNIUT042Z0Z_9 ));
    LocalMux I__2380 (
            .O(N__21300),
            .I(\ALU.r6_RNIUT042Z0Z_9 ));
    CascadeMux I__2379 (
            .O(N__21295),
            .I(\ALU.b_3_ns_1_9_cascade_ ));
    InMux I__2378 (
            .O(N__21292),
            .I(N__21289));
    LocalMux I__2377 (
            .O(N__21289),
            .I(N__21285));
    InMux I__2376 (
            .O(N__21288),
            .I(N__21282));
    Odrv12 I__2375 (
            .O(N__21285),
            .I(\ALU.r4_RNIM58R1Z0Z_9 ));
    LocalMux I__2374 (
            .O(N__21282),
            .I(\ALU.r4_RNIM58R1Z0Z_9 ));
    CascadeMux I__2373 (
            .O(N__21277),
            .I(\ALU.b_3_ns_1_10_cascade_ ));
    CascadeMux I__2372 (
            .O(N__21274),
            .I(\ALU.b_3_ns_1_11_cascade_ ));
    CascadeMux I__2371 (
            .O(N__21271),
            .I(\ALU.r5_RNIQGFS1Z0Z_11_cascade_ ));
    CascadeMux I__2370 (
            .O(N__21268),
            .I(\ALU.b_6_ns_1_10_cascade_ ));
    CascadeMux I__2369 (
            .O(N__21265),
            .I(\ALU.a12_b_0_cascade_ ));
    InMux I__2368 (
            .O(N__21262),
            .I(N__21258));
    InMux I__2367 (
            .O(N__21261),
            .I(N__21255));
    LocalMux I__2366 (
            .O(N__21258),
            .I(N__21250));
    LocalMux I__2365 (
            .O(N__21255),
            .I(N__21250));
    Odrv4 I__2364 (
            .O(N__21250),
            .I(\ALU.madd_263 ));
    CascadeMux I__2363 (
            .O(N__21247),
            .I(\ALU.madd_264_cascade_ ));
    InMux I__2362 (
            .O(N__21244),
            .I(N__21238));
    InMux I__2361 (
            .O(N__21243),
            .I(N__21238));
    LocalMux I__2360 (
            .O(N__21238),
            .I(\ALU.madd_288 ));
    InMux I__2359 (
            .O(N__21235),
            .I(N__21232));
    LocalMux I__2358 (
            .O(N__21232),
            .I(\ALU.a12_b_0 ));
    CascadeMux I__2357 (
            .O(N__21229),
            .I(N__21225));
    InMux I__2356 (
            .O(N__21228),
            .I(N__21220));
    InMux I__2355 (
            .O(N__21225),
            .I(N__21220));
    LocalMux I__2354 (
            .O(N__21220),
            .I(\ALU.a10_b_2 ));
    InMux I__2353 (
            .O(N__21217),
            .I(N__21214));
    LocalMux I__2352 (
            .O(N__21214),
            .I(\ALU.madd_259 ));
    CascadeMux I__2351 (
            .O(N__21211),
            .I(N__21207));
    InMux I__2350 (
            .O(N__21210),
            .I(N__21203));
    InMux I__2349 (
            .O(N__21207),
            .I(N__21198));
    InMux I__2348 (
            .O(N__21206),
            .I(N__21198));
    LocalMux I__2347 (
            .O(N__21203),
            .I(N__21195));
    LocalMux I__2346 (
            .O(N__21198),
            .I(\ALU.a7_b_5 ));
    Odrv4 I__2345 (
            .O(N__21195),
            .I(\ALU.a7_b_5 ));
    CascadeMux I__2344 (
            .O(N__21190),
            .I(\ALU.madd_259_cascade_ ));
    CascadeMux I__2343 (
            .O(N__21187),
            .I(N__21184));
    InMux I__2342 (
            .O(N__21184),
            .I(N__21180));
    InMux I__2341 (
            .O(N__21183),
            .I(N__21177));
    LocalMux I__2340 (
            .O(N__21180),
            .I(N__21174));
    LocalMux I__2339 (
            .O(N__21177),
            .I(N__21171));
    Span4Mux_s2_h I__2338 (
            .O(N__21174),
            .I(N__21166));
    Span4Mux_s3_v I__2337 (
            .O(N__21171),
            .I(N__21166));
    Odrv4 I__2336 (
            .O(N__21166),
            .I(\ALU.madd_284_0 ));
    InMux I__2335 (
            .O(N__21163),
            .I(N__21154));
    InMux I__2334 (
            .O(N__21162),
            .I(N__21154));
    InMux I__2333 (
            .O(N__21161),
            .I(N__21154));
    LocalMux I__2332 (
            .O(N__21154),
            .I(\ALU.madd_336 ));
    CascadeMux I__2331 (
            .O(N__21151),
            .I(N__21147));
    CascadeMux I__2330 (
            .O(N__21150),
            .I(N__21144));
    InMux I__2329 (
            .O(N__21147),
            .I(N__21136));
    InMux I__2328 (
            .O(N__21144),
            .I(N__21136));
    InMux I__2327 (
            .O(N__21143),
            .I(N__21136));
    LocalMux I__2326 (
            .O(N__21136),
            .I(N__21133));
    Odrv4 I__2325 (
            .O(N__21133),
            .I(\ALU.madd_335 ));
    InMux I__2324 (
            .O(N__21130),
            .I(N__21127));
    LocalMux I__2323 (
            .O(N__21127),
            .I(\ALU.madd_283 ));
    InMux I__2322 (
            .O(N__21124),
            .I(N__21121));
    LocalMux I__2321 (
            .O(N__21121),
            .I(N__21118));
    Odrv4 I__2320 (
            .O(N__21118),
            .I(\ALU.madd_124_0 ));
    CascadeMux I__2319 (
            .O(N__21115),
            .I(N__21112));
    InMux I__2318 (
            .O(N__21112),
            .I(N__21109));
    LocalMux I__2317 (
            .O(N__21109),
            .I(N__21106));
    Odrv4 I__2316 (
            .O(N__21106),
            .I(\ALU.madd_218_0_tz ));
    CascadeMux I__2315 (
            .O(N__21103),
            .I(\ALU.madd_218_cascade_ ));
    InMux I__2314 (
            .O(N__21100),
            .I(N__21097));
    LocalMux I__2313 (
            .O(N__21097),
            .I(\ALU.madd_346_1 ));
    InMux I__2312 (
            .O(N__21094),
            .I(N__21088));
    InMux I__2311 (
            .O(N__21093),
            .I(N__21088));
    LocalMux I__2310 (
            .O(N__21088),
            .I(N__21085));
    Odrv4 I__2309 (
            .O(N__21085),
            .I(\ALU.a2_b_10 ));
    CascadeMux I__2308 (
            .O(N__21082),
            .I(\ALU.a0_b_12_cascade_ ));
    InMux I__2307 (
            .O(N__21079),
            .I(N__21075));
    InMux I__2306 (
            .O(N__21078),
            .I(N__21072));
    LocalMux I__2305 (
            .O(N__21075),
            .I(N__21069));
    LocalMux I__2304 (
            .O(N__21072),
            .I(\ALU.madd_279_0 ));
    Odrv4 I__2303 (
            .O(N__21069),
            .I(\ALU.madd_279_0 ));
    InMux I__2302 (
            .O(N__21064),
            .I(N__21060));
    InMux I__2301 (
            .O(N__21063),
            .I(N__21056));
    LocalMux I__2300 (
            .O(N__21060),
            .I(N__21053));
    InMux I__2299 (
            .O(N__21059),
            .I(N__21050));
    LocalMux I__2298 (
            .O(N__21056),
            .I(\ALU.madd_331_0 ));
    Odrv12 I__2297 (
            .O(N__21053),
            .I(\ALU.madd_331_0 ));
    LocalMux I__2296 (
            .O(N__21050),
            .I(\ALU.madd_331_0 ));
    CascadeMux I__2295 (
            .O(N__21043),
            .I(N__21040));
    InMux I__2294 (
            .O(N__21040),
            .I(N__21037));
    LocalMux I__2293 (
            .O(N__21037),
            .I(N__21033));
    CascadeMux I__2292 (
            .O(N__21036),
            .I(N__21030));
    Span4Mux_s2_h I__2291 (
            .O(N__21033),
            .I(N__21025));
    InMux I__2290 (
            .O(N__21030),
            .I(N__21022));
    InMux I__2289 (
            .O(N__21029),
            .I(N__21017));
    InMux I__2288 (
            .O(N__21028),
            .I(N__21017));
    Odrv4 I__2287 (
            .O(N__21025),
            .I(\ALU.a0_b_12 ));
    LocalMux I__2286 (
            .O(N__21022),
            .I(\ALU.a0_b_12 ));
    LocalMux I__2285 (
            .O(N__21017),
            .I(\ALU.a0_b_12 ));
    InMux I__2284 (
            .O(N__21010),
            .I(N__21003));
    InMux I__2283 (
            .O(N__21009),
            .I(N__21003));
    InMux I__2282 (
            .O(N__21008),
            .I(N__20998));
    LocalMux I__2281 (
            .O(N__21003),
            .I(N__20995));
    InMux I__2280 (
            .O(N__21002),
            .I(N__20990));
    InMux I__2279 (
            .O(N__21001),
            .I(N__20990));
    LocalMux I__2278 (
            .O(N__20998),
            .I(\ALU.madd_218 ));
    Odrv12 I__2277 (
            .O(N__20995),
            .I(\ALU.madd_218 ));
    LocalMux I__2276 (
            .O(N__20990),
            .I(\ALU.madd_218 ));
    InMux I__2275 (
            .O(N__20983),
            .I(N__20979));
    InMux I__2274 (
            .O(N__20982),
            .I(N__20976));
    LocalMux I__2273 (
            .O(N__20979),
            .I(\ALU.madd_202 ));
    LocalMux I__2272 (
            .O(N__20976),
            .I(\ALU.madd_202 ));
    InMux I__2271 (
            .O(N__20971),
            .I(N__20967));
    InMux I__2270 (
            .O(N__20970),
            .I(N__20964));
    LocalMux I__2269 (
            .O(N__20967),
            .I(\ALU.madd_228 ));
    LocalMux I__2268 (
            .O(N__20964),
            .I(\ALU.madd_228 ));
    InMux I__2267 (
            .O(N__20959),
            .I(N__20956));
    LocalMux I__2266 (
            .O(N__20956),
            .I(N__20952));
    InMux I__2265 (
            .O(N__20955),
            .I(N__20949));
    Odrv12 I__2264 (
            .O(N__20952),
            .I(\ALU.madd_338 ));
    LocalMux I__2263 (
            .O(N__20949),
            .I(\ALU.madd_338 ));
    InMux I__2262 (
            .O(N__20944),
            .I(N__20941));
    LocalMux I__2261 (
            .O(N__20941),
            .I(N__20937));
    InMux I__2260 (
            .O(N__20940),
            .I(N__20934));
    Odrv12 I__2259 (
            .O(N__20937),
            .I(\ALU.madd_337 ));
    LocalMux I__2258 (
            .O(N__20934),
            .I(\ALU.madd_337 ));
    InMux I__2257 (
            .O(N__20929),
            .I(N__20926));
    LocalMux I__2256 (
            .O(N__20926),
            .I(\ALU.a0_b_13 ));
    InMux I__2255 (
            .O(N__20923),
            .I(N__20919));
    InMux I__2254 (
            .O(N__20922),
            .I(N__20916));
    LocalMux I__2253 (
            .O(N__20919),
            .I(\ALU.madd_335_0 ));
    LocalMux I__2252 (
            .O(N__20916),
            .I(\ALU.madd_335_0 ));
    InMux I__2251 (
            .O(N__20911),
            .I(N__20908));
    LocalMux I__2250 (
            .O(N__20908),
            .I(N__20904));
    InMux I__2249 (
            .O(N__20907),
            .I(N__20901));
    Odrv4 I__2248 (
            .O(N__20904),
            .I(\ALU.madd_233 ));
    LocalMux I__2247 (
            .O(N__20901),
            .I(\ALU.madd_233 ));
    CascadeMux I__2246 (
            .O(N__20896),
            .I(N__20893));
    InMux I__2245 (
            .O(N__20893),
            .I(N__20889));
    CascadeMux I__2244 (
            .O(N__20892),
            .I(N__20886));
    LocalMux I__2243 (
            .O(N__20889),
            .I(N__20882));
    InMux I__2242 (
            .O(N__20886),
            .I(N__20877));
    InMux I__2241 (
            .O(N__20885),
            .I(N__20877));
    Span4Mux_h I__2240 (
            .O(N__20882),
            .I(N__20874));
    LocalMux I__2239 (
            .O(N__20877),
            .I(N__20871));
    Odrv4 I__2238 (
            .O(N__20874),
            .I(\ALU.madd_238 ));
    Odrv4 I__2237 (
            .O(N__20871),
            .I(\ALU.madd_238 ));
    InMux I__2236 (
            .O(N__20866),
            .I(N__20860));
    InMux I__2235 (
            .O(N__20865),
            .I(N__20860));
    LocalMux I__2234 (
            .O(N__20860),
            .I(\ALU.madd_294 ));
    InMux I__2233 (
            .O(N__20857),
            .I(N__20852));
    InMux I__2232 (
            .O(N__20856),
            .I(N__20849));
    InMux I__2231 (
            .O(N__20855),
            .I(N__20846));
    LocalMux I__2230 (
            .O(N__20852),
            .I(\ALU.madd_304 ));
    LocalMux I__2229 (
            .O(N__20849),
            .I(\ALU.madd_304 ));
    LocalMux I__2228 (
            .O(N__20846),
            .I(\ALU.madd_304 ));
    InMux I__2227 (
            .O(N__20839),
            .I(N__20833));
    InMux I__2226 (
            .O(N__20838),
            .I(N__20833));
    LocalMux I__2225 (
            .O(N__20833),
            .I(N__20829));
    InMux I__2224 (
            .O(N__20832),
            .I(N__20826));
    Odrv4 I__2223 (
            .O(N__20829),
            .I(\ALU.madd_253 ));
    LocalMux I__2222 (
            .O(N__20826),
            .I(\ALU.madd_253 ));
    InMux I__2221 (
            .O(N__20821),
            .I(N__20817));
    CascadeMux I__2220 (
            .O(N__20820),
            .I(N__20814));
    LocalMux I__2219 (
            .O(N__20817),
            .I(N__20811));
    InMux I__2218 (
            .O(N__20814),
            .I(N__20808));
    Odrv4 I__2217 (
            .O(N__20811),
            .I(\ALU.madd_341 ));
    LocalMux I__2216 (
            .O(N__20808),
            .I(\ALU.madd_341 ));
    InMux I__2215 (
            .O(N__20803),
            .I(N__20800));
    LocalMux I__2214 (
            .O(N__20800),
            .I(\ALU.a4_b_8 ));
    CascadeMux I__2213 (
            .O(N__20797),
            .I(\ALU.a4_b_8_cascade_ ));
    InMux I__2212 (
            .O(N__20794),
            .I(N__20791));
    LocalMux I__2211 (
            .O(N__20791),
            .I(\ALU.madd_269 ));
    CascadeMux I__2210 (
            .O(N__20788),
            .I(N__20784));
    InMux I__2209 (
            .O(N__20787),
            .I(N__20781));
    InMux I__2208 (
            .O(N__20784),
            .I(N__20778));
    LocalMux I__2207 (
            .O(N__20781),
            .I(\ALU.madd_274 ));
    LocalMux I__2206 (
            .O(N__20778),
            .I(\ALU.madd_274 ));
    CascadeMux I__2205 (
            .O(N__20773),
            .I(\ALU.madd_269_cascade_ ));
    InMux I__2204 (
            .O(N__20770),
            .I(N__20765));
    InMux I__2203 (
            .O(N__20769),
            .I(N__20760));
    InMux I__2202 (
            .O(N__20768),
            .I(N__20760));
    LocalMux I__2201 (
            .O(N__20765),
            .I(N__20757));
    LocalMux I__2200 (
            .O(N__20760),
            .I(\ALU.madd_289 ));
    Odrv4 I__2199 (
            .O(N__20757),
            .I(\ALU.madd_289 ));
    CascadeMux I__2198 (
            .O(N__20752),
            .I(\ALU.madd_185_1_cascade_ ));
    InMux I__2197 (
            .O(N__20749),
            .I(N__20743));
    InMux I__2196 (
            .O(N__20748),
            .I(N__20743));
    LocalMux I__2195 (
            .O(N__20743),
            .I(N__20740));
    Odrv4 I__2194 (
            .O(N__20740),
            .I(\ALU.madd_106 ));
    CascadeMux I__2193 (
            .O(N__20737),
            .I(\ALU.g0_2_N_2L1_cascade_ ));
    CascadeMux I__2192 (
            .O(N__20734),
            .I(N__20731));
    InMux I__2191 (
            .O(N__20731),
            .I(N__20725));
    InMux I__2190 (
            .O(N__20730),
            .I(N__20725));
    LocalMux I__2189 (
            .O(N__20725),
            .I(\ALU.madd_186_0 ));
    CascadeMux I__2188 (
            .O(N__20722),
            .I(N__20719));
    InMux I__2187 (
            .O(N__20719),
            .I(N__20715));
    InMux I__2186 (
            .O(N__20718),
            .I(N__20712));
    LocalMux I__2185 (
            .O(N__20715),
            .I(\ALU.a6_b_2 ));
    LocalMux I__2184 (
            .O(N__20712),
            .I(\ALU.a6_b_2 ));
    CascadeMux I__2183 (
            .O(N__20707),
            .I(\ALU.a6_b_2_cascade_ ));
    InMux I__2182 (
            .O(N__20704),
            .I(N__20700));
    InMux I__2181 (
            .O(N__20703),
            .I(N__20697));
    LocalMux I__2180 (
            .O(N__20700),
            .I(\ALU.a7_b_1 ));
    LocalMux I__2179 (
            .O(N__20697),
            .I(\ALU.a7_b_1 ));
    CascadeMux I__2178 (
            .O(N__20692),
            .I(\ALU.madd_99_cascade_ ));
    InMux I__2177 (
            .O(N__20689),
            .I(N__20681));
    InMux I__2176 (
            .O(N__20688),
            .I(N__20681));
    InMux I__2175 (
            .O(N__20687),
            .I(N__20676));
    InMux I__2174 (
            .O(N__20686),
            .I(N__20676));
    LocalMux I__2173 (
            .O(N__20681),
            .I(\ALU.madd_149 ));
    LocalMux I__2172 (
            .O(N__20676),
            .I(\ALU.madd_149 ));
    InMux I__2171 (
            .O(N__20671),
            .I(N__20668));
    LocalMux I__2170 (
            .O(N__20668),
            .I(\ALU.madd_99 ));
    InMux I__2169 (
            .O(N__20665),
            .I(N__20659));
    InMux I__2168 (
            .O(N__20664),
            .I(N__20659));
    LocalMux I__2167 (
            .O(N__20659),
            .I(\ALU.madd_145 ));
    InMux I__2166 (
            .O(N__20656),
            .I(N__20653));
    LocalMux I__2165 (
            .O(N__20653),
            .I(\ALU.madd_244 ));
    CascadeMux I__2164 (
            .O(N__20650),
            .I(N__20647));
    InMux I__2163 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__2162 (
            .O(N__20644),
            .I(\ALU.madd_201 ));
    InMux I__2161 (
            .O(N__20641),
            .I(N__20636));
    InMux I__2160 (
            .O(N__20640),
            .I(N__20633));
    InMux I__2159 (
            .O(N__20639),
            .I(N__20630));
    LocalMux I__2158 (
            .O(N__20636),
            .I(N__20627));
    LocalMux I__2157 (
            .O(N__20633),
            .I(\ALU.madd_239 ));
    LocalMux I__2156 (
            .O(N__20630),
            .I(\ALU.madd_239 ));
    Odrv4 I__2155 (
            .O(N__20627),
            .I(\ALU.madd_239 ));
    CascadeMux I__2154 (
            .O(N__20620),
            .I(\ALU.a3_b_9_cascade_ ));
    InMux I__2153 (
            .O(N__20617),
            .I(N__20614));
    LocalMux I__2152 (
            .O(N__20614),
            .I(\ALU.a3_b_9 ));
    CascadeMux I__2151 (
            .O(N__20611),
            .I(\ALU.madd_155_cascade_ ));
    CascadeMux I__2150 (
            .O(N__20608),
            .I(\ALU.madd_109_0_tz_cascade_ ));
    CascadeMux I__2149 (
            .O(N__20605),
            .I(\ALU.madd_109_cascade_ ));
    InMux I__2148 (
            .O(N__20602),
            .I(N__20599));
    LocalMux I__2147 (
            .O(N__20599),
            .I(\ALU.N_687_0 ));
    InMux I__2146 (
            .O(N__20596),
            .I(N__20593));
    LocalMux I__2145 (
            .O(N__20593),
            .I(N__20590));
    Span4Mux_s0_v I__2144 (
            .O(N__20590),
            .I(N__20587));
    Odrv4 I__2143 (
            .O(N__20587),
            .I(\ALU.madd_159_N_2L1 ));
    CascadeMux I__2142 (
            .O(N__20584),
            .I(N__20581));
    InMux I__2141 (
            .O(N__20581),
            .I(N__20575));
    InMux I__2140 (
            .O(N__20580),
            .I(N__20575));
    LocalMux I__2139 (
            .O(N__20575),
            .I(\ALU.madd_159 ));
    CascadeMux I__2138 (
            .O(N__20572),
            .I(N__20569));
    InMux I__2137 (
            .O(N__20569),
            .I(N__20563));
    InMux I__2136 (
            .O(N__20568),
            .I(N__20563));
    LocalMux I__2135 (
            .O(N__20563),
            .I(N__20560));
    Odrv4 I__2134 (
            .O(N__20560),
            .I(\ALU.madd_150 ));
    InMux I__2133 (
            .O(N__20557),
            .I(N__20551));
    InMux I__2132 (
            .O(N__20556),
            .I(N__20551));
    LocalMux I__2131 (
            .O(N__20551),
            .I(\ALU.madd_155 ));
    CascadeMux I__2130 (
            .O(N__20548),
            .I(\ALU.a7_b_1_cascade_ ));
    CascadeMux I__2129 (
            .O(N__20545),
            .I(\ALU.r6_RNIC9GA2Z0Z_13_cascade_ ));
    CascadeMux I__2128 (
            .O(N__20542),
            .I(\ALU.b_13_cascade_ ));
    CascadeMux I__2127 (
            .O(N__20539),
            .I(TXbuffer_18_13_ns_1_4_cascade_));
    InMux I__2126 (
            .O(N__20536),
            .I(N__20533));
    LocalMux I__2125 (
            .O(N__20533),
            .I(N__20530));
    Span4Mux_v I__2124 (
            .O(N__20530),
            .I(N__20527));
    Odrv4 I__2123 (
            .O(N__20527),
            .I(TXbuffer_RNO_1Z0Z_4));
    CascadeMux I__2122 (
            .O(N__20524),
            .I(N__20521));
    InMux I__2121 (
            .O(N__20521),
            .I(N__20518));
    LocalMux I__2120 (
            .O(N__20518),
            .I(N__20515));
    Odrv12 I__2119 (
            .O(N__20515),
            .I(\ALU.N_661_0 ));
    CascadeMux I__2118 (
            .O(N__20512),
            .I(\ALU.a_15_cascade_ ));
    CascadeMux I__2117 (
            .O(N__20509),
            .I(\ALU.lshift_3_ns_1_15_cascade_ ));
    CascadeMux I__2116 (
            .O(N__20506),
            .I(\ALU.b_6_ns_1_13_cascade_ ));
    InMux I__2115 (
            .O(N__20503),
            .I(N__20500));
    LocalMux I__2114 (
            .O(N__20500),
            .I(N__20497));
    Odrv4 I__2113 (
            .O(N__20497),
            .I(TXbuffer_18_13_ns_1_3));
    InMux I__2112 (
            .O(N__20494),
            .I(N__20491));
    LocalMux I__2111 (
            .O(N__20491),
            .I(\ALU.r1_RNIAFSRZ0Z_15 ));
    CascadeMux I__2110 (
            .O(N__20488),
            .I(\ALU.r5_RNIJBVTZ0Z_15_cascade_ ));
    InMux I__2109 (
            .O(N__20485),
            .I(N__20482));
    LocalMux I__2108 (
            .O(N__20482),
            .I(\ALU.b_7_ns_1_15 ));
    InMux I__2107 (
            .O(N__20479),
            .I(N__20476));
    LocalMux I__2106 (
            .O(N__20476),
            .I(N__20473));
    Span4Mux_v I__2105 (
            .O(N__20473),
            .I(N__20470));
    Span4Mux_v I__2104 (
            .O(N__20470),
            .I(N__20467));
    Odrv4 I__2103 (
            .O(N__20467),
            .I(\ALU.madd_490_1 ));
    InMux I__2102 (
            .O(N__20464),
            .I(N__20461));
    LocalMux I__2101 (
            .O(N__20461),
            .I(N__20458));
    Span4Mux_v I__2100 (
            .O(N__20458),
            .I(N__20455));
    Span4Mux_s1_h I__2099 (
            .O(N__20455),
            .I(N__20452));
    Odrv4 I__2098 (
            .O(N__20452),
            .I(\ALU.madd_490_9 ));
    CascadeMux I__2097 (
            .O(N__20449),
            .I(\ALU.madd_490_0_cascade_ ));
    InMux I__2096 (
            .O(N__20446),
            .I(N__20443));
    LocalMux I__2095 (
            .O(N__20443),
            .I(\ALU.madd_490_13 ));
    InMux I__2094 (
            .O(N__20440),
            .I(N__20437));
    LocalMux I__2093 (
            .O(N__20437),
            .I(N__20434));
    Odrv4 I__2092 (
            .O(N__20434),
            .I(\ALU.madd_490_14 ));
    CascadeMux I__2091 (
            .O(N__20431),
            .I(\ALU.r2_RNIFR6TZ0Z_15_cascade_ ));
    CascadeMux I__2090 (
            .O(N__20428),
            .I(\ALU.b_15_cascade_ ));
    InMux I__2089 (
            .O(N__20425),
            .I(N__20422));
    LocalMux I__2088 (
            .O(N__20422),
            .I(N__20418));
    InMux I__2087 (
            .O(N__20421),
            .I(N__20415));
    Odrv4 I__2086 (
            .O(N__20418),
            .I(\ALU.a5_b_9 ));
    LocalMux I__2085 (
            .O(N__20415),
            .I(\ALU.a5_b_9 ));
    CascadeMux I__2084 (
            .O(N__20410),
            .I(\ALU.a6_b_8_cascade_ ));
    InMux I__2083 (
            .O(N__20407),
            .I(N__20401));
    InMux I__2082 (
            .O(N__20406),
            .I(N__20401));
    LocalMux I__2081 (
            .O(N__20401),
            .I(N__20398));
    Odrv4 I__2080 (
            .O(N__20398),
            .I(\ALU.madd_378 ));
    CascadeMux I__2079 (
            .O(N__20395),
            .I(\ALU.b_i_3_cascade_ ));
    InMux I__2078 (
            .O(N__20392),
            .I(N__20389));
    LocalMux I__2077 (
            .O(N__20389),
            .I(N__20386));
    Odrv12 I__2076 (
            .O(N__20386),
            .I(\ALU.a3_b_11 ));
    InMux I__2075 (
            .O(N__20383),
            .I(N__20380));
    LocalMux I__2074 (
            .O(N__20380),
            .I(\ALU.madd_382 ));
    InMux I__2073 (
            .O(N__20377),
            .I(N__20374));
    LocalMux I__2072 (
            .O(N__20374),
            .I(N__20370));
    InMux I__2071 (
            .O(N__20373),
            .I(N__20367));
    Odrv4 I__2070 (
            .O(N__20370),
            .I(\ALU.a4_b_10 ));
    LocalMux I__2069 (
            .O(N__20367),
            .I(\ALU.a4_b_10 ));
    CascadeMux I__2068 (
            .O(N__20362),
            .I(\ALU.a11_b_3_cascade_ ));
    InMux I__2067 (
            .O(N__20359),
            .I(N__20356));
    LocalMux I__2066 (
            .O(N__20356),
            .I(\ALU.madd_373 ));
    CascadeMux I__2065 (
            .O(N__20353),
            .I(N__20350));
    InMux I__2064 (
            .O(N__20350),
            .I(N__20347));
    LocalMux I__2063 (
            .O(N__20347),
            .I(\ALU.a11_b_3 ));
    InMux I__2062 (
            .O(N__20344),
            .I(N__20341));
    LocalMux I__2061 (
            .O(N__20341),
            .I(N__20338));
    Span4Mux_h I__2060 (
            .O(N__20338),
            .I(N__20335));
    Span4Mux_s0_h I__2059 (
            .O(N__20335),
            .I(N__20332));
    Odrv4 I__2058 (
            .O(N__20332),
            .I(\ALU.madd_392 ));
    InMux I__2057 (
            .O(N__20329),
            .I(N__20326));
    LocalMux I__2056 (
            .O(N__20326),
            .I(\ALU.madd_490_16 ));
    CascadeMux I__2055 (
            .O(N__20323),
            .I(\ALU.madd_490_15_cascade_ ));
    InMux I__2054 (
            .O(N__20320),
            .I(N__20317));
    LocalMux I__2053 (
            .O(N__20317),
            .I(\ALU.madd_490_19 ));
    InMux I__2052 (
            .O(N__20314),
            .I(N__20311));
    LocalMux I__2051 (
            .O(N__20311),
            .I(N__20308));
    Span4Mux_v I__2050 (
            .O(N__20308),
            .I(N__20305));
    Odrv4 I__2049 (
            .O(N__20305),
            .I(\ALU.madd_339 ));
    CascadeMux I__2048 (
            .O(N__20302),
            .I(N__20299));
    InMux I__2047 (
            .O(N__20299),
            .I(N__20296));
    LocalMux I__2046 (
            .O(N__20296),
            .I(\ALU.madd_340_0 ));
    CascadeMux I__2045 (
            .O(N__20293),
            .I(\ALU.a7_b_7_cascade_ ));
    InMux I__2044 (
            .O(N__20290),
            .I(N__20287));
    LocalMux I__2043 (
            .O(N__20287),
            .I(N__20282));
    InMux I__2042 (
            .O(N__20286),
            .I(N__20277));
    InMux I__2041 (
            .O(N__20285),
            .I(N__20277));
    Odrv4 I__2040 (
            .O(N__20282),
            .I(\ALU.madd_383 ));
    LocalMux I__2039 (
            .O(N__20277),
            .I(\ALU.madd_383 ));
    CascadeMux I__2038 (
            .O(N__20272),
            .I(\ALU.b_9_cascade_ ));
    CascadeMux I__2037 (
            .O(N__20269),
            .I(N__20266));
    InMux I__2036 (
            .O(N__20266),
            .I(N__20263));
    LocalMux I__2035 (
            .O(N__20263),
            .I(\ALU.madd_326_0 ));
    CascadeMux I__2034 (
            .O(N__20260),
            .I(\ALU.a5_b_9_cascade_ ));
    InMux I__2033 (
            .O(N__20257),
            .I(N__20254));
    LocalMux I__2032 (
            .O(N__20254),
            .I(N__20251));
    Odrv4 I__2031 (
            .O(N__20251),
            .I(\ALU.a6_b_8 ));
    InMux I__2030 (
            .O(N__20248),
            .I(N__20242));
    InMux I__2029 (
            .O(N__20247),
            .I(N__20242));
    LocalMux I__2028 (
            .O(N__20242),
            .I(\ALU.madd_413_0 ));
    CascadeMux I__2027 (
            .O(N__20239),
            .I(\ALU.madd_418_cascade_ ));
    CascadeMux I__2026 (
            .O(N__20236),
            .I(N__20233));
    InMux I__2025 (
            .O(N__20233),
            .I(N__20227));
    InMux I__2024 (
            .O(N__20232),
            .I(N__20227));
    LocalMux I__2023 (
            .O(N__20227),
            .I(N__20224));
    Odrv12 I__2022 (
            .O(N__20224),
            .I(\ALU.madd_293 ));
    InMux I__2021 (
            .O(N__20221),
            .I(N__20215));
    InMux I__2020 (
            .O(N__20220),
            .I(N__20215));
    LocalMux I__2019 (
            .O(N__20215),
            .I(\ALU.madd_336_0 ));
    InMux I__2018 (
            .O(N__20212),
            .I(N__20208));
    InMux I__2017 (
            .O(N__20211),
            .I(N__20205));
    LocalMux I__2016 (
            .O(N__20208),
            .I(\ALU.madd_351 ));
    LocalMux I__2015 (
            .O(N__20205),
            .I(\ALU.madd_351 ));
    InMux I__2014 (
            .O(N__20200),
            .I(N__20197));
    LocalMux I__2013 (
            .O(N__20197),
            .I(\ALU.madd_346 ));
    InMux I__2012 (
            .O(N__20194),
            .I(N__20190));
    InMux I__2011 (
            .O(N__20193),
            .I(N__20187));
    LocalMux I__2010 (
            .O(N__20190),
            .I(\ALU.madd_172 ));
    LocalMux I__2009 (
            .O(N__20187),
            .I(\ALU.madd_172 ));
    CascadeMux I__2008 (
            .O(N__20182),
            .I(\ALU.madd_346_cascade_ ));
    InMux I__2007 (
            .O(N__20179),
            .I(N__20175));
    InMux I__2006 (
            .O(N__20178),
            .I(N__20172));
    LocalMux I__2005 (
            .O(N__20175),
            .I(\ALU.madd_298_0 ));
    LocalMux I__2004 (
            .O(N__20172),
            .I(\ALU.madd_298_0 ));
    InMux I__2003 (
            .O(N__20167),
            .I(N__20161));
    InMux I__2002 (
            .O(N__20166),
            .I(N__20161));
    LocalMux I__2001 (
            .O(N__20161),
            .I(\ALU.madd_360 ));
    InMux I__2000 (
            .O(N__20158),
            .I(N__20155));
    LocalMux I__1999 (
            .O(N__20155),
            .I(\ALU.madd_190 ));
    CascadeMux I__1998 (
            .O(N__20152),
            .I(N__20149));
    InMux I__1997 (
            .O(N__20149),
            .I(N__20146));
    LocalMux I__1996 (
            .O(N__20146),
            .I(\ALU.madd_330_0_tz ));
    InMux I__1995 (
            .O(N__20143),
            .I(N__20140));
    LocalMux I__1994 (
            .O(N__20140),
            .I(\ALU.madd_326 ));
    CascadeMux I__1993 (
            .O(N__20137),
            .I(\ALU.madd_326_cascade_ ));
    InMux I__1992 (
            .O(N__20134),
            .I(N__20131));
    LocalMux I__1991 (
            .O(N__20131),
            .I(\ALU.madd_350_0 ));
    InMux I__1990 (
            .O(N__20128),
            .I(N__20125));
    LocalMux I__1989 (
            .O(N__20125),
            .I(\ALU.madd_355 ));
    InMux I__1988 (
            .O(N__20122),
            .I(N__20118));
    InMux I__1987 (
            .O(N__20121),
            .I(N__20115));
    LocalMux I__1986 (
            .O(N__20118),
            .I(\ALU.madd_408 ));
    LocalMux I__1985 (
            .O(N__20115),
            .I(\ALU.madd_408 ));
    CascadeMux I__1984 (
            .O(N__20110),
            .I(\ALU.madd_350_0_cascade_ ));
    InMux I__1983 (
            .O(N__20107),
            .I(N__20104));
    LocalMux I__1982 (
            .O(N__20104),
            .I(N__20101));
    Odrv4 I__1981 (
            .O(N__20101),
            .I(\ALU.madd_422 ));
    InMux I__1980 (
            .O(N__20098),
            .I(N__20095));
    LocalMux I__1979 (
            .O(N__20095),
            .I(\ALU.madd_356 ));
    CascadeMux I__1978 (
            .O(N__20092),
            .I(N__20089));
    InMux I__1977 (
            .O(N__20089),
            .I(N__20083));
    InMux I__1976 (
            .O(N__20088),
            .I(N__20083));
    LocalMux I__1975 (
            .O(N__20083),
            .I(\ALU.madd_303_0 ));
    CascadeMux I__1974 (
            .O(N__20080),
            .I(\ALU.madd_356_cascade_ ));
    InMux I__1973 (
            .O(N__20077),
            .I(N__20071));
    InMux I__1972 (
            .O(N__20076),
            .I(N__20071));
    LocalMux I__1971 (
            .O(N__20071),
            .I(\ALU.madd_175 ));
    InMux I__1970 (
            .O(N__20068),
            .I(N__20065));
    LocalMux I__1969 (
            .O(N__20065),
            .I(N__20062));
    Span4Mux_s2_h I__1968 (
            .O(N__20062),
            .I(N__20059));
    Odrv4 I__1967 (
            .O(N__20059),
            .I(\ALU.madd_388_0 ));
    InMux I__1966 (
            .O(N__20056),
            .I(N__20053));
    LocalMux I__1965 (
            .O(N__20053),
            .I(N__20050));
    Odrv4 I__1964 (
            .O(N__20050),
            .I(\ALU.madd_393 ));
    InMux I__1963 (
            .O(N__20047),
            .I(N__20044));
    LocalMux I__1962 (
            .O(N__20044),
            .I(N__20040));
    InMux I__1961 (
            .O(N__20043),
            .I(N__20037));
    Span4Mux_v I__1960 (
            .O(N__20040),
            .I(N__20032));
    LocalMux I__1959 (
            .O(N__20037),
            .I(N__20032));
    Odrv4 I__1958 (
            .O(N__20032),
            .I(\ALU.madd_340 ));
    CascadeMux I__1957 (
            .O(N__20029),
            .I(\ALU.madd_355_cascade_ ));
    InMux I__1956 (
            .O(N__20026),
            .I(N__20023));
    LocalMux I__1955 (
            .O(N__20023),
            .I(\ALU.madd_418 ));
    CascadeMux I__1954 (
            .O(N__20020),
            .I(N__20017));
    InMux I__1953 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__1952 (
            .O(N__20014),
            .I(N__20010));
    InMux I__1951 (
            .O(N__20013),
            .I(N__20007));
    Odrv12 I__1950 (
            .O(N__20010),
            .I(\ALU.madd_181_0 ));
    LocalMux I__1949 (
            .O(N__20007),
            .I(\ALU.madd_181_0 ));
    CascadeMux I__1948 (
            .O(N__20002),
            .I(N__19999));
    InMux I__1947 (
            .O(N__19999),
            .I(N__19995));
    InMux I__1946 (
            .O(N__19998),
            .I(N__19992));
    LocalMux I__1945 (
            .O(N__19995),
            .I(N__19989));
    LocalMux I__1944 (
            .O(N__19992),
            .I(N__19986));
    Span4Mux_h I__1943 (
            .O(N__19989),
            .I(N__19983));
    Odrv12 I__1942 (
            .O(N__19986),
            .I(\ALU.madd_315_0 ));
    Odrv4 I__1941 (
            .O(N__19983),
            .I(\ALU.madd_315_0 ));
    InMux I__1940 (
            .O(N__19978),
            .I(N__19974));
    InMux I__1939 (
            .O(N__19977),
            .I(N__19971));
    LocalMux I__1938 (
            .O(N__19974),
            .I(N__19968));
    LocalMux I__1937 (
            .O(N__19971),
            .I(N__19965));
    Odrv4 I__1936 (
            .O(N__19968),
            .I(\ALU.madd_320 ));
    Odrv4 I__1935 (
            .O(N__19965),
            .I(\ALU.madd_320 ));
    CascadeMux I__1934 (
            .O(N__19960),
            .I(\ALU.madd_393_cascade_ ));
    InMux I__1933 (
            .O(N__19957),
            .I(N__19954));
    LocalMux I__1932 (
            .O(N__19954),
            .I(N__19951));
    Span4Mux_v I__1931 (
            .O(N__19951),
            .I(N__19948));
    Odrv4 I__1930 (
            .O(N__19948),
            .I(\ALU.madd_412 ));
    InMux I__1929 (
            .O(N__19945),
            .I(N__19939));
    InMux I__1928 (
            .O(N__19944),
            .I(N__19939));
    LocalMux I__1927 (
            .O(N__19939),
            .I(N__19936));
    Odrv4 I__1926 (
            .O(N__19936),
            .I(\ALU.madd_308_0_tz_0 ));
    CascadeMux I__1925 (
            .O(N__19933),
            .I(N__19930));
    InMux I__1924 (
            .O(N__19930),
            .I(N__19924));
    InMux I__1923 (
            .O(N__19929),
            .I(N__19924));
    LocalMux I__1922 (
            .O(N__19924),
            .I(\ALU.madd_299 ));
    InMux I__1921 (
            .O(N__19921),
            .I(N__19917));
    InMux I__1920 (
            .O(N__19920),
            .I(N__19914));
    LocalMux I__1919 (
            .O(N__19917),
            .I(\ALU.madd_209 ));
    LocalMux I__1918 (
            .O(N__19914),
            .I(\ALU.madd_209 ));
    InMux I__1917 (
            .O(N__19909),
            .I(N__19903));
    InMux I__1916 (
            .O(N__19908),
            .I(N__19903));
    LocalMux I__1915 (
            .O(N__19903),
            .I(\ALU.madd_243 ));
    CascadeMux I__1914 (
            .O(N__19900),
            .I(\ALU.a0_b_13_cascade_ ));
    InMux I__1913 (
            .O(N__19897),
            .I(N__19894));
    LocalMux I__1912 (
            .O(N__19894),
            .I(N__19891));
    Sp12to4 I__1911 (
            .O(N__19891),
            .I(N__19888));
    Odrv12 I__1910 (
            .O(N__19888),
            .I(\ALU.g2_0_1 ));
    InMux I__1909 (
            .O(N__19885),
            .I(N__19880));
    CascadeMux I__1908 (
            .O(N__19884),
            .I(N__19877));
    CascadeMux I__1907 (
            .O(N__19883),
            .I(N__19874));
    LocalMux I__1906 (
            .O(N__19880),
            .I(N__19871));
    InMux I__1905 (
            .O(N__19877),
            .I(N__19866));
    InMux I__1904 (
            .O(N__19874),
            .I(N__19866));
    Span4Mux_s1_v I__1903 (
            .O(N__19871),
            .I(N__19863));
    LocalMux I__1902 (
            .O(N__19866),
            .I(N__19860));
    Odrv4 I__1901 (
            .O(N__19863),
            .I(\ALU.madd_182_0 ));
    Odrv4 I__1900 (
            .O(N__19860),
            .I(\ALU.madd_182_0 ));
    CascadeMux I__1899 (
            .O(N__19855),
            .I(N__19851));
    InMux I__1898 (
            .O(N__19854),
            .I(N__19847));
    InMux I__1897 (
            .O(N__19851),
            .I(N__19842));
    InMux I__1896 (
            .O(N__19850),
            .I(N__19842));
    LocalMux I__1895 (
            .O(N__19847),
            .I(\ALU.a3_b_7 ));
    LocalMux I__1894 (
            .O(N__19842),
            .I(\ALU.a3_b_7 ));
    CascadeMux I__1893 (
            .O(N__19837),
            .I(N__19834));
    InMux I__1892 (
            .O(N__19834),
            .I(N__19830));
    InMux I__1891 (
            .O(N__19833),
            .I(N__19827));
    LocalMux I__1890 (
            .O(N__19830),
            .I(N__19824));
    LocalMux I__1889 (
            .O(N__19827),
            .I(\ALU.a2_b_8 ));
    Odrv4 I__1888 (
            .O(N__19824),
            .I(\ALU.a2_b_8 ));
    InMux I__1887 (
            .O(N__19819),
            .I(N__19816));
    LocalMux I__1886 (
            .O(N__19816),
            .I(N__19810));
    InMux I__1885 (
            .O(N__19815),
            .I(N__19803));
    InMux I__1884 (
            .O(N__19814),
            .I(N__19803));
    InMux I__1883 (
            .O(N__19813),
            .I(N__19803));
    Odrv4 I__1882 (
            .O(N__19810),
            .I(\ALU.madd_177 ));
    LocalMux I__1881 (
            .O(N__19803),
            .I(\ALU.madd_177 ));
    InMux I__1880 (
            .O(N__19798),
            .I(N__19792));
    InMux I__1879 (
            .O(N__19797),
            .I(N__19792));
    LocalMux I__1878 (
            .O(N__19792),
            .I(\ALU.madd_229 ));
    CascadeMux I__1877 (
            .O(N__19789),
            .I(\ALU.madd_243_cascade_ ));
    InMux I__1876 (
            .O(N__19786),
            .I(N__19778));
    InMux I__1875 (
            .O(N__19785),
            .I(N__19778));
    InMux I__1874 (
            .O(N__19784),
            .I(N__19773));
    InMux I__1873 (
            .O(N__19783),
            .I(N__19773));
    LocalMux I__1872 (
            .O(N__19778),
            .I(\ALU.madd_219_0 ));
    LocalMux I__1871 (
            .O(N__19773),
            .I(\ALU.madd_219_0 ));
    CascadeMux I__1870 (
            .O(N__19768),
            .I(N__19764));
    InMux I__1869 (
            .O(N__19767),
            .I(N__19759));
    InMux I__1868 (
            .O(N__19764),
            .I(N__19759));
    LocalMux I__1867 (
            .O(N__19759),
            .I(\ALU.madd_192_0 ));
    InMux I__1866 (
            .O(N__19756),
            .I(N__19747));
    InMux I__1865 (
            .O(N__19755),
            .I(N__19747));
    InMux I__1864 (
            .O(N__19754),
            .I(N__19747));
    LocalMux I__1863 (
            .O(N__19747),
            .I(\ALU.madd_144 ));
    InMux I__1862 (
            .O(N__19744),
            .I(N__19741));
    LocalMux I__1861 (
            .O(N__19741),
            .I(\ALU.g0_1 ));
    CascadeMux I__1860 (
            .O(N__19738),
            .I(N__19735));
    InMux I__1859 (
            .O(N__19735),
            .I(N__19732));
    LocalMux I__1858 (
            .O(N__19732),
            .I(N__19729));
    Odrv4 I__1857 (
            .O(N__19729),
            .I(\ALU.N_695_0 ));
    InMux I__1856 (
            .O(N__19726),
            .I(N__19723));
    LocalMux I__1855 (
            .O(N__19723),
            .I(\ALU.g0_4 ));
    InMux I__1854 (
            .O(N__19720),
            .I(N__19714));
    InMux I__1853 (
            .O(N__19719),
            .I(N__19714));
    LocalMux I__1852 (
            .O(N__19714),
            .I(\ALU.madd_197 ));
    InMux I__1851 (
            .O(N__19711),
            .I(N__19707));
    InMux I__1850 (
            .O(N__19710),
            .I(N__19704));
    LocalMux I__1849 (
            .O(N__19707),
            .I(\ALU.madd_112 ));
    LocalMux I__1848 (
            .O(N__19704),
            .I(\ALU.madd_112 ));
    InMux I__1847 (
            .O(N__19699),
            .I(N__19692));
    InMux I__1846 (
            .O(N__19698),
            .I(N__19692));
    InMux I__1845 (
            .O(N__19697),
            .I(N__19689));
    LocalMux I__1844 (
            .O(N__19692),
            .I(N__19686));
    LocalMux I__1843 (
            .O(N__19689),
            .I(\ALU.madd_191 ));
    Odrv4 I__1842 (
            .O(N__19686),
            .I(\ALU.madd_191 ));
    InMux I__1841 (
            .O(N__19681),
            .I(N__19678));
    LocalMux I__1840 (
            .O(N__19678),
            .I(N__19675));
    Odrv4 I__1839 (
            .O(N__19675),
            .I(\ALU.madd_234 ));
    CascadeMux I__1838 (
            .O(N__19672),
            .I(\ALU.madd_112_cascade_ ));
    InMux I__1837 (
            .O(N__19669),
            .I(N__19665));
    InMux I__1836 (
            .O(N__19668),
            .I(N__19660));
    LocalMux I__1835 (
            .O(N__19665),
            .I(N__19657));
    InMux I__1834 (
            .O(N__19664),
            .I(N__19654));
    InMux I__1833 (
            .O(N__19663),
            .I(N__19651));
    LocalMux I__1832 (
            .O(N__19660),
            .I(\ALU.madd_196_0 ));
    Odrv4 I__1831 (
            .O(N__19657),
            .I(\ALU.madd_196_0 ));
    LocalMux I__1830 (
            .O(N__19654),
            .I(\ALU.madd_196_0 ));
    LocalMux I__1829 (
            .O(N__19651),
            .I(\ALU.madd_196_0 ));
    InMux I__1828 (
            .O(N__19642),
            .I(N__19636));
    InMux I__1827 (
            .O(N__19641),
            .I(N__19631));
    InMux I__1826 (
            .O(N__19640),
            .I(N__19631));
    InMux I__1825 (
            .O(N__19639),
            .I(N__19628));
    LocalMux I__1824 (
            .O(N__19636),
            .I(\ALU.madd_187 ));
    LocalMux I__1823 (
            .O(N__19631),
            .I(\ALU.madd_187 ));
    LocalMux I__1822 (
            .O(N__19628),
            .I(\ALU.madd_187 ));
    InMux I__1821 (
            .O(N__19621),
            .I(N__19615));
    InMux I__1820 (
            .O(N__19620),
            .I(N__19615));
    LocalMux I__1819 (
            .O(N__19615),
            .I(\ALU.madd_154 ));
    InMux I__1818 (
            .O(N__19612),
            .I(N__19606));
    InMux I__1817 (
            .O(N__19611),
            .I(N__19606));
    LocalMux I__1816 (
            .O(N__19606),
            .I(\ALU.madd_134 ));
    InMux I__1815 (
            .O(N__19603),
            .I(clkdiv_cry_22));
    IoInMux I__1814 (
            .O(N__19600),
            .I(N__19597));
    LocalMux I__1813 (
            .O(N__19597),
            .I(N__19594));
    Span12Mux_s8_v I__1812 (
            .O(N__19594),
            .I(N__19590));
    InMux I__1811 (
            .O(N__19593),
            .I(N__19587));
    Odrv12 I__1810 (
            .O(N__19590),
            .I(GPIO3_c));
    LocalMux I__1809 (
            .O(N__19587),
            .I(GPIO3_c));
    CascadeMux I__1808 (
            .O(N__19582),
            .I(\ALU.madd_154_cascade_ ));
    CascadeMux I__1807 (
            .O(N__19579),
            .I(\ALU.N_703_1_cascade_ ));
    CascadeMux I__1806 (
            .O(N__19576),
            .I(\ALU.g0_cascade_ ));
    InMux I__1805 (
            .O(N__19573),
            .I(N__19567));
    InMux I__1804 (
            .O(N__19572),
            .I(N__19567));
    LocalMux I__1803 (
            .O(N__19567),
            .I(\ALU.madd_206 ));
    CascadeMux I__1802 (
            .O(N__19564),
            .I(\ALU.madd_334_cascade_ ));
    InMux I__1801 (
            .O(N__19561),
            .I(N__19558));
    LocalMux I__1800 (
            .O(N__19558),
            .I(\ALU.N_724_0_0_0 ));
    InMux I__1799 (
            .O(N__19555),
            .I(N__19552));
    LocalMux I__1798 (
            .O(N__19552),
            .I(clkdivZ0Z_14));
    InMux I__1797 (
            .O(N__19549),
            .I(clkdiv_cry_13));
    InMux I__1796 (
            .O(N__19546),
            .I(N__19543));
    LocalMux I__1795 (
            .O(N__19543),
            .I(clkdivZ0Z_15));
    InMux I__1794 (
            .O(N__19540),
            .I(clkdiv_cry_14));
    InMux I__1793 (
            .O(N__19537),
            .I(N__19534));
    LocalMux I__1792 (
            .O(N__19534),
            .I(clkdivZ0Z_16));
    InMux I__1791 (
            .O(N__19531),
            .I(bfn_1_17_0_));
    InMux I__1790 (
            .O(N__19528),
            .I(N__19525));
    LocalMux I__1789 (
            .O(N__19525),
            .I(clkdivZ0Z_17));
    InMux I__1788 (
            .O(N__19522),
            .I(clkdiv_cry_16));
    InMux I__1787 (
            .O(N__19519),
            .I(N__19516));
    LocalMux I__1786 (
            .O(N__19516),
            .I(clkdivZ0Z_18));
    InMux I__1785 (
            .O(N__19513),
            .I(clkdiv_cry_17));
    InMux I__1784 (
            .O(N__19510),
            .I(N__19507));
    LocalMux I__1783 (
            .O(N__19507),
            .I(clkdivZ0Z_19));
    InMux I__1782 (
            .O(N__19504),
            .I(clkdiv_cry_18));
    InMux I__1781 (
            .O(N__19501),
            .I(N__19498));
    LocalMux I__1780 (
            .O(N__19498),
            .I(clkdivZ0Z_20));
    InMux I__1779 (
            .O(N__19495),
            .I(clkdiv_cry_19));
    InMux I__1778 (
            .O(N__19492),
            .I(N__19489));
    LocalMux I__1777 (
            .O(N__19489),
            .I(clkdivZ0Z_21));
    InMux I__1776 (
            .O(N__19486),
            .I(clkdiv_cry_20));
    InMux I__1775 (
            .O(N__19483),
            .I(N__19480));
    LocalMux I__1774 (
            .O(N__19480),
            .I(clkdivZ0Z_22));
    InMux I__1773 (
            .O(N__19477),
            .I(clkdiv_cry_21));
    InMux I__1772 (
            .O(N__19474),
            .I(clkdiv_cry_5));
    InMux I__1771 (
            .O(N__19471),
            .I(clkdiv_cry_6));
    InMux I__1770 (
            .O(N__19468),
            .I(N__19465));
    LocalMux I__1769 (
            .O(N__19465),
            .I(clkdivZ0Z_8));
    InMux I__1768 (
            .O(N__19462),
            .I(bfn_1_16_0_));
    InMux I__1767 (
            .O(N__19459),
            .I(N__19456));
    LocalMux I__1766 (
            .O(N__19456),
            .I(clkdivZ0Z_9));
    InMux I__1765 (
            .O(N__19453),
            .I(clkdiv_cry_8));
    InMux I__1764 (
            .O(N__19450),
            .I(N__19447));
    LocalMux I__1763 (
            .O(N__19447),
            .I(clkdivZ0Z_10));
    InMux I__1762 (
            .O(N__19444),
            .I(clkdiv_cry_9));
    InMux I__1761 (
            .O(N__19441),
            .I(N__19438));
    LocalMux I__1760 (
            .O(N__19438),
            .I(clkdivZ0Z_11));
    InMux I__1759 (
            .O(N__19435),
            .I(clkdiv_cry_10));
    InMux I__1758 (
            .O(N__19432),
            .I(N__19429));
    LocalMux I__1757 (
            .O(N__19429),
            .I(clkdivZ0Z_12));
    InMux I__1756 (
            .O(N__19426),
            .I(clkdiv_cry_11));
    InMux I__1755 (
            .O(N__19423),
            .I(N__19420));
    LocalMux I__1754 (
            .O(N__19420),
            .I(clkdivZ0Z_13));
    InMux I__1753 (
            .O(N__19417),
            .I(clkdiv_cry_12));
    InMux I__1752 (
            .O(N__19414),
            .I(N__19411));
    LocalMux I__1751 (
            .O(N__19411),
            .I(TXbuffer_RNO_1Z0Z_3));
    InMux I__1750 (
            .O(N__19408),
            .I(bfn_1_15_0_));
    InMux I__1749 (
            .O(N__19405),
            .I(clkdiv_cry_0));
    InMux I__1748 (
            .O(N__19402),
            .I(clkdiv_cry_1));
    InMux I__1747 (
            .O(N__19399),
            .I(clkdiv_cry_2));
    InMux I__1746 (
            .O(N__19396),
            .I(clkdiv_cry_3));
    InMux I__1745 (
            .O(N__19393),
            .I(clkdiv_cry_4));
    CascadeMux I__1744 (
            .O(N__19390),
            .I(TXbuffer_RNO_5Z0Z_4_cascade_));
    CascadeMux I__1743 (
            .O(N__19387),
            .I(TXbuffer_18_15_ns_1_4_cascade_));
    InMux I__1742 (
            .O(N__19384),
            .I(N__19381));
    LocalMux I__1741 (
            .O(N__19381),
            .I(TXbuffer_RNO_1Z0Z_0));
    CascadeMux I__1740 (
            .O(N__19378),
            .I(TXbuffer_18_15_ns_1_0_cascade_));
    CascadeMux I__1739 (
            .O(N__19375),
            .I(TXbuffer_18_10_ns_1_3_cascade_));
    CascadeMux I__1738 (
            .O(N__19372),
            .I(TXbuffer_RNO_0Z0Z_3_cascade_));
    CascadeMux I__1737 (
            .O(N__19369),
            .I(TXbuffer_18_10_ns_1_4_cascade_));
    InMux I__1736 (
            .O(N__19366),
            .I(N__19363));
    LocalMux I__1735 (
            .O(N__19363),
            .I(N__19360));
    Odrv4 I__1734 (
            .O(N__19360),
            .I(TXbuffer_RNO_0Z0Z_4));
    CascadeMux I__1733 (
            .O(N__19357),
            .I(\ALU.a6_b_9_cascade_ ));
    CascadeMux I__1732 (
            .O(N__19354),
            .I(\ALU.madd_490_10_cascade_ ));
    CascadeMux I__1731 (
            .O(N__19351),
            .I(\ALU.madd_490_7_cascade_ ));
    InMux I__1730 (
            .O(N__19348),
            .I(N__19345));
    LocalMux I__1729 (
            .O(N__19345),
            .I(\ALU.madd_490_11 ));
    InMux I__1728 (
            .O(N__19342),
            .I(N__19339));
    LocalMux I__1727 (
            .O(N__19339),
            .I(\ALU.a2_b_13 ));
    CascadeMux I__1726 (
            .O(N__19336),
            .I(TXbuffer_18_13_ns_1_0_cascade_));
    CascadeMux I__1725 (
            .O(N__19333),
            .I(TXbuffer_18_6_ns_1_2_cascade_));
    CascadeMux I__1724 (
            .O(N__19330),
            .I(TXbuffer_RNO_6Z0Z_2_cascade_));
    InMux I__1723 (
            .O(N__19327),
            .I(N__19324));
    LocalMux I__1722 (
            .O(N__19324),
            .I(N__19321));
    Odrv4 I__1721 (
            .O(N__19321),
            .I(\ALU.madd_417 ));
    CascadeMux I__1720 (
            .O(N__19318),
            .I(\ALU.madd_490_1_0_cascade_ ));
    CascadeMux I__1719 (
            .O(N__19315),
            .I(N__19312));
    InMux I__1718 (
            .O(N__19312),
            .I(N__19309));
    LocalMux I__1717 (
            .O(N__19309),
            .I(N__19306));
    Span4Mux_v I__1716 (
            .O(N__19306),
            .I(N__19303));
    Odrv4 I__1715 (
            .O(N__19303),
            .I(\ALU.madd_378_0 ));
    InMux I__1714 (
            .O(N__19300),
            .I(N__19297));
    LocalMux I__1713 (
            .O(N__19297),
            .I(N__19294));
    Odrv4 I__1712 (
            .O(N__19294),
            .I(\ALU.madd_388 ));
    CascadeMux I__1711 (
            .O(N__19291),
            .I(\ALU.madd_402_cascade_ ));
    InMux I__1710 (
            .O(N__19288),
            .I(N__19285));
    LocalMux I__1709 (
            .O(N__19285),
            .I(N__19280));
    InMux I__1708 (
            .O(N__19284),
            .I(N__19275));
    InMux I__1707 (
            .O(N__19283),
            .I(N__19275));
    Odrv12 I__1706 (
            .O(N__19280),
            .I(\ALU.madd_330 ));
    LocalMux I__1705 (
            .O(N__19275),
            .I(\ALU.madd_330 ));
    InMux I__1704 (
            .O(N__19270),
            .I(N__19267));
    LocalMux I__1703 (
            .O(N__19267),
            .I(\ALU.madd_490_21 ));
    InMux I__1702 (
            .O(N__19264),
            .I(N__19261));
    LocalMux I__1701 (
            .O(N__19261),
            .I(N__19258));
    Odrv4 I__1700 (
            .O(N__19258),
            .I(\ALU.madd_397 ));
    CascadeMux I__1699 (
            .O(N__19255),
            .I(\ALU.madd_388_cascade_ ));
    CascadeMux I__1698 (
            .O(N__19252),
            .I(\ALU.madd_403_cascade_ ));
    CascadeMux I__1697 (
            .O(N__19249),
            .I(N__19246));
    InMux I__1696 (
            .O(N__19246),
            .I(N__19243));
    LocalMux I__1695 (
            .O(N__19243),
            .I(\ALU.a1_b_13 ));
    CascadeMux I__1694 (
            .O(N__19240),
            .I(\ALU.madd_403_0_cascade_ ));
    CascadeMux I__1693 (
            .O(N__19237),
            .I(\ALU.a_6_ns_1_2_cascade_ ));
    CascadeMux I__1692 (
            .O(N__19234),
            .I(TXbuffer_18_13_ns_1_2_cascade_));
    CascadeMux I__1691 (
            .O(N__19231),
            .I(\ALU.madd_311_cascade_ ));
    InMux I__1690 (
            .O(N__19228),
            .I(N__19225));
    LocalMux I__1689 (
            .O(N__19225),
            .I(\ALU.madd_268 ));
    CascadeMux I__1688 (
            .O(N__19222),
            .I(\ALU.madd_268_cascade_ ));
    InMux I__1687 (
            .O(N__19219),
            .I(N__19216));
    LocalMux I__1686 (
            .O(N__19216),
            .I(\ALU.madd_311 ));
    InMux I__1685 (
            .O(N__19213),
            .I(N__19207));
    InMux I__1684 (
            .O(N__19212),
            .I(N__19207));
    LocalMux I__1683 (
            .O(N__19207),
            .I(\ALU.madd_316 ));
    InMux I__1682 (
            .O(N__19204),
            .I(N__19198));
    InMux I__1681 (
            .O(N__19203),
            .I(N__19198));
    LocalMux I__1680 (
            .O(N__19198),
            .I(\ALU.a8_b_5 ));
    CascadeMux I__1679 (
            .O(N__19195),
            .I(\ALU.a1_b_13_cascade_ ));
    InMux I__1678 (
            .O(N__19192),
            .I(N__19189));
    LocalMux I__1677 (
            .O(N__19189),
            .I(\ALU.madd_171_0_tz ));
    CascadeMux I__1676 (
            .O(N__19186),
            .I(\ALU.madd_171_cascade_ ));
    CascadeMux I__1675 (
            .O(N__19183),
            .I(\ALU.madd_315_0_tz_cascade_ ));
    InMux I__1674 (
            .O(N__19180),
            .I(N__19176));
    InMux I__1673 (
            .O(N__19179),
            .I(N__19173));
    LocalMux I__1672 (
            .O(N__19176),
            .I(\ALU.madd_214 ));
    LocalMux I__1671 (
            .O(N__19173),
            .I(\ALU.madd_214 ));
    CascadeMux I__1670 (
            .O(N__19168),
            .I(\ALU.madd_234_cascade_ ));
    CascadeMux I__1669 (
            .O(N__19165),
            .I(\ALU.a7_b_8_cascade_ ));
    InMux I__1668 (
            .O(N__19162),
            .I(N__19159));
    LocalMux I__1667 (
            .O(N__19159),
            .I(\ALU.madd_490_3 ));
    CascadeMux I__1666 (
            .O(N__19156),
            .I(\ALU.madd_171_0_tz_cascade_ ));
    InMux I__1665 (
            .O(N__19153),
            .I(N__19150));
    LocalMux I__1664 (
            .O(N__19150),
            .I(\ALU.madd_97 ));
    CascadeMux I__1663 (
            .O(N__19147),
            .I(\ALU.madd_171_x_cascade_ ));
    InMux I__1662 (
            .O(N__19144),
            .I(N__19141));
    LocalMux I__1661 (
            .O(N__19141),
            .I(\ALU.g0_2 ));
    CascadeMux I__1660 (
            .O(N__19138),
            .I(\ALU.a5_b_4_cascade_ ));
    InMux I__1659 (
            .O(N__19135),
            .I(N__19126));
    InMux I__1658 (
            .O(N__19134),
            .I(N__19126));
    InMux I__1657 (
            .O(N__19133),
            .I(N__19126));
    LocalMux I__1656 (
            .O(N__19126),
            .I(\ALU.madd_139 ));
    CascadeMux I__1655 (
            .O(N__19123),
            .I(\ALU.a2_b_8_cascade_ ));
    CascadeMux I__1654 (
            .O(N__19120),
            .I(\ALU.madd_181_cascade_ ));
    InMux I__1653 (
            .O(N__19117),
            .I(N__19110));
    InMux I__1652 (
            .O(N__19116),
            .I(N__19110));
    InMux I__1651 (
            .O(N__19115),
            .I(N__19107));
    LocalMux I__1650 (
            .O(N__19110),
            .I(\ALU.a3_b_8 ));
    LocalMux I__1649 (
            .O(N__19107),
            .I(\ALU.a3_b_8 ));
    CascadeMux I__1648 (
            .O(N__19102),
            .I(\ALU.a3_b_8_cascade_ ));
    CascadeMux I__1647 (
            .O(N__19099),
            .I(N__19095));
    InMux I__1646 (
            .O(N__19098),
            .I(N__19092));
    InMux I__1645 (
            .O(N__19095),
            .I(N__19089));
    LocalMux I__1644 (
            .O(N__19092),
            .I(\ALU.madd_181 ));
    LocalMux I__1643 (
            .O(N__19089),
            .I(\ALU.madd_181 ));
    CascadeMux I__1642 (
            .O(N__19084),
            .I(\ALU.N_675_0_0_cascade_ ));
    CascadeMux I__1641 (
            .O(N__19081),
            .I(\ALU.N_703_0_0_0_cascade_ ));
    InMux I__1640 (
            .O(N__19078),
            .I(N__19075));
    LocalMux I__1639 (
            .O(N__19075),
            .I(N__19072));
    Odrv4 I__1638 (
            .O(N__19072),
            .I(\ALU.N_681_0_0_0 ));
    CascadeMux I__1637 (
            .O(N__19069),
            .I(\ALU.g0_0_2_cascade_ ));
    InMux I__1636 (
            .O(N__19066),
            .I(N__19063));
    LocalMux I__1635 (
            .O(N__19063),
            .I(\ALU.N_699_0 ));
    CascadeMux I__1634 (
            .O(N__19060),
            .I(\ALU.madd_167_cascade_ ));
    InMux I__1633 (
            .O(N__19057),
            .I(N__19051));
    InMux I__1632 (
            .O(N__19056),
            .I(N__19051));
    LocalMux I__1631 (
            .O(N__19051),
            .I(\ALU.madd_167 ));
    INV \INVFTDI.baudAcc_0C  (
            .O(\INVFTDI.baudAcc_0C_net ),
            .I(N__56247));
    INV \INVFTDI.TXstate_3C  (
            .O(\INVFTDI.TXstate_3C_net ),
            .I(N__56244));
    INV \INVFTDI.TXstate_0C  (
            .O(\INVFTDI.TXstate_0C_net ),
            .I(N__56238));
    INV \INVFTDI.TXshift_0C  (
            .O(\INVFTDI.TXshift_0C_net ),
            .I(N__56243));
    INV \INVFTDI.TXstate_2C  (
            .O(\INVFTDI.TXstate_2C_net ),
            .I(N__56237));
    INV \INVFTDI.TXstate_1C  (
            .O(\INVFTDI.TXstate_1C_net ),
            .I(N__56235));
    INV \INVFTDI.TXshift_4C  (
            .O(\INVFTDI.TXshift_4C_net ),
            .I(N__56239));
    INV \INVFTDI.TXshift_1C  (
            .O(\INVFTDI.TXshift_1C_net ),
            .I(N__56236));
    INV \INVFTDI.TXshift_7C  (
            .O(\INVFTDI.TXshift_7C_net ),
            .I(N__56233));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(\ALU.r0_12_prm_2_7_s1 ),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\ALU.r0_12_prm_2_7_s0 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(\ALU.r0_12_prm_2_6_s1 ),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_13_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_3_0_));
    defparam IN_MUX_bfv_13_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_4_0_ (
            .carryinitin(\ALU.r0_12_prm_2_6_s0 ),
            .carryinitout(bfn_13_4_0_));
    defparam IN_MUX_bfv_13_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_5_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(\ALU.r0_12_prm_2_4 ),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_16_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_5_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(\ALU.r0_12_prm_2_3 ),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_14_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_1_0_));
    defparam IN_MUX_bfv_14_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_2_0_ (
            .carryinitin(\ALU.r0_12_prm_2_2 ),
            .carryinitout(bfn_14_2_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\ALU.r0_12_prm_2_1 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_18_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_6_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\ALU.r0_12_prm_2_9_s1 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\ALU.r0_12_prm_2_9_s0 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\ALU.r0_12_prm_2_8_s1 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\ALU.r0_12_prm_2_8_s0 ),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\ALU.r0_12_prm_2_5_s1 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\ALU.r0_12_prm_2_5_s0 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\ALU.r0_12_prm_2_15_s1 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\ALU.r0_12_prm_2_15_s0 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\ALU.r0_12_prm_2_14_s1 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\ALU.r0_12_prm_2_14_s0 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\ALU.r0_12_prm_2_13_s1 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_6_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_16_0_ (
            .carryinitin(\ALU.r0_12_prm_2_13_s0 ),
            .carryinitout(bfn_6_16_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\ALU.r0_12_prm_2_12_s1 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\ALU.r0_12_prm_2_12_s0 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(\ALU.r0_12_prm_2_11_s1 ),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\ALU.r0_12_prm_2_11_s0 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\ALU.r0_12_prm_2_10_s1 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\ALU.r0_12_prm_2_10_s0 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(\ALU.r0_12_s1_0 ),
            .carryinitout(bfn_12_3_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\ALU.r0_12_s0_0 ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\ALU.madd_cry_7 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(clkdiv_cry_7),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(clkdiv_cry_15),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\ALU.un9_addsub_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\ALU.un2_addsub_cry_7 ),
            .carryinitout(bfn_10_10_0_));
    ICE_GB clkdiv_RNIQAHO1_0_0 (
            .USERSIGNALTOGLOBALBUFFER(N__26956),
            .GLOBALBUFFEROUTPUT(params5_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \ALU.mult_madd_159_N_2L1_LC_1_1_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_159_N_2L1_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_159_N_2L1_LC_1_1_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ALU.mult_madd_159_N_2L1_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(N__46375),
            .in2(_gnd_net_),
            .in3(N__48612),
            .lcout(\ALU.madd_159_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_134_LC_1_1_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_134_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_134_LC_1_1_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_madd_134_LC_1_1_1  (
            .in0(N__22123),
            .in1(N__38018),
            .in2(N__23050),
            .in3(N__52275),
            .lcout(\ALU.madd_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_17_LC_1_1_2 .C_ON=1'b0;
    defparam \ALU.mult_g0_17_LC_1_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_17_LC_1_1_2 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_g0_17_LC_1_1_2  (
            .in0(N__47424),
            .in1(N__49003),
            .in2(N__20524),
            .in3(N__22096),
            .lcout(\ALU.N_681_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_20_LC_1_1_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_20_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_20_LC_1_1_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_g0_20_LC_1_1_3  (
            .in0(N__22122),
            .in1(N__38019),
            .in2(N__23049),
            .in3(N__52276),
            .lcout(),
            .ltout(\ALU.N_675_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_15_LC_1_1_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_15_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_15_LC_1_1_4 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_g0_15_LC_1_1_4  (
            .in0(N__19897),
            .in1(N__19639),
            .in2(N__19084),
            .in3(N__21535),
            .lcout(),
            .ltout(\ALU.N_703_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_1_LC_1_1_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_1_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_1_LC_1_1_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_1_LC_1_1_5  (
            .in0(N__20641),
            .in1(N__19066),
            .in2(N__19081),
            .in3(N__19144),
            .lcout(),
            .ltout(\ALU.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_14_LC_1_1_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_14_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_14_LC_1_1_6 .LUT_INIT=16'b0000111101111000;
    LogicCell40 \ALU.mult_g0_14_LC_1_1_6  (
            .in0(N__19819),
            .in1(N__19078),
            .in2(N__19069),
            .in3(N__19668),
            .lcout(\ALU.N_724_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_18_LC_1_2_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_18_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_18_LC_1_2_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_g0_18_LC_1_2_0  (
            .in0(N__19057),
            .in1(N__19135),
            .in2(_gnd_net_),
            .in3(N__19756),
            .lcout(\ALU.N_699_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_167_LC_1_2_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_167_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_167_LC_1_2_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ALU.mult_madd_167_LC_1_2_1  (
            .in0(N__22189),
            .in1(N__52253),
            .in2(_gnd_net_),
            .in3(N__46796),
            .lcout(\ALU.madd_167 ),
            .ltout(\ALU.madd_167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_187_LC_1_2_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_187_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_187_LC_1_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_187_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(N__19133),
            .in2(N__19060),
            .in3(N__19754),
            .lcout(\ALU.madd_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_1_0_LC_1_2_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_1_0_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_1_0_LC_1_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_g0_1_0_LC_1_2_3  (
            .in0(N__19116),
            .in1(N__19785),
            .in2(_gnd_net_),
            .in3(N__21741),
            .lcout(\ALU.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_191_LC_1_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_191_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_191_LC_1_2_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_191_LC_1_2_4  (
            .in0(N__19056),
            .in1(N__19134),
            .in2(_gnd_net_),
            .in3(N__19755),
            .lcout(\ALU.madd_191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_2_0_LC_1_2_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_2_0_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_2_0_LC_1_2_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_2_0_LC_1_2_5  (
            .in0(N__19117),
            .in1(N__19786),
            .in2(N__19099),
            .in3(N__21742),
            .lcout(\ALU.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_4_LC_1_2_6 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_4_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_4_LC_1_2_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a5_b_4_LC_1_2_6  (
            .in0(N__29101),
            .in1(N__29013),
            .in2(N__29245),
            .in3(N__40530),
            .lcout(),
            .ltout(\ALU.a5_b_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_139_LC_1_2_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_139_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_139_LC_1_2_7 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_139_LC_1_2_7  (
            .in0(N__43393),
            .in1(N__21874),
            .in2(N__19138),
            .in3(N__44349),
            .lcout(\ALU.madd_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_10_LC_1_3_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_10_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_10_LC_1_3_0 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_g0_10_LC_1_3_0  (
            .in0(N__42827),
            .in1(N__43637),
            .in2(N__19855),
            .in3(N__19833),
            .lcout(\ALU.N_695_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_7_LC_1_3_1 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_7_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_7_LC_1_3_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a3_b_7_LC_1_3_1  (
            .in0(N__44723),
            .in1(N__31922),
            .in2(N__36769),
            .in3(N__31834),
            .lcout(\ALU.a3_b_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_8_LC_1_3_2 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_8_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_8_LC_1_3_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a2_b_8_LC_1_3_2  (
            .in0(N__32665),
            .in1(N__32590),
            .in2(N__29244),
            .in3(N__46334),
            .lcout(\ALU.a2_b_8 ),
            .ltout(\ALU.a2_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_181_LC_1_3_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_181_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_181_LC_1_3_3 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_181_LC_1_3_3  (
            .in0(N__43636),
            .in1(N__19850),
            .in2(N__19123),
            .in3(N__42826),
            .lcout(\ALU.madd_181 ),
            .ltout(\ALU.madd_181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_238_LC_1_3_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_238_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_238_LC_1_3_4 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \ALU.mult_madd_238_LC_1_3_4  (
            .in0(N__21734),
            .in1(N__19783),
            .in2(N__19120),
            .in3(N__19115),
            .lcout(\ALU.madd_238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_8_LC_1_3_5 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_8_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_8_LC_1_3_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a3_b_8_LC_1_3_5  (
            .in0(N__46335),
            .in1(N__31923),
            .in2(N__32262),
            .in3(N__31835),
            .lcout(\ALU.a3_b_8 ),
            .ltout(\ALU.a3_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_234_LC_1_3_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_234_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_234_LC_1_3_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_234_LC_1_3_6  (
            .in0(N__21735),
            .in1(N__19784),
            .in2(N__19102),
            .in3(N__19098),
            .lcout(\ALU.madd_234 ),
            .ltout(\ALU.madd_234_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_248_LC_1_3_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_248_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_248_LC_1_3_7 .LUT_INIT=16'b1111101011101000;
    LogicCell40 \ALU.mult_madd_248_LC_1_3_7  (
            .in0(N__19697),
            .in1(N__19663),
            .in2(N__19168),
            .in3(N__19710),
            .lcout(\ALU.madd_308_0_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a7_b_8_LC_1_4_0 .C_ON=1'b0;
    defparam \ALU.mult_a7_b_8_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a7_b_8_LC_1_4_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a7_b_8_LC_1_4_0  (
            .in0(N__46433),
            .in1(N__23107),
            .in2(N__32278),
            .in3(N__30723),
            .lcout(),
            .ltout(\ALU.a7_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_9_LC_1_4_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_9_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_9_LC_1_4_1 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_490_9_LC_1_4_1  (
            .in0(N__19162),
            .in1(N__43631),
            .in2(N__19165),
            .in3(N__52199),
            .lcout(\ALU.madd_490_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_3_LC_1_4_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_3_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_3_LC_1_4_2 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.mult_madd_490_3_LC_1_4_2  (
            .in0(N__46795),
            .in1(N__44783),
            .in2(N__47071),
            .in3(N__46139),
            .lcout(\ALU.madd_490_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_1_LC_1_4_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_1_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_1_LC_1_4_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_490_1_LC_1_4_3  (
            .in0(N__43950),
            .in1(N__41570),
            .in2(N__45249),
            .in3(N__51810),
            .lcout(\ALU.madd_490_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_170_LC_1_4_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_170_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_170_LC_1_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_170_LC_1_4_4  (
            .in0(N__46793),
            .in1(N__46135),
            .in2(N__52254),
            .in3(N__43949),
            .lcout(\ALU.madd_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_171_0_tz_LC_1_4_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_171_0_tz_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_171_0_tz_LC_1_4_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_171_0_tz_LC_1_4_5  (
            .in0(N__43948),
            .in1(N__52198),
            .in2(N__46189),
            .in3(N__46794),
            .lcout(\ALU.madd_171_0_tz ),
            .ltout(\ALU.madd_171_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_171_x_LC_1_4_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_171_x_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_171_x_LC_1_4_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \ALU.mult_madd_171_x_LC_1_4_6  (
            .in0(N__51809),
            .in1(_gnd_net_),
            .in2(N__19156),
            .in3(N__38017),
            .lcout(),
            .ltout(\ALU.madd_171_x_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_229_LC_1_4_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_229_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_229_LC_1_4_7 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \ALU.mult_madd_229_LC_1_4_7  (
            .in0(N__19153),
            .in1(N__19179),
            .in2(N__19147),
            .in3(N__19920),
            .lcout(\ALU.madd_229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a8_b_5_LC_1_5_0 .C_ON=1'b0;
    defparam \ALU.mult_a8_b_5_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a8_b_5_LC_1_5_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a8_b_5_LC_1_5_0  (
            .in0(N__45194),
            .in1(N__23410),
            .in2(N__36763),
            .in3(N__30622),
            .lcout(\ALU.a8_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_171_LC_1_5_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_171_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_171_LC_1_5_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_madd_171_LC_1_5_1  (
            .in0(N__51811),
            .in1(N__19192),
            .in2(N__22066),
            .in3(N__37896),
            .lcout(),
            .ltout(\ALU.madd_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_233_LC_1_5_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_233_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_233_LC_1_5_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_233_LC_1_5_2  (
            .in0(N__19180),
            .in1(_gnd_net_),
            .in2(N__19186),
            .in3(N__19921),
            .lcout(\ALU.madd_233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_378_0_LC_1_5_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_378_0_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_378_0_LC_1_5_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_378_0_LC_1_5_3  (
            .in0(N__43376),
            .in1(N__46456),
            .in2(N__43666),
            .in3(N__46188),
            .lcout(\ALU.madd_378_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_315_0_tz_LC_1_5_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_315_0_tz_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_315_0_tz_LC_1_5_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \ALU.mult_madd_315_0_tz_LC_1_5_4  (
            .in0(N__40987),
            .in1(N__43937),
            .in2(N__41364),
            .in3(N__46805),
            .lcout(),
            .ltout(\ALU.madd_315_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_315_0_LC_1_5_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_315_0_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_315_0_LC_1_5_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \ALU.mult_madd_315_0_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__41566),
            .in2(N__19183),
            .in3(N__37895),
            .lcout(\ALU.madd_315_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_214_LC_1_5_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_214_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_214_LC_1_5_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALU.mult_madd_214_LC_1_5_6  (
            .in0(N__45195),
            .in1(N__24415),
            .in2(_gnd_net_),
            .in3(N__43375),
            .lcout(\ALU.madd_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_314_LC_1_5_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_314_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_314_LC_1_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_314_LC_1_5_7  (
            .in0(N__46806),
            .in1(N__41339),
            .in2(N__43954),
            .in3(N__40988),
            .lcout(\ALU.madd_181_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_297_LC_1_6_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_297_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_297_LC_1_6_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \ALU.mult_madd_297_LC_1_6_0  (
            .in0(N__20885),
            .in1(N__21009),
            .in2(N__21043),
            .in3(N__22231),
            .lcout(\ALU.madd_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_311_LC_1_6_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_311_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_311_LC_1_6_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ALU.mult_madd_311_LC_1_6_1  (
            .in0(N__46807),
            .in1(_gnd_net_),
            .in2(N__41365),
            .in3(N__24445),
            .lcout(\ALU.madd_311 ),
            .ltout(\ALU.madd_311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_340_LC_1_6_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_340_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_340_LC_1_6_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_340_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__19213),
            .in2(N__19231),
            .in3(N__19228),
            .lcout(\ALU.madd_340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_268_LC_1_6_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_268_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_268_LC_1_6_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_268_LC_1_6_3  (
            .in0(N__22207),
            .in1(N__23256),
            .in2(_gnd_net_),
            .in3(N__21210),
            .lcout(\ALU.madd_268 ),
            .ltout(\ALU.madd_268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_336_LC_1_6_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_336_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_336_LC_1_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_336_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__19212),
            .in2(N__19222),
            .in3(N__19219),
            .lcout(\ALU.madd_336_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_316_LC_1_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_316_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_316_LC_1_6_5 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_316_LC_1_6_5  (
            .in0(N__19203),
            .in1(N__51742),
            .in2(N__23196),
            .in3(N__44344),
            .lcout(\ALU.madd_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_298_0_LC_1_6_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_298_0_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_298_0_LC_1_6_6 .LUT_INIT=16'b1010001010101000;
    LogicCell40 \ALU.mult_madd_298_0_LC_1_6_6  (
            .in0(N__20907),
            .in1(N__21010),
            .in2(N__20892),
            .in3(N__21079),
            .lcout(\ALU.madd_298_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_320_LC_1_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_320_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_320_LC_1_6_7 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_320_LC_1_6_7  (
            .in0(N__19204),
            .in1(N__51743),
            .in2(N__23197),
            .in3(N__44345),
            .lcout(\ALU.madd_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_330_LC_1_7_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_330_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_330_LC_1_7_0 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \ALU.mult_madd_330_LC_1_7_0  (
            .in0(N__20158),
            .in1(N__47352),
            .in2(N__20152),
            .in3(N__42843),
            .lcout(\ALU.madd_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a1_b_13_LC_1_7_1 .C_ON=1'b0;
    defparam \ALU.mult_a1_b_13_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a1_b_13_LC_1_7_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a1_b_13_LC_1_7_1  (
            .in0(N__35374),
            .in1(N__31655),
            .in2(N__32202),
            .in3(N__31741),
            .lcout(\ALU.a1_b_13 ),
            .ltout(\ALU.a1_b_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_388_LC_1_7_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_388_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_388_LC_1_7_2 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_388_LC_1_7_2  (
            .in0(N__39863),
            .in1(N__22159),
            .in2(N__19195),
            .in3(N__48391),
            .lcout(\ALU.madd_388 ),
            .ltout(\ALU.madd_388_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_403_LC_1_7_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_403_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_403_LC_1_7_3 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \ALU.mult_madd_403_LC_1_7_3  (
            .in0(N__20286),
            .in1(N__19284),
            .in2(N__19255),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ALU.madd_403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_417_LC_1_7_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_417_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_417_LC_1_7_4 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_madd_417_LC_1_7_4  (
            .in0(N__27280),
            .in1(N__20407),
            .in2(N__19252),
            .in3(N__21672),
            .lcout(\ALU.madd_417 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_392_LC_1_7_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_392_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_392_LC_1_7_5 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_392_LC_1_7_5  (
            .in0(N__48390),
            .in1(N__39862),
            .in2(N__19249),
            .in3(N__22158),
            .lcout(\ALU.madd_392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_403_0_LC_1_7_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_403_0_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_403_0_LC_1_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_403_0_LC_1_7_6  (
            .in0(N__22157),
            .in1(N__20068),
            .in2(_gnd_net_),
            .in3(N__20285),
            .lcout(),
            .ltout(\ALU.madd_403_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_413_0_LC_1_7_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_413_0_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_413_0_LC_1_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_413_0_LC_1_7_7  (
            .in0(N__20406),
            .in1(N__19283),
            .in2(N__19240),
            .in3(N__27279),
            .lcout(\ALU.madd_413_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIS0G71_2_LC_1_8_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIS0G71_2_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIS0G71_2_LC_1_8_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r2_RNIS0G71_2_LC_1_8_0  (
            .in0(N__23378),
            .in1(N__25012),
            .in2(N__23361),
            .in3(N__31096),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIBF8D2_2_LC_1_8_1 .C_ON=1'b0;
    defparam \ALU.r6_RNIBF8D2_2_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIBF8D2_2_LC_1_8_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIBF8D2_2_LC_1_8_1  (
            .in0(N__28089),
            .in1(N__39167),
            .in2(N__19237),
            .in3(N__30926),
            .lcout(\ALU.r6_RNIBF8D2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_2_LC_1_8_2 .C_ON=1'b0;
    defparam \ALU.r2_2_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_2_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_2_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40296),
            .lcout(r2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56279),
            .ce(N__47712),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_2_LC_1_8_3.C_ON=1'b0;
    defparam TXbuffer_RNO_4_2_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_2_LC_1_8_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_4_2_LC_1_8_3 (
            .in0(N__30040),
            .in1(N__22390),
            .in2(N__30387),
            .in3(N__23357),
            .lcout(),
            .ltout(TXbuffer_18_13_ns_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_2_LC_1_8_4.C_ON=1'b0;
    defparam TXbuffer_RNO_1_2_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_2_LC_1_8_4.LUT_INIT=16'b1100101100001011;
    LogicCell40 TXbuffer_RNO_1_2_LC_1_8_4 (
            .in0(N__22684),
            .in1(N__30041),
            .in2(N__19234),
            .in3(N__28090),
            .lcout(TXbuffer_RNO_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_2_LC_1_8_5.C_ON=1'b0;
    defparam TXbuffer_RNO_8_2_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_2_LC_1_8_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_8_2_LC_1_8_5 (
            .in0(N__30042),
            .in1(N__22297),
            .in2(N__30388),
            .in3(N__23379),
            .lcout(),
            .ltout(TXbuffer_18_6_ns_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_2_LC_1_8_6.C_ON=1'b0;
    defparam TXbuffer_RNO_6_2_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_2_LC_1_8_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 TXbuffer_RNO_6_2_LC_1_8_6 (
            .in0(N__39168),
            .in1(N__30043),
            .in2(N__19333),
            .in3(N__22572),
            .lcout(),
            .ltout(TXbuffer_RNO_6Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_2_LC_1_8_7.C_ON=1'b0;
    defparam TXbuffer_RNO_2_2_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_2_LC_1_8_7.LUT_INIT=16'b0011001100011101;
    LogicCell40 TXbuffer_RNO_2_2_LC_1_8_7 (
            .in0(N__22603),
            .in1(N__29670),
            .in2(N__19330),
            .in3(N__49932),
            .lcout(TXbuffer_18_15_ns_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_1_0_LC_1_9_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_1_0_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_1_0_LC_1_9_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.mult_madd_490_1_0_LC_1_9_0  (
            .in0(N__19264),
            .in1(N__19270),
            .in2(_gnd_net_),
            .in3(N__19957),
            .lcout(),
            .ltout(\ALU.madd_490_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_LC_1_9_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_LC_1_9_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \ALU.mult_madd_490_LC_1_9_1  (
            .in0(N__20107),
            .in1(N__19327),
            .in2(N__19318),
            .in3(N__20320),
            .lcout(\ALU.madd_340_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_402_LC_1_9_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_402_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_402_LC_1_9_2 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \ALU.mult_madd_402_LC_1_9_2  (
            .in0(N__20359),
            .in1(N__20425),
            .in2(N__19315),
            .in3(N__24511),
            .lcout(),
            .ltout(\ALU.madd_402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_21_LC_1_9_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_21_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_21_LC_1_9_3 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \ALU.mult_madd_490_21_LC_1_9_3  (
            .in0(N__20290),
            .in1(N__19300),
            .in2(N__19291),
            .in3(N__19288),
            .lcout(\ALU.madd_490_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_397_LC_1_9_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_397_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_397_LC_1_9_4 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \ALU.mult_madd_397_LC_1_9_4  (
            .in0(N__19978),
            .in1(N__21790),
            .in2(N__20020),
            .in3(N__19998),
            .lcout(\ALU.madd_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r3_2_LC_1_10_0 .C_ON=1'b0;
    defparam \ALU.r3_2_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_2_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_2_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40300),
            .lcout(r3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56287),
            .ce(N__47763),
            .sr(_gnd_net_));
    defparam \ALU.r3_3_LC_1_10_1 .C_ON=1'b0;
    defparam \ALU.r3_3_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_3_LC_1_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_3_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50199),
            .lcout(r3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56287),
            .ce(N__47763),
            .sr(_gnd_net_));
    defparam \ALU.mult_a6_b_9_LC_1_11_0 .C_ON=1'b0;
    defparam \ALU.mult_a6_b_9_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a6_b_9_LC_1_11_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a6_b_9_LC_1_11_0  (
            .in0(N__47425),
            .in1(N__26513),
            .in2(N__36767),
            .in3(N__26449),
            .lcout(),
            .ltout(\ALU.a6_b_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_10_LC_1_11_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_10_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_10_LC_1_11_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_490_10_LC_1_11_1  (
            .in0(N__40113),
            .in1(N__31954),
            .in2(N__19357),
            .in3(N__38021),
            .lcout(),
            .ltout(\ALU.madd_490_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_13_LC_1_11_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_13_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_13_LC_1_11_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_490_13_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19354),
            .in3(N__19348),
            .lcout(\ALU.madd_490_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_7_LC_1_11_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_7_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_7_LC_1_11_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_490_7_LC_1_11_3  (
            .in0(N__39925),
            .in1(N__49013),
            .in2(N__47139),
            .in3(N__48613),
            .lcout(),
            .ltout(\ALU.madd_490_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_11_LC_1_11_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_11_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_11_LC_1_11_4 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_490_11_LC_1_11_4  (
            .in0(N__39837),
            .in1(N__19342),
            .in2(N__19351),
            .in3(N__49418),
            .lcout(\ALU.madd_490_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_13_LC_1_11_5 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_13_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_13_LC_1_11_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a2_b_13_LC_1_11_5  (
            .in0(N__35373),
            .in1(N__32655),
            .in2(N__36766),
            .in3(N__32578),
            .lcout(\ALU.a2_b_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_0_LC_1_12_1.C_ON=1'b0;
    defparam TXbuffer_RNO_4_0_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_0_LC_1_12_1.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_4_0_LC_1_12_1 (
            .in0(N__29969),
            .in1(N__23547),
            .in2(N__30310),
            .in3(N__28838),
            .lcout(),
            .ltout(TXbuffer_18_13_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_0_LC_1_12_2.C_ON=1'b0;
    defparam TXbuffer_RNO_1_0_LC_1_12_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_0_LC_1_12_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_1_0_LC_1_12_2 (
            .in0(N__29971),
            .in1(N__27826),
            .in2(N__19336),
            .in3(N__23326),
            .lcout(TXbuffer_RNO_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_4_LC_1_12_3.C_ON=1'b0;
    defparam TXbuffer_RNO_5_4_LC_1_12_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_4_LC_1_12_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_5_4_LC_1_12_3 (
            .in0(N__29970),
            .in1(N__25452),
            .in2(N__22588),
            .in3(N__34300),
            .lcout(),
            .ltout(TXbuffer_RNO_5Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_4_LC_1_12_4.C_ON=1'b0;
    defparam TXbuffer_RNO_2_4_LC_1_12_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_4_LC_1_12_4.LUT_INIT=16'b0010001101100111;
    LogicCell40 TXbuffer_RNO_2_4_LC_1_12_4 (
            .in0(N__49937),
            .in1(N__29661),
            .in2(N__19390),
            .in3(N__25231),
            .lcout(),
            .ltout(TXbuffer_18_15_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_4_LC_1_12_5.C_ON=1'b0;
    defparam TXbuffer_4_LC_1_12_5.SEQ_MODE=4'b1000;
    defparam TXbuffer_4_LC_1_12_5.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_4_LC_1_12_5 (
            .in0(N__49939),
            .in1(N__20536),
            .in2(N__19387),
            .in3(N__19366),
            .lcout(TXbufferZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56296),
            .ce(N__56037),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_0_LC_1_12_6.C_ON=1'b0;
    defparam TXbuffer_RNO_2_0_LC_1_12_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_0_LC_1_12_6.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_2_0_LC_1_12_6 (
            .in0(N__49936),
            .in1(N__21523),
            .in2(N__29674),
            .in3(N__27655),
            .lcout(),
            .ltout(TXbuffer_18_15_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_0_LC_1_12_7.C_ON=1'b0;
    defparam TXbuffer_0_LC_1_12_7.SEQ_MODE=4'b1000;
    defparam TXbuffer_0_LC_1_12_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_0_LC_1_12_7 (
            .in0(N__49938),
            .in1(N__19384),
            .in2(N__19378),
            .in3(N__27607),
            .lcout(TXbufferZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56296),
            .ce(N__56037),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_3_LC_1_13_0.C_ON=1'b0;
    defparam TXbuffer_RNO_3_3_LC_1_13_0.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_3_LC_1_13_0.LUT_INIT=16'b0000010110111011;
    LogicCell40 TXbuffer_RNO_3_3_LC_1_13_0 (
            .in0(N__29887),
            .in1(N__33244),
            .in2(N__25212),
            .in3(N__30240),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_3_LC_1_13_1.C_ON=1'b0;
    defparam TXbuffer_RNO_0_3_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_3_LC_1_13_1.LUT_INIT=16'b1000111110000101;
    LogicCell40 TXbuffer_RNO_0_3_LC_1_13_1 (
            .in0(N__29885),
            .in1(N__33610),
            .in2(N__19375),
            .in3(N__26118),
            .lcout(),
            .ltout(TXbuffer_RNO_0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_3_LC_1_13_2.C_ON=1'b0;
    defparam TXbuffer_3_LC_1_13_2.SEQ_MODE=4'b1000;
    defparam TXbuffer_3_LC_1_13_2.LUT_INIT=16'b1010000011011101;
    LogicCell40 TXbuffer_3_LC_1_13_2 (
            .in0(N__49902),
            .in1(N__19414),
            .in2(N__19372),
            .in3(N__24844),
            .lcout(TXbufferZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56300),
            .ce(N__56036),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_4_LC_1_13_5.C_ON=1'b0;
    defparam TXbuffer_RNO_3_4_LC_1_13_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_4_LC_1_13_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_3_4_LC_1_13_5 (
            .in0(N__29884),
            .in1(N__25171),
            .in2(N__30304),
            .in3(N__33478),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_4_LC_1_13_6.C_ON=1'b0;
    defparam TXbuffer_RNO_0_4_LC_1_13_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_4_LC_1_13_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_0_4_LC_1_13_6 (
            .in0(N__29886),
            .in1(N__26083),
            .in2(N__19369),
            .in3(N__33574),
            .lcout(TXbuffer_RNO_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXstart_LC_1_14_1.C_ON=1'b0;
    defparam TXstart_LC_1_14_1.SEQ_MODE=4'b1000;
    defparam TXstart_LC_1_14_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 TXstart_LC_1_14_1 (
            .in0(N__27075),
            .in1(N__26976),
            .in2(N__27015),
            .in3(N__27051),
            .lcout(TXstartZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56302),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI7AQC9_0_15_LC_1_14_4 .C_ON=1'b0;
    defparam \ALU.r2_RNI7AQC9_0_15_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI7AQC9_0_15_LC_1_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.r2_RNI7AQC9_0_15_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__40084),
            .in2(_gnd_net_),
            .in3(N__39973),
            .lcout(\ALU.r2_RNI7AQC9_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_3_LC_1_14_5.C_ON=1'b0;
    defparam TXbuffer_RNO_1_3_LC_1_14_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_3_LC_1_14_5.LUT_INIT=16'b1000100011110101;
    LogicCell40 TXbuffer_RNO_1_3_LC_1_14_5 (
            .in0(N__29859),
            .in1(N__28060),
            .in2(N__22651),
            .in3(N__20503),
            .lcout(TXbuffer_RNO_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_0_LC_1_15_0.C_ON=1'b1;
    defparam clkdiv_0_LC_1_15_0.SEQ_MODE=4'b1000;
    defparam clkdiv_0_LC_1_15_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_0_LC_1_15_0 (
            .in0(_gnd_net_),
            .in1(N__26975),
            .in2(_gnd_net_),
            .in3(N__19408),
            .lcout(clkdivZ0Z_0),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(clkdiv_cry_0),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_1_LC_1_15_1.C_ON=1'b1;
    defparam clkdiv_1_LC_1_15_1.SEQ_MODE=4'b1000;
    defparam clkdiv_1_LC_1_15_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_1_LC_1_15_1 (
            .in0(_gnd_net_),
            .in1(N__27074),
            .in2(_gnd_net_),
            .in3(N__19405),
            .lcout(clkdivZ0Z_1),
            .ltout(),
            .carryin(clkdiv_cry_0),
            .carryout(clkdiv_cry_1),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_2_LC_1_15_2.C_ON=1'b1;
    defparam clkdiv_2_LC_1_15_2.SEQ_MODE=4'b1000;
    defparam clkdiv_2_LC_1_15_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_2_LC_1_15_2 (
            .in0(_gnd_net_),
            .in1(N__27050),
            .in2(_gnd_net_),
            .in3(N__19402),
            .lcout(clkdivZ0Z_2),
            .ltout(),
            .carryin(clkdiv_cry_1),
            .carryout(clkdiv_cry_2),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_3_LC_1_15_3.C_ON=1'b1;
    defparam clkdiv_3_LC_1_15_3.SEQ_MODE=4'b1000;
    defparam clkdiv_3_LC_1_15_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_3_LC_1_15_3 (
            .in0(_gnd_net_),
            .in1(N__27008),
            .in2(_gnd_net_),
            .in3(N__19399),
            .lcout(clkdivZ0Z_3),
            .ltout(),
            .carryin(clkdiv_cry_2),
            .carryout(clkdiv_cry_3),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_4_LC_1_15_4.C_ON=1'b1;
    defparam clkdiv_4_LC_1_15_4.SEQ_MODE=4'b1000;
    defparam clkdiv_4_LC_1_15_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_4_LC_1_15_4 (
            .in0(_gnd_net_),
            .in1(N__49853),
            .in2(_gnd_net_),
            .in3(N__19396),
            .lcout(clkdivZ0Z_4),
            .ltout(),
            .carryin(clkdiv_cry_3),
            .carryout(clkdiv_cry_4),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_5_LC_1_15_5.C_ON=1'b1;
    defparam clkdiv_5_LC_1_15_5.SEQ_MODE=4'b1000;
    defparam clkdiv_5_LC_1_15_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_5_LC_1_15_5 (
            .in0(_gnd_net_),
            .in1(N__29622),
            .in2(_gnd_net_),
            .in3(N__19393),
            .lcout(clkdivZ0Z_5),
            .ltout(),
            .carryin(clkdiv_cry_4),
            .carryout(clkdiv_cry_5),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_6_LC_1_15_6.C_ON=1'b1;
    defparam clkdiv_6_LC_1_15_6.SEQ_MODE=4'b1000;
    defparam clkdiv_6_LC_1_15_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_6_LC_1_15_6 (
            .in0(_gnd_net_),
            .in1(N__29842),
            .in2(_gnd_net_),
            .in3(N__19474),
            .lcout(clkdivZ0Z_6),
            .ltout(),
            .carryin(clkdiv_cry_5),
            .carryout(clkdiv_cry_6),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_7_LC_1_15_7.C_ON=1'b1;
    defparam clkdiv_7_LC_1_15_7.SEQ_MODE=4'b1000;
    defparam clkdiv_7_LC_1_15_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_7_LC_1_15_7 (
            .in0(_gnd_net_),
            .in1(N__30209),
            .in2(_gnd_net_),
            .in3(N__19471),
            .lcout(clkdivZ0Z_7),
            .ltout(),
            .carryin(clkdiv_cry_6),
            .carryout(clkdiv_cry_7),
            .clk(N__56303),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_8_LC_1_16_0.C_ON=1'b1;
    defparam clkdiv_8_LC_1_16_0.SEQ_MODE=4'b1000;
    defparam clkdiv_8_LC_1_16_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_8_LC_1_16_0 (
            .in0(_gnd_net_),
            .in1(N__19468),
            .in2(_gnd_net_),
            .in3(N__19462),
            .lcout(clkdivZ0Z_8),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(clkdiv_cry_8),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_9_LC_1_16_1.C_ON=1'b1;
    defparam clkdiv_9_LC_1_16_1.SEQ_MODE=4'b1000;
    defparam clkdiv_9_LC_1_16_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_9_LC_1_16_1 (
            .in0(_gnd_net_),
            .in1(N__19459),
            .in2(_gnd_net_),
            .in3(N__19453),
            .lcout(clkdivZ0Z_9),
            .ltout(),
            .carryin(clkdiv_cry_8),
            .carryout(clkdiv_cry_9),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_10_LC_1_16_2.C_ON=1'b1;
    defparam clkdiv_10_LC_1_16_2.SEQ_MODE=4'b1000;
    defparam clkdiv_10_LC_1_16_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_10_LC_1_16_2 (
            .in0(_gnd_net_),
            .in1(N__19450),
            .in2(_gnd_net_),
            .in3(N__19444),
            .lcout(clkdivZ0Z_10),
            .ltout(),
            .carryin(clkdiv_cry_9),
            .carryout(clkdiv_cry_10),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_11_LC_1_16_3.C_ON=1'b1;
    defparam clkdiv_11_LC_1_16_3.SEQ_MODE=4'b1000;
    defparam clkdiv_11_LC_1_16_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_11_LC_1_16_3 (
            .in0(_gnd_net_),
            .in1(N__19441),
            .in2(_gnd_net_),
            .in3(N__19435),
            .lcout(clkdivZ0Z_11),
            .ltout(),
            .carryin(clkdiv_cry_10),
            .carryout(clkdiv_cry_11),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_12_LC_1_16_4.C_ON=1'b1;
    defparam clkdiv_12_LC_1_16_4.SEQ_MODE=4'b1000;
    defparam clkdiv_12_LC_1_16_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_12_LC_1_16_4 (
            .in0(_gnd_net_),
            .in1(N__19432),
            .in2(_gnd_net_),
            .in3(N__19426),
            .lcout(clkdivZ0Z_12),
            .ltout(),
            .carryin(clkdiv_cry_11),
            .carryout(clkdiv_cry_12),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_13_LC_1_16_5.C_ON=1'b1;
    defparam clkdiv_13_LC_1_16_5.SEQ_MODE=4'b1000;
    defparam clkdiv_13_LC_1_16_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_13_LC_1_16_5 (
            .in0(_gnd_net_),
            .in1(N__19423),
            .in2(_gnd_net_),
            .in3(N__19417),
            .lcout(clkdivZ0Z_13),
            .ltout(),
            .carryin(clkdiv_cry_12),
            .carryout(clkdiv_cry_13),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_14_LC_1_16_6.C_ON=1'b1;
    defparam clkdiv_14_LC_1_16_6.SEQ_MODE=4'b1000;
    defparam clkdiv_14_LC_1_16_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_14_LC_1_16_6 (
            .in0(_gnd_net_),
            .in1(N__19555),
            .in2(_gnd_net_),
            .in3(N__19549),
            .lcout(clkdivZ0Z_14),
            .ltout(),
            .carryin(clkdiv_cry_13),
            .carryout(clkdiv_cry_14),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_15_LC_1_16_7.C_ON=1'b1;
    defparam clkdiv_15_LC_1_16_7.SEQ_MODE=4'b1000;
    defparam clkdiv_15_LC_1_16_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_15_LC_1_16_7 (
            .in0(_gnd_net_),
            .in1(N__19546),
            .in2(_gnd_net_),
            .in3(N__19540),
            .lcout(clkdivZ0Z_15),
            .ltout(),
            .carryin(clkdiv_cry_14),
            .carryout(clkdiv_cry_15),
            .clk(N__56304),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_16_LC_1_17_0.C_ON=1'b1;
    defparam clkdiv_16_LC_1_17_0.SEQ_MODE=4'b1000;
    defparam clkdiv_16_LC_1_17_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_16_LC_1_17_0 (
            .in0(_gnd_net_),
            .in1(N__19537),
            .in2(_gnd_net_),
            .in3(N__19531),
            .lcout(clkdivZ0Z_16),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(clkdiv_cry_16),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_17_LC_1_17_1.C_ON=1'b1;
    defparam clkdiv_17_LC_1_17_1.SEQ_MODE=4'b1000;
    defparam clkdiv_17_LC_1_17_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_17_LC_1_17_1 (
            .in0(_gnd_net_),
            .in1(N__19528),
            .in2(_gnd_net_),
            .in3(N__19522),
            .lcout(clkdivZ0Z_17),
            .ltout(),
            .carryin(clkdiv_cry_16),
            .carryout(clkdiv_cry_17),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_18_LC_1_17_2.C_ON=1'b1;
    defparam clkdiv_18_LC_1_17_2.SEQ_MODE=4'b1000;
    defparam clkdiv_18_LC_1_17_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_18_LC_1_17_2 (
            .in0(_gnd_net_),
            .in1(N__19519),
            .in2(_gnd_net_),
            .in3(N__19513),
            .lcout(clkdivZ0Z_18),
            .ltout(),
            .carryin(clkdiv_cry_17),
            .carryout(clkdiv_cry_18),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_19_LC_1_17_3.C_ON=1'b1;
    defparam clkdiv_19_LC_1_17_3.SEQ_MODE=4'b1000;
    defparam clkdiv_19_LC_1_17_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_19_LC_1_17_3 (
            .in0(_gnd_net_),
            .in1(N__19510),
            .in2(_gnd_net_),
            .in3(N__19504),
            .lcout(clkdivZ0Z_19),
            .ltout(),
            .carryin(clkdiv_cry_18),
            .carryout(clkdiv_cry_19),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_20_LC_1_17_4.C_ON=1'b1;
    defparam clkdiv_20_LC_1_17_4.SEQ_MODE=4'b1000;
    defparam clkdiv_20_LC_1_17_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_20_LC_1_17_4 (
            .in0(_gnd_net_),
            .in1(N__19501),
            .in2(_gnd_net_),
            .in3(N__19495),
            .lcout(clkdivZ0Z_20),
            .ltout(),
            .carryin(clkdiv_cry_19),
            .carryout(clkdiv_cry_20),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_21_LC_1_17_5.C_ON=1'b1;
    defparam clkdiv_21_LC_1_17_5.SEQ_MODE=4'b1000;
    defparam clkdiv_21_LC_1_17_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_21_LC_1_17_5 (
            .in0(_gnd_net_),
            .in1(N__19492),
            .in2(_gnd_net_),
            .in3(N__19486),
            .lcout(clkdivZ0Z_21),
            .ltout(),
            .carryin(clkdiv_cry_20),
            .carryout(clkdiv_cry_21),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_22_LC_1_17_6.C_ON=1'b1;
    defparam clkdiv_22_LC_1_17_6.SEQ_MODE=4'b1000;
    defparam clkdiv_22_LC_1_17_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_22_LC_1_17_6 (
            .in0(_gnd_net_),
            .in1(N__19483),
            .in2(_gnd_net_),
            .in3(N__19477),
            .lcout(clkdivZ0Z_22),
            .ltout(),
            .carryin(clkdiv_cry_21),
            .carryout(clkdiv_cry_22),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_23_LC_1_17_7.C_ON=1'b0;
    defparam clkdiv_23_LC_1_17_7.SEQ_MODE=4'b1000;
    defparam clkdiv_23_LC_1_17_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 clkdiv_23_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(N__19593),
            .in2(_gnd_net_),
            .in3(N__19603),
            .lcout(GPIO3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56305),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_154_LC_2_1_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_154_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_154_LC_2_1_0 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \ALU.mult_madd_154_LC_2_1_0  (
            .in0(N__22841),
            .in1(N__21871),
            .in2(N__31575),
            .in3(N__21549),
            .lcout(\ALU.madd_154 ),
            .ltout(\ALU.madd_154_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_LC_2_1_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_LC_2_1_1 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_g0_0_LC_2_1_1  (
            .in0(N__19885),
            .in1(N__23128),
            .in2(N__19582),
            .in3(N__19642),
            .lcout(),
            .ltout(\ALU.N_703_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_LC_2_1_2 .C_ON=1'b0;
    defparam \ALU.mult_g0_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_LC_2_1_2 .LUT_INIT=16'b1110000100011110;
    LogicCell40 \ALU.mult_g0_LC_2_1_2  (
            .in0(N__19669),
            .in1(N__19711),
            .in2(N__19579),
            .in3(N__19726),
            .lcout(),
            .ltout(\ALU.g0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_10_LC_2_1_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_10_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_10_LC_2_1_3 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_axb_10_LC_2_1_3  (
            .in0(N__19572),
            .in1(N__26319),
            .in2(N__19576),
            .in3(N__26304),
            .lcout(\ALU.madd_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_150_LC_2_1_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_150_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_150_LC_2_1_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_150_LC_2_1_4  (
            .in0(N__22842),
            .in1(N__21872),
            .in2(N__31576),
            .in3(N__21550),
            .lcout(\ALU.madd_150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_206_LC_2_1_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_206_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_206_LC_2_1_5 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_madd_206_LC_2_1_5  (
            .in0(N__20689),
            .in1(N__19767),
            .in2(N__20584),
            .in3(N__19720),
            .lcout(\ALU.madd_206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_202_LC_2_1_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_202_LC_2_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_202_LC_2_1_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_202_LC_2_1_6  (
            .in0(N__19719),
            .in1(N__20580),
            .in2(N__19768),
            .in3(N__20688),
            .lcout(\ALU.madd_334 ),
            .ltout(\ALU.madd_334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_13_LC_2_1_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_13_LC_2_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_13_LC_2_1_7 .LUT_INIT=16'b1110101010000000;
    LogicCell40 \ALU.mult_g0_13_LC_2_1_7  (
            .in0(N__19573),
            .in1(N__20602),
            .in2(N__19564),
            .in3(N__19561),
            .lcout(\ALU.g0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_192_0_LC_2_2_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_192_0_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_192_0_LC_2_2_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_192_0_LC_2_2_0  (
            .in0(N__19815),
            .in1(_gnd_net_),
            .in2(N__47269),
            .in3(N__24394),
            .lcout(\ALU.madd_192_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_144_LC_2_2_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_144_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_144_LC_2_2_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ALU.mult_madd_144_LC_2_2_1  (
            .in0(N__21883),
            .in1(N__22888),
            .in2(N__43649),
            .in3(N__49361),
            .lcout(\ALU.madd_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_3_LC_2_2_2 .C_ON=1'b0;
    defparam \ALU.mult_g0_3_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_3_LC_2_2_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_3_LC_2_2_2  (
            .in0(N__19744),
            .in1(N__19698),
            .in2(N__19738),
            .in3(N__20639),
            .lcout(\ALU.g0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_197_LC_2_2_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_197_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_197_LC_2_2_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_197_LC_2_2_3  (
            .in0(N__19640),
            .in1(N__19620),
            .in2(N__19883),
            .in3(N__19611),
            .lcout(\ALU.madd_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_195_LC_2_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_195_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_195_LC_2_2_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_madd_195_LC_2_2_4  (
            .in0(N__19813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20686),
            .lcout(\ALU.madd_112 ),
            .ltout(\ALU.madd_112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_244_LC_2_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_244_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_244_LC_2_2_5 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ALU.mult_madd_244_LC_2_2_5  (
            .in0(N__19699),
            .in1(N__19681),
            .in2(N__19672),
            .in3(N__19664),
            .lcout(\ALU.madd_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_196_0_LC_2_2_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_196_0_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_196_0_LC_2_2_6 .LUT_INIT=16'b0011110000101000;
    LogicCell40 \ALU.mult_madd_196_0_LC_2_2_6  (
            .in0(N__19814),
            .in1(N__24393),
            .in2(N__47268),
            .in3(N__20687),
            .lcout(\ALU.madd_196_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_201_LC_2_2_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_201_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_201_LC_2_2_7 .LUT_INIT=16'b1000111011101000;
    LogicCell40 \ALU.mult_madd_201_LC_2_2_7  (
            .in0(N__19641),
            .in1(N__19621),
            .in2(N__19884),
            .in3(N__19612),
            .lcout(\ALU.madd_201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_239_LC_2_3_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_239_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_239_LC_2_3_0 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ALU.mult_madd_239_LC_2_3_0  (
            .in0(N__20748),
            .in1(N__19797),
            .in2(N__23164),
            .in3(N__20730),
            .lcout(\ALU.madd_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g2_0_1_LC_2_3_1 .C_ON=1'b0;
    defparam \ALU.mult_g2_0_1_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g2_0_1_LC_2_3_1 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_g2_0_1_LC_2_3_1  (
            .in0(N__51988),
            .in1(N__48928),
            .in2(N__47457),
            .in3(N__48570),
            .lcout(\ALU.g2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_182_0_LC_2_3_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_182_0_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_182_0_LC_2_3_2 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_182_0_LC_2_3_2  (
            .in0(N__48569),
            .in1(N__47423),
            .in2(N__48988),
            .in3(N__51987),
            .lcout(\ALU.madd_182_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_0_LC_2_3_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_0_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_0_LC_2_3_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_axb_0_LC_2_3_3  (
            .in0(N__38020),
            .in1(N__48571),
            .in2(N__46823),
            .in3(N__48932),
            .lcout(\ALU.mult_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_177_LC_2_3_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_177_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_177_LC_2_3_4 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_177_LC_2_3_4  (
            .in0(N__42753),
            .in1(N__19854),
            .in2(N__19837),
            .in3(N__43635),
            .lcout(\ALU.madd_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_243_LC_2_3_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_243_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_243_LC_2_3_5 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \ALU.mult_madd_243_LC_2_3_5  (
            .in0(N__19798),
            .in1(N__23163),
            .in2(N__20734),
            .in3(N__20749),
            .lcout(\ALU.madd_243 ),
            .ltout(\ALU.madd_243_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_299_LC_2_3_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_299_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_299_LC_2_3_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_299_LC_2_3_6  (
            .in0(N__21183),
            .in1(N__20770),
            .in2(N__19789),
            .in3(N__22871),
            .lcout(\ALU.madd_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_219_0_LC_2_3_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_219_0_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_219_0_LC_2_3_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_219_0_LC_2_3_7  (
            .in0(N__44766),
            .in1(N__45461),
            .in2(N__43664),
            .in3(N__42752),
            .lcout(\ALU.madd_219_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_304_LC_2_4_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_304_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_304_LC_2_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_304_LC_2_4_0  (
            .in0(N__20865),
            .in1(N__19944),
            .in2(_gnd_net_),
            .in3(N__19929),
            .lcout(\ALU.madd_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_303_0_LC_2_4_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_303_0_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_303_0_LC_2_4_1 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \ALU.mult_madd_303_0_LC_2_4_1  (
            .in0(N__22873),
            .in1(N__20769),
            .in2(N__21187),
            .in3(N__19909),
            .lcout(\ALU.madd_303_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_293_LC_2_4_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_293_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_293_LC_2_4_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_293_LC_2_4_2  (
            .in0(N__20794),
            .in1(_gnd_net_),
            .in2(N__20788),
            .in3(N__20970),
            .lcout(\ALU.madd_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_393_LC_2_4_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_393_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_393_LC_2_4_3 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \ALU.mult_madd_393_LC_2_4_3  (
            .in0(N__20013),
            .in1(N__21786),
            .in2(N__20002),
            .in3(N__19977),
            .lcout(\ALU.madd_393 ),
            .ltout(\ALU.madd_393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_412_LC_2_4_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_412_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_412_LC_2_4_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_412_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__20047),
            .in2(N__19960),
            .in3(N__20923),
            .lcout(\ALU.madd_412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_308_LC_2_4_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_308_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_308_LC_2_4_5 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_308_LC_2_4_5  (
            .in0(N__19945),
            .in1(_gnd_net_),
            .in2(N__19933),
            .in3(N__20866),
            .lcout(\ALU.madd_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_209_LC_2_4_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_209_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_209_LC_2_4_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALU.mult_madd_209_LC_2_4_6  (
            .in0(N__51808),
            .in1(N__23011),
            .in2(_gnd_net_),
            .in3(N__46789),
            .lcout(\ALU.madd_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_302_LC_2_4_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_302_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_302_LC_2_4_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_302_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(N__20768),
            .in2(_gnd_net_),
            .in3(N__19908),
            .lcout(\ALU.madd_175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_365_LC_2_5_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_365_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_365_LC_2_5_0 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \ALU.mult_madd_365_LC_2_5_0  (
            .in0(N__20212),
            .in1(N__20098),
            .in2(N__20092),
            .in3(N__20077),
            .lcout(\ALU.madd_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_13_LC_2_5_1 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_13_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_13_LC_2_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a0_b_13_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__35387),
            .in2(_gnd_net_),
            .in3(N__49004),
            .lcout(\ALU.a0_b_13 ),
            .ltout(\ALU.a0_b_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_331_LC_2_5_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_331_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_331_LC_2_5_2 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ALU.mult_madd_331_LC_2_5_2  (
            .in0(N__48608),
            .in1(N__39813),
            .in2(N__19900),
            .in3(N__21261),
            .lcout(\ALU.madd_331_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_356_LC_2_5_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_356_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_356_LC_2_5_3 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ALU.mult_madd_356_LC_2_5_3  (
            .in0(N__20194),
            .in1(N__20200),
            .in2(N__20820),
            .in3(N__20178),
            .lcout(\ALU.madd_356 ),
            .ltout(\ALU.madd_356_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_361_LC_2_5_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_361_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_361_LC_2_5_4 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ALU.mult_madd_361_LC_2_5_4  (
            .in0(N__20088),
            .in1(N__20211),
            .in2(N__20080),
            .in3(N__20076),
            .lcout(\ALU.madd_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_388_0_LC_2_5_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_388_0_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_388_0_LC_2_5_5 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.mult_madd_388_0_LC_2_5_5  (
            .in0(N__48365),
            .in1(N__35388),
            .in2(N__39849),
            .in3(N__48609),
            .lcout(\ALU.madd_388_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_1_c_RNO_LC_2_5_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_3_1_c_RNO_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_1_c_RNO_LC_2_5_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_3_1_c_RNO_LC_2_5_6  (
            .in0(N__55162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41823),
            .lcout(\ALU.r0_12_prm_3_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_RNO_4_LC_2_5_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_1_c_RNO_4_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_RNO_4_LC_2_5_7 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \ALU.r0_12_prm_8_1_c_RNO_4_LC_2_5_7  (
            .in0(N__48366),
            .in1(N__53516),
            .in2(N__54478),
            .in3(N__48610),
            .lcout(\ALU.rshift_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_427_LC_2_6_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_427_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_427_LC_2_6_0 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_madd_427_LC_2_6_0  (
            .in0(N__20248),
            .in1(N__20026),
            .in2(N__21673),
            .in3(N__20167),
            .lcout(\ALU.madd_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_408_LC_2_6_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_408_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_408_LC_2_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_408_LC_2_6_1  (
            .in0(N__20056),
            .in1(N__20922),
            .in2(_gnd_net_),
            .in3(N__20043),
            .lcout(\ALU.madd_408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_355_LC_2_6_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_355_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_355_LC_2_6_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_355_LC_2_6_2  (
            .in0(N__20220),
            .in1(N__20232),
            .in2(_gnd_net_),
            .in3(N__21243),
            .lcout(\ALU.madd_355 ),
            .ltout(\ALU.madd_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_418_LC_2_6_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_418_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_418_LC_2_6_3 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \ALU.mult_madd_418_LC_2_6_3  (
            .in0(N__20982),
            .in1(N__20121),
            .in2(N__20029),
            .in3(N__20134),
            .lcout(\ALU.madd_418 ),
            .ltout(\ALU.madd_418_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_423_LC_2_6_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_423_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_423_LC_2_6_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_423_LC_2_6_4  (
            .in0(N__20247),
            .in1(N__21668),
            .in2(N__20239),
            .in3(N__20166),
            .lcout(\ALU.madd_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_351_LC_2_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_351_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_351_LC_2_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_351_LC_2_6_5  (
            .in0(N__21244),
            .in1(_gnd_net_),
            .in2(N__20236),
            .in3(N__20221),
            .lcout(\ALU.madd_351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_346_LC_2_6_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_346_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_346_LC_2_6_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.mult_madd_346_LC_2_6_6  (
            .in0(N__20143),
            .in1(N__21059),
            .in2(_gnd_net_),
            .in3(N__21100),
            .lcout(\ALU.madd_346 ),
            .ltout(\ALU.madd_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_360_LC_2_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_360_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_360_LC_2_6_7 .LUT_INIT=16'b1111101011101000;
    LogicCell40 \ALU.mult_madd_360_LC_2_6_7  (
            .in0(N__20821),
            .in1(N__20193),
            .in2(N__20182),
            .in3(N__20179),
            .lcout(\ALU.madd_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_329_LC_2_7_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_329_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_329_LC_2_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_329_LC_2_7_0  (
            .in0(N__49364),
            .in1(N__51919),
            .in2(N__35540),
            .in3(N__48364),
            .lcout(\ALU.madd_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_330_0_tz_LC_2_7_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_330_0_tz_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_330_0_tz_LC_2_7_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \ALU.mult_madd_330_0_tz_LC_2_7_1  (
            .in0(N__48363),
            .in1(N__35500),
            .in2(N__51958),
            .in3(N__49365),
            .lcout(\ALU.madd_330_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_326_LC_2_7_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_326_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_326_LC_2_7_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ALU.mult_madd_326_LC_2_7_2  (
            .in0(N__35496),
            .in1(_gnd_net_),
            .in2(N__20269),
            .in3(N__48362),
            .lcout(\ALU.madd_326 ),
            .ltout(\ALU.madd_326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_350_0_LC_2_7_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_350_0_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_350_0_LC_2_7_3 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \ALU.mult_madd_350_0_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__21130),
            .in2(N__20137),
            .in3(N__21064),
            .lcout(\ALU.madd_350_0 ),
            .ltout(\ALU.madd_350_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_422_LC_2_7_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_422_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_422_LC_2_7_4 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \ALU.mult_madd_422_LC_2_7_4  (
            .in0(N__20128),
            .in1(N__20122),
            .in2(N__20110),
            .in3(N__20983),
            .lcout(\ALU.madd_422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a7_b_7_LC_2_7_5 .C_ON=1'b0;
    defparam \ALU.mult_a7_b_7_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a7_b_7_LC_2_7_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a7_b_7_LC_2_7_5  (
            .in0(N__44776),
            .in1(N__23102),
            .in2(N__32201),
            .in3(N__30722),
            .lcout(\ALU.a7_b_7 ),
            .ltout(\ALU.a7_b_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_383_LC_2_7_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_383_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_383_LC_2_7_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ALU.mult_madd_383_LC_2_7_6  (
            .in0(N__49363),
            .in1(N__35539),
            .in2(N__20293),
            .in3(N__20373),
            .lcout(\ALU.madd_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a4_b_10_LC_2_7_7 .C_ON=1'b0;
    defparam \ALU.mult_a4_b_10_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a4_b_10_LC_2_7_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a4_b_10_LC_2_7_7  (
            .in0(N__51918),
            .in1(N__32464),
            .in2(N__32200),
            .in3(N__32372),
            .lcout(\ALU.a4_b_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIU2J74_9_LC_2_8_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIU2J74_9_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIU2J74_9_LC_2_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIU2J74_9_LC_2_8_0  (
            .in0(N__24630),
            .in1(N__21306),
            .in2(_gnd_net_),
            .in3(N__21288),
            .lcout(\ALU.b_9 ),
            .ltout(\ALU.b_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_326_0_LC_2_8_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_326_0_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_326_0_LC_2_8_1 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.mult_madd_326_0_LC_2_8_1  (
            .in0(N__42842),
            .in1(N__51917),
            .in2(N__20272),
            .in3(N__49362),
            .lcout(\ALU.madd_326_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_11_LC_2_8_2 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_11_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_11_LC_2_8_2 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \ALU.mult_a3_b_11_LC_2_8_2  (
            .in0(N__35501),
            .in1(N__31921),
            .in2(N__31833),
            .in3(N__32199),
            .lcout(\ALU.a3_b_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_9_LC_2_8_3 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_9_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_9_LC_2_8_3 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \ALU.mult_a5_b_9_LC_2_8_3  (
            .in0(N__29003),
            .in1(N__29077),
            .in2(N__32237),
            .in3(N__47342),
            .lcout(\ALU.a5_b_9 ),
            .ltout(\ALU.a5_b_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_382_LC_2_8_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_382_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_382_LC_2_8_4 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_382_LC_2_8_4  (
            .in0(N__20257),
            .in1(N__43651),
            .in2(N__20260),
            .in3(N__46173),
            .lcout(\ALU.madd_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a6_b_8_LC_2_8_5 .C_ON=1'b0;
    defparam \ALU.mult_a6_b_8_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a6_b_8_LC_2_8_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a6_b_8_LC_2_8_5  (
            .in0(N__26504),
            .in1(N__26435),
            .in2(N__32238),
            .in3(N__46432),
            .lcout(\ALU.a6_b_8 ),
            .ltout(\ALU.a6_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_378_LC_2_8_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_378_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_378_LC_2_8_6 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_378_LC_2_8_6  (
            .in0(N__20421),
            .in1(N__43650),
            .in2(N__20410),
            .in3(N__46172),
            .lcout(\ALU.madd_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNILIOQ3_3_LC_2_9_0 .C_ON=1'b0;
    defparam \ALU.r4_RNILIOQ3_3_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNILIOQ3_3_LC_2_9_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.r4_RNILIOQ3_3_LC_2_9_0  (
            .in0(N__32883),
            .in1(N__24336),
            .in2(_gnd_net_),
            .in3(N__33036),
            .lcout(\ALU.b_i_3 ),
            .ltout(\ALU.b_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNINFAJC_3_LC_2_9_1 .C_ON=1'b0;
    defparam \ALU.r4_RNINFAJC_3_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNINFAJC_3_LC_2_9_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.r4_RNINFAJC_3_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20395),
            .in3(N__24307),
            .lcout(\ALU.r4_RNINFAJCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_16_LC_2_9_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_16_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_16_LC_2_9_3 .LUT_INIT=16'b0011011001101100;
    LogicCell40 \ALU.mult_madd_490_16_LC_2_9_3  (
            .in0(N__20392),
            .in1(N__20383),
            .in2(N__48061),
            .in3(N__20377),
            .lcout(\ALU.madd_490_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a11_b_3_LC_2_9_4 .C_ON=1'b0;
    defparam \ALU.mult_a11_b_3_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a11_b_3_LC_2_9_4 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a11_b_3_LC_2_9_4  (
            .in0(N__24337),
            .in1(N__33037),
            .in2(N__32895),
            .in3(N__40892),
            .lcout(\ALU.a11_b_3 ),
            .ltout(\ALU.a11_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_373_LC_2_9_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_373_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_373_LC_2_9_5 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_373_LC_2_9_5  (
            .in0(N__36486),
            .in1(N__45222),
            .in2(N__20362),
            .in3(N__52299),
            .lcout(\ALU.madd_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_15_LC_2_9_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_15_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_15_LC_2_9_6 .LUT_INIT=16'b0011011001101100;
    LogicCell40 \ALU.mult_madd_490_15_LC_2_9_6  (
            .in0(N__27306),
            .in1(N__24484),
            .in2(N__20353),
            .in3(N__36487),
            .lcout(),
            .ltout(\ALU.madd_490_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_19_LC_2_9_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_19_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_19_LC_2_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_490_19_LC_2_9_7  (
            .in0(N__20344),
            .in1(N__20329),
            .in2(N__20323),
            .in3(N__20440),
            .lcout(\ALU.madd_490_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_14_LC_2_10_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_14_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_14_LC_2_10_1 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_axb_14_LC_2_10_1  (
            .in0(N__20314),
            .in1(N__20959),
            .in2(N__20302),
            .in3(N__20944),
            .lcout(\ALU.madd_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIE0AK8_1_11_LC_2_10_2 .C_ON=1'b0;
    defparam \ALU.r5_RNIE0AK8_1_11_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIE0AK8_1_11_LC_2_10_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ALU.r5_RNIE0AK8_1_11_LC_2_10_2  (
            .in0(N__40957),
            .in1(_gnd_net_),
            .in2(N__35592),
            .in3(_gnd_net_),
            .lcout(\ALU.r5_RNIE0AK8_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIAFSR_15_LC_2_10_3 .C_ON=1'b0;
    defparam \ALU.r1_RNIAFSR_15_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIAFSR_15_LC_2_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r1_RNIAFSR_15_LC_2_10_3  (
            .in0(N__30480),
            .in1(N__30117),
            .in2(_gnd_net_),
            .in3(N__29507),
            .lcout(\ALU.r1_RNIAFSRZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_0_LC_2_10_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_0_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_0_LC_2_10_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_490_0_LC_2_10_5  (
            .in0(N__40521),
            .in1(N__44361),
            .in2(N__41362),
            .in3(N__40956),
            .lcout(),
            .ltout(\ALU.madd_490_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_14_LC_2_10_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_14_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_14_LC_2_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_490_14_LC_2_10_6  (
            .in0(N__20479),
            .in1(N__20464),
            .in2(N__20449),
            .in3(N__20446),
            .lcout(\ALU.madd_490_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNISP2L9_2_12_LC_2_10_7 .C_ON=1'b0;
    defparam \ALU.r5_RNISP2L9_2_12_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNISP2L9_2_12_LC_2_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r5_RNISP2L9_2_12_LC_2_10_7  (
            .in0(N__39826),
            .in1(_gnd_net_),
            .in2(N__41363),
            .in3(_gnd_net_),
            .lcout(\ALU.r5_RNISP2L9_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIFR6T_15_LC_2_11_1 .C_ON=1'b0;
    defparam \ALU.r2_RNIFR6T_15_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIFR6T_15_LC_2_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r2_RNIFR6T_15_LC_2_11_1  (
            .in0(N__25079),
            .in1(N__22511),
            .in2(_gnd_net_),
            .in3(N__22431),
            .lcout(),
            .ltout(\ALU.r2_RNIFR6TZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI418R4_15_LC_2_11_2 .C_ON=1'b0;
    defparam \ALU.r2_RNI418R4_15_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI418R4_15_LC_2_11_2 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \ALU.r2_RNI418R4_15_LC_2_11_2  (
            .in0(N__32892),
            .in1(N__21406),
            .in2(N__20431),
            .in3(N__20485),
            .lcout(\ALU.b_15 ),
            .ltout(\ALU.b_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_15_s1_c_RNO_LC_2_11_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_15_s1_c_RNO_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_15_s1_c_RNO_LC_2_11_3 .LUT_INIT=16'b1010010101010101;
    LogicCell40 \ALU.r0_12_prm_7_15_s1_c_RNO_LC_2_11_3  (
            .in0(N__53254),
            .in1(_gnd_net_),
            .in2(N__20428),
            .in3(N__40114),
            .lcout(\ALU.r0_12_prm_7_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_7_LC_2_11_4.C_ON=1'b0;
    defparam TXbuffer_RNO_4_7_LC_2_11_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_7_LC_2_11_4.LUT_INIT=16'b0001000111001111;
    LogicCell40 TXbuffer_RNO_4_7_LC_2_11_4 (
            .in0(N__22512),
            .in1(N__29975),
            .in2(N__22486),
            .in3(N__30281),
            .lcout(TXbuffer_18_13_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_3_LC_2_11_5.C_ON=1'b0;
    defparam TXbuffer_RNO_4_3_LC_2_11_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_3_LC_2_11_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_4_3_LC_2_11_5 (
            .in0(N__29976),
            .in1(N__22362),
            .in2(N__30336),
            .in3(N__23658),
            .lcout(TXbuffer_18_13_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIJBVT_15_LC_2_11_6 .C_ON=1'b0;
    defparam \ALU.r5_RNIJBVT_15_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIJBVT_15_LC_2_11_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r5_RNIJBVT_15_LC_2_11_6  (
            .in0(N__30447),
            .in1(N__25078),
            .in2(_gnd_net_),
            .in3(N__29721),
            .lcout(),
            .ltout(\ALU.r5_RNIJBVTZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIJING2_15_LC_2_11_7 .C_ON=1'b0;
    defparam \ALU.r1_RNIJING2_15_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIJING2_15_LC_2_11_7 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.r1_RNIJING2_15_LC_2_11_7  (
            .in0(N__24641),
            .in1(N__20494),
            .in2(N__20488),
            .in3(N__21963),
            .lcout(\ALU.b_7_ns_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_11_s1_c_RNO_LC_2_12_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_11_s1_c_RNO_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_11_s1_c_RNO_LC_2_12_0 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_11_s1_c_RNO_LC_2_12_0  (
            .in0(N__35568),
            .in1(N__53238),
            .in2(N__54780),
            .in3(N__40960),
            .lcout(\ALU.r0_12_prm_5_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIE0AK8_2_11_LC_2_12_3 .C_ON=1'b0;
    defparam \ALU.r5_RNIE0AK8_2_11_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIE0AK8_2_11_LC_2_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r5_RNIE0AK8_2_11_LC_2_12_3  (
            .in0(N__40961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35566),
            .lcout(\ALU.r5_RNIE0AK8_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_9_s0_c_RNO_LC_2_12_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_9_s0_c_RNO_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_9_s0_c_RNO_LC_2_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_9_s0_c_RNO_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__55968),
            .in2(_gnd_net_),
            .in3(N__42448),
            .lcout(\ALU.r0_12_prm_2_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIUF9K8_2_10_LC_2_12_5 .C_ON=1'b0;
    defparam \ALU.r5_RNIUF9K8_2_10_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIUF9K8_2_10_LC_2_12_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \ALU.r5_RNIUF9K8_2_10_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__51983),
            .in2(_gnd_net_),
            .in3(N__51836),
            .lcout(\ALU.r5_RNIUF9K8_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_11_s1_c_RNO_LC_2_12_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_11_s1_c_RNO_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_11_s1_c_RNO_LC_2_12_6 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \ALU.r0_12_prm_7_11_s1_c_RNO_LC_2_12_6  (
            .in0(N__35567),
            .in1(N__53237),
            .in2(_gnd_net_),
            .in3(N__40959),
            .lcout(\ALU.r0_12_prm_7_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIAG9A9_15_LC_2_12_7 .C_ON=1'b0;
    defparam \ALU.r5_RNIAG9A9_15_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIAG9A9_15_LC_2_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r5_RNIAG9A9_15_LC_2_12_7  (
            .in0(N__53680),
            .in1(N__40054),
            .in2(_gnd_net_),
            .in3(N__47046),
            .lcout(\ALU.r5_RNIAG9A9Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIE0AK8_0_11_LC_2_13_0 .C_ON=1'b0;
    defparam \ALU.r5_RNIE0AK8_0_11_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIE0AK8_0_11_LC_2_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.r5_RNIE0AK8_0_11_LC_2_13_0  (
            .in0(N__35569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40958),
            .lcout(\ALU.r5_RNIE0AK8_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_15_s1_c_RNO_LC_2_13_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_15_s1_c_RNO_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_15_s1_c_RNO_LC_2_13_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r0_12_prm_4_15_s1_c_RNO_LC_2_13_2  (
            .in0(N__40086),
            .in1(N__53256),
            .in2(N__54778),
            .in3(N__53685),
            .lcout(\ALU.r0_12_prm_4_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_15_s1_c_RNO_LC_2_13_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_15_s1_c_RNO_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_15_s1_c_RNO_LC_2_13_3 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_15_s1_c_RNO_LC_2_13_3  (
            .in0(N__39957),
            .in1(N__53255),
            .in2(N__53899),
            .in3(N__40085),
            .lcout(\ALU.r0_12_prm_6_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI39IH4_15_LC_2_13_4 .C_ON=1'b0;
    defparam \ALU.r5_RNI39IH4_15_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI39IH4_15_LC_2_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.r5_RNI39IH4_15_LC_2_13_4  (
            .in0(N__25492),
            .in1(N__36764),
            .in2(_gnd_net_),
            .in3(N__21412),
            .lcout(\ALU.a_15 ),
            .ltout(\ALU.a_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNINNEH9_15_LC_2_13_5 .C_ON=1'b0;
    defparam \ALU.r5_RNINNEH9_15_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNINNEH9_15_LC_2_13_5 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.r5_RNINNEH9_15_LC_2_13_5  (
            .in0(N__53681),
            .in1(N__47033),
            .in2(N__20512),
            .in3(N__54585),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIVF7TI_13_LC_2_13_6 .C_ON=1'b0;
    defparam \ALU.r5_RNIVF7TI_13_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIVF7TI_13_LC_2_13_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r5_RNIVF7TI_13_LC_2_13_6  (
            .in0(N__54586),
            .in1(N__41520),
            .in2(N__20509),
            .in3(N__41317),
            .lcout(\ALU.r5_RNIVF7TIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_11_s1_c_RNO_LC_2_13_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_11_s1_c_RNO_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_11_s1_c_RNO_LC_2_13_7 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \ALU.r0_12_prm_1_11_s1_c_RNO_LC_2_13_7  (
            .in0(N__53686),
            .in1(N__55969),
            .in2(_gnd_net_),
            .in3(N__35768),
            .lcout(\ALU.r0_12_prm_1_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_13_LC_2_14_0 .C_ON=1'b0;
    defparam \ALU.r2_13_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_13_LC_2_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_13_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26281),
            .lcout(r2_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56301),
            .ce(N__47707),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINFOB1_13_LC_2_14_1 .C_ON=1'b0;
    defparam \ALU.r2_RNINFOB1_13_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINFOB1_13_LC_2_14_1 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r2_RNINFOB1_13_LC_2_14_1  (
            .in0(N__25066),
            .in1(N__24106),
            .in2(N__22000),
            .in3(N__23906),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIC9GA2_13_LC_2_14_2 .C_ON=1'b0;
    defparam \ALU.r6_RNIC9GA2_13_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIC9GA2_13_LC_2_14_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIC9GA2_13_LC_2_14_2  (
            .in0(N__23988),
            .in1(N__24078),
            .in2(N__20506),
            .in3(N__21999),
            .lcout(),
            .ltout(\ALU.r6_RNIC9GA2Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIR9125_13_LC_2_14_3 .C_ON=1'b0;
    defparam \ALU.r5_RNIR9125_13_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIR9125_13_LC_2_14_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.r5_RNIR9125_13_LC_2_14_3  (
            .in0(N__21421),
            .in1(_gnd_net_),
            .in2(N__20545),
            .in3(N__32896),
            .lcout(\ALU.b_13 ),
            .ltout(\ALU.b_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNID2JJ9_2_13_LC_2_14_4 .C_ON=1'b0;
    defparam \ALU.r5_RNID2JJ9_2_13_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNID2JJ9_2_13_LC_2_14_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \ALU.r5_RNID2JJ9_2_13_LC_2_14_4  (
            .in0(N__41544),
            .in1(_gnd_net_),
            .in2(N__20542),
            .in3(_gnd_net_),
            .lcout(\ALU.r5_RNID2JJ9_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNID2JJ9_0_13_LC_2_14_5 .C_ON=1'b0;
    defparam \ALU.r5_RNID2JJ9_0_13_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNID2JJ9_0_13_LC_2_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.r5_RNID2JJ9_0_13_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__35347),
            .in2(_gnd_net_),
            .in3(N__41542),
            .lcout(\ALU.r5_RNID2JJ9_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNID2JJ9_1_13_LC_2_14_7 .C_ON=1'b0;
    defparam \ALU.r5_RNID2JJ9_1_13_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNID2JJ9_1_13_LC_2_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r5_RNID2JJ9_1_13_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__35348),
            .in2(_gnd_net_),
            .in3(N__41543),
            .lcout(\ALU.r5_RNID2JJ9_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_4_LC_2_15_2.C_ON=1'b0;
    defparam TXbuffer_RNO_4_4_LC_2_15_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_4_LC_2_15_2.LUT_INIT=16'b0001000110101111;
    LogicCell40 TXbuffer_RNO_4_4_LC_2_15_2 (
            .in0(N__29934),
            .in1(N__23872),
            .in2(N__24958),
            .in3(N__30208),
            .lcout(),
            .ltout(TXbuffer_18_13_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_4_LC_2_15_3.C_ON=1'b0;
    defparam TXbuffer_RNO_1_4_LC_2_15_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_4_LC_2_15_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_1_4_LC_2_15_3 (
            .in0(N__29844),
            .in1(N__23622),
            .in2(N__20539),
            .in3(N__28027),
            .lcout(TXbuffer_RNO_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_6_LC_2_15_7.C_ON=1'b0;
    defparam TXbuffer_RNO_8_6_LC_2_15_7.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_6_LC_2_15_7.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_8_6_LC_2_15_7 (
            .in0(N__29843),
            .in1(N__25861),
            .in2(N__30268),
            .in3(N__23745),
            .lcout(TXbuffer_18_6_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_5_LC_2_17_0.C_ON=1'b0;
    defparam TXbuffer_RNO_7_5_LC_2_17_0.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_5_LC_2_17_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_7_5_LC_2_17_0 (
            .in0(N__29903),
            .in1(N__26212),
            .in2(N__30360),
            .in3(N__22333),
            .lcout(TXbuffer_18_3_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_4_LC_3_1_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_4_LC_3_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_4_LC_3_1_0 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_g0_4_LC_3_1_0  (
            .in0(N__46204),
            .in1(N__20704),
            .in2(N__20722),
            .in3(N__37964),
            .lcout(\ALU.N_661_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_155_LC_3_1_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_155_LC_3_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_155_LC_3_1_1 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \ALU.mult_madd_155_LC_3_1_1  (
            .in0(N__21607),
            .in1(N__48576),
            .in2(N__46431),
            .in3(N__20665),
            .lcout(\ALU.madd_155 ),
            .ltout(\ALU.madd_155_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_160_LC_3_1_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_160_LC_3_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_160_LC_3_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_160_LC_3_1_2  (
            .in0(_gnd_net_),
            .in1(N__20568),
            .in2(N__20611),
            .in3(N__22814),
            .lcout(\ALU.madd_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_109_0_tz_LC_3_1_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_109_0_tz_LC_3_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_109_0_tz_LC_3_1_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_madd_109_0_tz_LC_3_1_3  (
            .in0(N__44750),
            .in1(N__46383),
            .in2(N__48987),
            .in3(N__48575),
            .lcout(),
            .ltout(\ALU.madd_109_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_109_LC_3_1_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_109_LC_3_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_109_LC_3_1_4 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \ALU.mult_madd_109_LC_3_1_4  (
            .in0(N__43570),
            .in1(N__48351),
            .in2(N__20608),
            .in3(N__21625),
            .lcout(\ALU.madd_109 ),
            .ltout(\ALU.madd_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_5_LC_3_1_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_5_LC_3_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_5_LC_3_1_5 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \ALU.mult_g0_5_LC_3_1_5  (
            .in0(N__22816),
            .in1(N__21850),
            .in2(N__20605),
            .in3(N__20557),
            .lcout(\ALU.N_687_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_159_LC_3_1_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_159_LC_3_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_159_LC_3_1_6 .LUT_INIT=16'b1000001011101011;
    LogicCell40 \ALU.mult_madd_159_LC_3_1_6  (
            .in0(N__20664),
            .in1(N__20596),
            .in2(N__21619),
            .in3(N__21631),
            .lcout(\ALU.madd_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_164_LC_3_1_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_164_LC_3_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_164_LC_3_1_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_164_LC_3_1_7  (
            .in0(N__22815),
            .in1(_gnd_net_),
            .in2(N__20572),
            .in3(N__20556),
            .lcout(\ALU.madd_333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a4_b_5_LC_3_2_0 .C_ON=1'b0;
    defparam \ALU.mult_a4_b_5_LC_3_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a4_b_5_LC_3_2_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a4_b_5_LC_3_2_0  (
            .in0(N__32470),
            .in1(N__32376),
            .in2(N__29226),
            .in3(N__45180),
            .lcout(\ALU.a4_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a7_b_1_LC_3_2_1 .C_ON=1'b0;
    defparam \ALU.mult_a7_b_1_LC_3_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a7_b_1_LC_3_2_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a7_b_1_LC_3_2_1  (
            .in0(_gnd_net_),
            .in1(N__44549),
            .in2(_gnd_net_),
            .in3(N__46750),
            .lcout(\ALU.a7_b_1 ),
            .ltout(\ALU.a7_b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_95_LC_3_2_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_95_LC_3_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_95_LC_3_2_2 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_95_LC_3_2_2  (
            .in0(N__46153),
            .in1(N__20718),
            .in2(N__20548),
            .in3(N__37966),
            .lcout(\ALU.madd_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a6_b_2_LC_3_2_3 .C_ON=1'b0;
    defparam \ALU.mult_a6_b_2_LC_3_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a6_b_2_LC_3_2_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a6_b_2_LC_3_2_3  (
            .in0(N__26512),
            .in1(N__26448),
            .in2(N__29227),
            .in3(N__43928),
            .lcout(\ALU.a6_b_2 ),
            .ltout(\ALU.a6_b_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_99_LC_3_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_99_LC_3_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_99_LC_3_2_4 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_99_LC_3_2_4  (
            .in0(N__46152),
            .in1(N__37965),
            .in2(N__20707),
            .in3(N__20703),
            .lcout(\ALU.madd_99 ),
            .ltout(\ALU.madd_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_149_LC_3_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_149_LC_3_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_149_LC_3_2_5 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_149_LC_3_2_5  (
            .in0(N__48926),
            .in1(N__47413),
            .in2(N__20692),
            .in3(N__22091),
            .lcout(\ALU.madd_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_145_LC_3_2_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_145_LC_3_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_145_LC_3_2_6 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \ALU.mult_madd_145_LC_3_2_6  (
            .in0(N__22092),
            .in1(N__20671),
            .in2(N__47455),
            .in3(N__48927),
            .lcout(\ALU.madd_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_253_LC_3_2_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_253_LC_3_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_253_LC_3_2_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_253_LC_3_2_7  (
            .in0(N__20656),
            .in1(_gnd_net_),
            .in2(N__20650),
            .in3(N__20640),
            .lcout(\ALU.madd_253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_9_LC_3_3_0 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_9_LC_3_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_9_LC_3_3_0 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \ALU.mult_a3_b_9_LC_3_3_0  (
            .in0(N__47436),
            .in1(N__31924),
            .in2(N__31840),
            .in3(N__36759),
            .lcout(\ALU.a3_b_9 ),
            .ltout(\ALU.a3_b_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_274_LC_3_3_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_274_LC_3_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_274_LC_3_3_1 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_274_LC_3_3_1  (
            .in0(N__21093),
            .in1(N__35573),
            .in2(N__20620),
            .in3(N__48568),
            .lcout(\ALU.madd_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_278_LC_3_3_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_278_LC_3_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_278_LC_3_3_2 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \ALU.mult_madd_278_LC_3_3_2  (
            .in0(N__48567),
            .in1(N__20617),
            .in2(N__35593),
            .in3(N__21094),
            .lcout(\ALU.madd_278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_11_l_fx_LC_3_3_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_11_l_fx_LC_3_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_11_l_fx_LC_3_3_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.mult_madd_axb_11_l_fx_LC_3_3_3  (
            .in0(N__20832),
            .in1(N__27480),
            .in2(_gnd_net_),
            .in3(N__20855),
            .lcout(\ALU.madd_axb_11_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_273_LC_3_3_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_273_LC_3_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_273_LC_3_3_4 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_273_LC_3_3_4  (
            .in0(N__43394),
            .in1(N__43639),
            .in2(N__21760),
            .in3(N__20803),
            .lcout(\ALU.madd_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a4_b_8_LC_3_3_5 .C_ON=1'b0;
    defparam \ALU.mult_a4_b_8_LC_3_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a4_b_8_LC_3_3_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a4_b_8_LC_3_3_5  (
            .in0(N__32471),
            .in1(N__32377),
            .in2(N__36778),
            .in3(N__46336),
            .lcout(\ALU.a4_b_8 ),
            .ltout(\ALU.a4_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_269_LC_3_3_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_269_LC_3_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_269_LC_3_3_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ALU.mult_madd_269_LC_3_3_6  (
            .in0(N__43395),
            .in1(N__43638),
            .in2(N__20797),
            .in3(N__21759),
            .lcout(\ALU.madd_269 ),
            .ltout(\ALU.madd_269_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_289_LC_3_3_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_289_LC_3_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_289_LC_3_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_289_LC_3_3_7  (
            .in0(_gnd_net_),
            .in1(N__20787),
            .in2(N__20773),
            .in3(N__20971),
            .lcout(\ALU.madd_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_185_1_LC_3_4_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_185_1_LC_3_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_185_1_LC_3_4_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ALU.mult_madd_185_1_LC_3_4_1  (
            .in0(_gnd_net_),
            .in1(N__37973),
            .in2(_gnd_net_),
            .in3(N__52222),
            .lcout(),
            .ltout(\ALU.madd_185_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_185_LC_3_4_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_185_LC_3_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_185_LC_3_4_2 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \ALU.mult_madd_185_LC_3_4_2  (
            .in0(N__21799),
            .in1(N__23037),
            .in2(N__20752),
            .in3(N__22113),
            .lcout(\ALU.madd_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_2_N_2L1_LC_3_4_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_2_N_2L1_LC_3_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_2_N_2L1_LC_3_4_3 .LUT_INIT=16'b0101001111111111;
    LogicCell40 \ALU.mult_g0_2_N_2L1_LC_3_4_3  (
            .in0(N__21313),
            .in1(N__21292),
            .in2(N__24655),
            .in3(N__48553),
            .lcout(),
            .ltout(\ALU.g0_2_N_2L1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_2_LC_3_4_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_2_LC_3_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_2_LC_3_4_4 .LUT_INIT=16'b0000111100000001;
    LogicCell40 \ALU.mult_g0_2_LC_3_4_4  (
            .in0(N__22129),
            .in1(N__22009),
            .in2(N__20737),
            .in3(N__22135),
            .lcout(\ALU.madd_186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_218_0_tz_LC_3_4_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_218_0_tz_LC_3_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_218_0_tz_LC_3_4_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_218_0_tz_LC_3_4_5  (
            .in0(N__45206),
            .in1(N__40509),
            .in2(N__43425),
            .in3(N__44551),
            .lcout(\ALU.madd_218_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_228_LC_3_4_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_228_LC_3_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_228_LC_3_4_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ALU.mult_madd_228_LC_3_4_6  (
            .in0(N__22963),
            .in1(N__22102),
            .in2(N__47456),
            .in3(N__48307),
            .lcout(\ALU.madd_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_217_LC_3_4_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_217_LC_3_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_217_LC_3_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_217_LC_3_4_7  (
            .in0(N__45205),
            .in1(N__40508),
            .in2(N__43424),
            .in3(N__44550),
            .lcout(\ALU.madd_124_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_13_l_ofx_LC_3_5_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_13_l_ofx_LC_3_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_13_l_ofx_LC_3_5_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.mult_madd_axb_13_l_ofx_LC_3_5_0  (
            .in0(N__20955),
            .in1(N__21163),
            .in2(N__21151),
            .in3(N__20940),
            .lcout(\ALU.madd_axb_13_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_335_LC_3_5_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_335_LC_3_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_335_LC_3_5_1 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \ALU.mult_madd_335_LC_3_5_1  (
            .in0(N__20929),
            .in1(N__21262),
            .in2(N__39850),
            .in3(N__48611),
            .lcout(\ALU.madd_335_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_12_ma_LC_3_5_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_12_ma_LC_3_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_12_ma_LC_3_5_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_cry_12_ma_LC_3_5_2  (
            .in0(_gnd_net_),
            .in1(N__20838),
            .in2(_gnd_net_),
            .in3(N__20856),
            .lcout(\ALU.madd_cry_12_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_294_LC_3_5_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_294_LC_3_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_294_LC_3_5_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_294_LC_3_5_3  (
            .in0(N__20911),
            .in1(N__21008),
            .in2(N__20896),
            .in3(N__21078),
            .lcout(\ALU.madd_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_12_l_ofx_LC_3_5_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_12_l_ofx_LC_3_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_12_l_ofx_LC_3_5_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_axb_12_l_ofx_LC_3_5_4  (
            .in0(N__20857),
            .in1(N__20839),
            .in2(N__21150),
            .in3(N__21161),
            .lcout(\ALU.madd_axb_12_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_5_s0_c_RNO_LC_3_5_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_5_s0_c_RNO_LC_3_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_5_s0_c_RNO_LC_3_5_5 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \ALU.r0_12_prm_7_5_s0_c_RNO_LC_3_5_5  (
            .in0(N__47255),
            .in1(N__53145),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_7_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_341_LC_3_5_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_341_LC_3_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_341_LC_3_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_341_LC_3_5_6  (
            .in0(N__21708),
            .in1(N__22032),
            .in2(_gnd_net_),
            .in3(N__21691),
            .lcout(\ALU.madd_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_13_ma_LC_3_5_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_13_ma_LC_3_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_13_ma_LC_3_5_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_madd_cry_13_ma_LC_3_5_7  (
            .in0(N__21162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21143),
            .lcout(\ALU.madd_cry_13_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_283_LC_3_6_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_283_LC_3_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_283_LC_3_6_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_283_LC_3_6_0  (
            .in0(N__22226),
            .in1(N__21029),
            .in2(_gnd_net_),
            .in3(N__21001),
            .lcout(\ALU.madd_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_218_LC_3_6_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_218_LC_3_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_218_LC_3_6_1 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \ALU.mult_madd_218_LC_3_6_1  (
            .in0(N__21124),
            .in1(N__46103),
            .in2(N__21115),
            .in3(N__44343),
            .lcout(\ALU.madd_218 ),
            .ltout(\ALU.madd_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_346_1_LC_3_6_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_346_1_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_346_1_LC_3_6_2 .LUT_INIT=16'b0000010101011111;
    LogicCell40 \ALU.mult_madd_346_1_LC_3_6_2  (
            .in0(N__22225),
            .in1(_gnd_net_),
            .in2(N__21103),
            .in3(N__21028),
            .lcout(\ALU.madd_346_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_10_LC_3_6_3 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_10_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_10_LC_3_6_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a2_b_10_LC_3_6_3  (
            .in0(N__51908),
            .in1(N__32666),
            .in2(N__36755),
            .in3(N__32570),
            .lcout(\ALU.a2_b_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_12_LC_3_6_4 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_12_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_12_LC_3_6_4 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \ALU.mult_a0_b_12_LC_3_6_4  (
            .in0(N__21445),
            .in1(N__21454),
            .in2(N__32894),
            .in3(N__48916),
            .lcout(\ALU.a0_b_12 ),
            .ltout(\ALU.a0_b_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_279_0_LC_3_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_279_0_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_279_0_LC_3_6_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_279_0_LC_3_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21082),
            .in3(N__22224),
            .lcout(\ALU.madd_279_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_349_LC_3_6_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_349_LC_3_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_349_LC_3_6_6 .LUT_INIT=16'b1100100010000000;
    LogicCell40 \ALU.mult_madd_349_LC_3_6_6  (
            .in0(N__22227),
            .in1(N__21063),
            .in2(N__21036),
            .in3(N__21002),
            .lcout(\ALU.madd_202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a7_b_5_LC_3_6_7 .C_ON=1'b0;
    defparam \ALU.mult_a7_b_5_LC_3_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a7_b_5_LC_3_6_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a7_b_5_LC_3_6_7  (
            .in0(N__45106),
            .in1(N__23106),
            .in2(N__36754),
            .in3(N__30724),
            .lcout(\ALU.a7_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a12_b_0_LC_3_7_0 .C_ON=1'b0;
    defparam \ALU.mult_a12_b_0_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a12_b_0_LC_3_7_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a12_b_0_LC_3_7_0  (
            .in0(N__41276),
            .in1(N__32748),
            .in2(N__32864),
            .in3(N__32719),
            .lcout(\ALU.a12_b_0 ),
            .ltout(\ALU.a12_b_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_263_LC_3_7_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_263_LC_3_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_263_LC_3_7_1 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_263_LC_3_7_1  (
            .in0(N__21228),
            .in1(N__40876),
            .in2(N__21265),
            .in3(N__46780),
            .lcout(\ALU.madd_263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a10_b_2_LC_3_7_2 .C_ON=1'b0;
    defparam \ALU.mult_a10_b_2_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a10_b_2_LC_3_7_2 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.mult_a10_b_2_LC_3_7_2  (
            .in0(N__29364),
            .in1(N__51747),
            .in2(N__32863),
            .in3(N__33348),
            .lcout(\ALU.a10_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_264_LC_3_7_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_264_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_264_LC_3_7_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_264_LC_3_7_3  (
            .in0(N__22205),
            .in1(_gnd_net_),
            .in2(N__21211),
            .in3(N__23262),
            .lcout(),
            .ltout(\ALU.madd_264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_288_LC_3_7_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_288_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_288_LC_3_7_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_288_LC_3_7_4  (
            .in0(_gnd_net_),
            .in1(N__21217),
            .in2(N__21247),
            .in3(N__22872),
            .lcout(\ALU.madd_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_259_LC_3_7_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_259_LC_3_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_259_LC_3_7_5 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_259_LC_3_7_5  (
            .in0(N__21235),
            .in1(N__40877),
            .in2(N__21229),
            .in3(N__46781),
            .lcout(\ALU.madd_259 ),
            .ltout(\ALU.madd_259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_284_0_LC_3_7_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_284_0_LC_3_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_284_0_LC_3_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_284_0_LC_3_7_6  (
            .in0(N__23263),
            .in1(N__21206),
            .in2(N__21190),
            .in3(N__22206),
            .lcout(\ALU.madd_284_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIUOP24_10_LC_3_7_7 .C_ON=1'b0;
    defparam \ALU.r5_RNIUOP24_10_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIUOP24_10_LC_3_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r5_RNIUOP24_10_LC_3_7_7  (
            .in0(N__24654),
            .in1(N__21834),
            .in2(_gnd_net_),
            .in3(N__21810),
            .lcout(\ALU.b_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIRP8Q_9_LC_3_8_0 .C_ON=1'b0;
    defparam \ALU.r0_RNIRP8Q_9_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIRP8Q_9_LC_3_8_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r0_RNIRP8Q_9_LC_3_8_0  (
            .in0(N__29486),
            .in1(N__31011),
            .in2(N__26858),
            .in3(N__31146),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIM58R1_9_LC_3_8_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIM58R1_9_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIM58R1_9_LC_3_8_1 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.r4_RNIM58R1_9_LC_3_8_1  (
            .in0(N__33687),
            .in1(N__21968),
            .in2(N__21295),
            .in3(N__34405),
            .lcout(\ALU.r4_RNIM58R1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_0_rep2_LC_3_8_2.C_ON=1'b0;
    defparam b_0_rep2_LC_3_8_2.SEQ_MODE=4'b1000;
    defparam b_0_rep2_LC_3_8_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 b_0_rep2_LC_3_8_2 (
            .in0(N__29489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_0_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56270),
            .ce(N__56043),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIB9GU_10_LC_3_8_3 .C_ON=1'b0;
    defparam \ALU.r1_RNIB9GU_10_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIB9GU_10_LC_3_8_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r1_RNIB9GU_10_LC_3_8_3  (
            .in0(N__28123),
            .in1(N__26844),
            .in2(N__27973),
            .in3(N__29487),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIMCFS1_10_LC_3_8_4 .C_ON=1'b0;
    defparam \ALU.r5_RNIMCFS1_10_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIMCFS1_10_LC_3_8_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r5_RNIMCFS1_10_LC_3_8_4  (
            .in0(N__21969),
            .in1(N__27937),
            .in2(N__21277),
            .in3(N__25483),
            .lcout(\ALU.r5_RNIMCFS1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIDBGU_11_LC_3_8_5 .C_ON=1'b0;
    defparam \ALU.r1_RNIDBGU_11_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIDBGU_11_LC_3_8_5 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r1_RNIDBGU_11_LC_3_8_5  (
            .in0(N__24539),
            .in1(N__29488),
            .in2(N__25216),
            .in3(N__26845),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIQGFS1_11_LC_3_8_6 .C_ON=1'b0;
    defparam \ALU.r5_RNIQGFS1_11_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIQGFS1_11_LC_3_8_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r5_RNIQGFS1_11_LC_3_8_6  (
            .in0(N__21970),
            .in1(N__26119),
            .in2(N__21274),
            .in3(N__24736),
            .lcout(),
            .ltout(\ALU.r5_RNIQGFS1Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI61Q24_11_LC_3_8_7 .C_ON=1'b0;
    defparam \ALU.r5_RNI61Q24_11_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI61Q24_11_LC_3_8_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.r5_RNI61Q24_11_LC_3_8_7  (
            .in0(_gnd_net_),
            .in1(N__24631),
            .in2(N__21271),
            .in3(N__21325),
            .lcout(\ALU.b_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIFP8V_10_LC_3_9_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIFP8V_10_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIFP8V_10_LC_3_9_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \ALU.r2_RNIFP8V_10_LC_3_9_0  (
            .in0(N__22290),
            .in1(N__26856),
            .in2(N__29516),
            .in3(N__22385),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIUC0U1_10_LC_3_9_1 .C_ON=1'b0;
    defparam \ALU.r6_RNIUC0U1_10_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIUC0U1_10_LC_3_9_1 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.r6_RNIUC0U1_10_LC_3_9_1  (
            .in0(N__22680),
            .in1(N__21943),
            .in2(N__21268),
            .in3(N__22573),
            .lcout(\ALU.r6_RNIUC0U1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_10_LC_3_9_2 .C_ON=1'b0;
    defparam \ALU.r2_10_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_10_LC_3_9_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ALU.r2_10_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__28192),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r2_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56275),
            .ce(N__47716),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIHR8V_11_LC_3_9_3 .C_ON=1'b0;
    defparam \ALU.r2_RNIHR8V_11_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIHR8V_11_LC_3_9_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r2_RNIHR8V_11_LC_3_9_3  (
            .in0(N__29481),
            .in1(N__22361),
            .in2(N__26860),
            .in3(N__24816),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI2H0U1_11_LC_3_9_4 .C_ON=1'b0;
    defparam \ALU.r6_RNI2H0U1_11_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI2H0U1_11_LC_3_9_4 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.r6_RNI2H0U1_11_LC_3_9_4  (
            .in0(N__24768),
            .in1(N__21934),
            .in2(N__21328),
            .in3(N__22649),
            .lcout(\ALU.r6_RNI2H0U1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_11_LC_3_9_5 .C_ON=1'b0;
    defparam \ALU.r2_11_LC_3_9_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_11_LC_3_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_11_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26172),
            .lcout(r2_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56275),
            .ce(N__47716),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIV5LU_9_LC_3_9_6 .C_ON=1'b0;
    defparam \ALU.r2_RNIV5LU_9_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIV5LU_9_LC_3_9_6 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \ALU.r2_RNIV5LU_9_LC_3_9_6  (
            .in0(N__27581),
            .in1(N__29482),
            .in2(N__23710),
            .in3(N__26857),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIUT042_9_LC_3_9_7 .C_ON=1'b0;
    defparam \ALU.r6_RNIUT042_9_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIUT042_9_LC_3_9_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNIUT042_9_LC_3_9_7  (
            .in0(N__21935),
            .in1(N__27795),
            .in2(N__21316),
            .in3(N__22255),
            .lcout(\ALU.r6_RNIUT042Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIDP6T_14_LC_3_10_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIDP6T_14_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIDP6T_14_LC_3_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r2_RNIDP6T_14_LC_3_10_0  (
            .in0(N__25830),
            .in1(N__25857),
            .in2(_gnd_net_),
            .in3(N__25076),
            .lcout(\ALU.r2_RNIDP6TZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNILPNU_14_LC_3_10_1 .C_ON=1'b0;
    defparam \ALU.r6_RNILPNU_14_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNILPNU_14_LC_3_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r6_RNILPNU_14_LC_3_10_1  (
            .in0(N__25075),
            .in1(N__25798),
            .in2(_gnd_net_),
            .in3(N__25763),
            .lcout(\ALU.r6_RNILPNUZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIH9VT_14_LC_3_10_2 .C_ON=1'b0;
    defparam \ALU.r5_RNIH9VT_14_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIH9VT_14_LC_3_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r5_RNIH9VT_14_LC_3_10_2  (
            .in0(N__26026),
            .in1(N__25887),
            .in2(_gnd_net_),
            .in3(N__25074),
            .lcout(\ALU.r5_RNIH9VTZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNI8DSR_14_LC_3_10_3 .C_ON=1'b0;
    defparam \ALU.r1_RNI8DSR_14_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNI8DSR_14_LC_3_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.r1_RNI8DSR_14_LC_3_10_3  (
            .in0(N__25719),
            .in1(N__28245),
            .in2(_gnd_net_),
            .in3(N__29508),
            .lcout(),
            .ltout(\ALU.r1_RNI8DSRZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIFENG2_14_LC_3_10_4 .C_ON=1'b0;
    defparam \ALU.r1_RNIFENG2_14_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIFENG2_14_LC_3_10_4 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \ALU.r1_RNIFENG2_14_LC_3_10_4  (
            .in0(N__24649),
            .in1(N__21379),
            .in2(N__21373),
            .in3(N__21964),
            .lcout(),
            .ltout(\ALU.b_7_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNISO7R4_14_LC_3_10_5 .C_ON=1'b0;
    defparam \ALU.r2_RNISO7R4_14_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNISO7R4_14_LC_3_10_5 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r2_RNISO7R4_14_LC_3_10_5  (
            .in0(N__32887),
            .in1(N__21370),
            .in2(N__21364),
            .in3(N__21361),
            .lcout(\ALU.b_14 ),
            .ltout(\ALU.b_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINPPC9_2_14_LC_3_10_6 .C_ON=1'b0;
    defparam \ALU.r2_RNINPPC9_2_14_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINPPC9_2_14_LC_3_10_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \ALU.r2_RNINPPC9_2_14_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21355),
            .in3(N__47045),
            .lcout(\ALU.r2_RNINPPC9_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_2_LC_3_10_7.C_ON=1'b0;
    defparam b_2_LC_3_10_7.SEQ_MODE=4'b1000;
    defparam b_2_LC_3_10_7.LUT_INIT=16'b0101101011110000;
    LogicCell40 b_2_LC_3_10_7 (
            .in0(N__25077),
            .in1(_gnd_net_),
            .in2(N__21991),
            .in3(N__32893),
            .lcout(bZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56280),
            .ce(N__56041),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_0_LC_3_11_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_0_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_0_LC_3_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_11_s1_c_RNO_0_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__34234),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\ALU.r0_12_prm_8_11_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s1_c_LC_3_11_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_11_s1_c_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s1_c_LC_3_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_11_s1_c_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__34444),
            .in2(N__31120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_11_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_11_s1_c_LC_3_11_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_11_s1_c_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_11_s1_c_LC_3_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_11_s1_c_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__21498),
            .in2(N__21352),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_11_s1 ),
            .carryout(\ALU.r0_12_prm_7_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_11_s1_c_LC_3_11_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_11_s1_c_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_11_s1_c_LC_3_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_11_s1_c_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__35145),
            .in2(N__22783),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_11_s1 ),
            .carryout(\ALU.r0_12_prm_6_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_11_s1_c_LC_3_11_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_11_s1_c_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_11_s1_c_LC_3_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_11_s1_c_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__21471),
            .in2(N__21340),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_11_s1 ),
            .carryout(\ALU.r0_12_prm_5_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_11_s1_c_LC_3_11_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_11_s1_c_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_11_s1_c_LC_3_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_11_s1_c_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(N__21601),
            .in2(N__22711),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_11_s1 ),
            .carryout(\ALU.r0_12_prm_4_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_11_s1_c_LC_3_11_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_11_s1_c_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_11_s1_c_LC_3_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_11_s1_c_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(N__56398),
            .in2(N__55259),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_11_s1 ),
            .carryout(\ALU.r0_12_prm_3_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_11_s1_c_LC_3_11_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_11_s1_c_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_11_s1_c_LC_3_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_11_s1_c_LC_3_11_7  (
            .in0(_gnd_net_),
            .in1(N__35844),
            .in2(N__35806),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_11_s1 ),
            .carryout(\ALU.r0_12_prm_2_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_11_s1_c_LC_3_12_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_11_s1_c_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_11_s1_c_LC_3_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_11_s1_c_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__35772),
            .in2(N__21394),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\ALU.r0_12_s1_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_11_s0_c_RNI9L4SLH1_LC_3_12_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_11_s0_c_RNI9L4SLH1_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_11_s0_c_RNI9L4SLH1_LC_3_12_1 .LUT_INIT=16'b1011111010000010;
    LogicCell40 \ALU.r0_12_prm_1_11_s0_c_RNI9L4SLH1_LC_3_12_1  (
            .in0(N__21574),
            .in1(N__27534),
            .in2(N__27508),
            .in3(N__21385),
            .lcout(\ALU.r0_12_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_11_LC_3_12_2 .C_ON=1'b0;
    defparam \ALU.r0_11_LC_3_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_11_LC_3_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_11_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26154),
            .lcout(r0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56288),
            .ce(N__49733),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIHTVA1_12_LC_3_13_0 .C_ON=1'b0;
    defparam \ALU.r1_RNIHTVA1_12_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIHTVA1_12_LC_3_13_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r1_RNIHTVA1_12_LC_3_13_0  (
            .in0(N__25047),
            .in1(N__25170),
            .in2(N__21995),
            .in3(N__28373),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI05V82_12_LC_3_13_1 .C_ON=1'b0;
    defparam \ALU.r5_RNI05V82_12_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI05V82_12_LC_3_13_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r5_RNI05V82_12_LC_3_13_1  (
            .in0(N__26079),
            .in1(N__25453),
            .in2(N__21382),
            .in3(N__21984),
            .lcout(\ALU.r5_RNI05V82Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNILDOB1_12_LC_3_13_2 .C_ON=1'b0;
    defparam \ALU.r2_RNILDOB1_12_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNILDOB1_12_LC_3_13_2 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.r2_RNILDOB1_12_LC_3_13_2  (
            .in0(N__21980),
            .in1(N__23871),
            .in2(N__25073),
            .in3(N__25317),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI85GA2_12_LC_3_13_3 .C_ON=1'b0;
    defparam \ALU.r6_RNI85GA2_12_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI85GA2_12_LC_3_13_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNI85GA2_12_LC_3_13_3  (
            .in0(N__23623),
            .in1(N__25257),
            .in2(N__21457),
            .in3(N__21985),
            .lcout(\ALU.r6_RNI85GA2Z0Z_12 ),
            .ltout(\ALU.r6_RNI85GA2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIJ1125_12_LC_3_13_4 .C_ON=1'b0;
    defparam \ALU.r5_RNIJ1125_12_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIJ1125_12_LC_3_13_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.r5_RNIJ1125_12_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__21438),
            .in2(N__21427),
            .in3(N__32891),
            .lcout(\ALU.b_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_0_LC_3_13_5.C_ON=1'b0;
    defparam b_0_LC_3_13_5.SEQ_MODE=4'b1000;
    defparam b_0_LC_3_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 b_0_LC_3_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25051),
            .lcout(bZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56292),
            .ce(N__56040),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIJVVA1_13_LC_3_13_6 .C_ON=1'b0;
    defparam \ALU.r1_RNIJVVA1_13_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIJVVA1_13_LC_3_13_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r1_RNIJVVA1_13_LC_3_13_6  (
            .in0(N__25046),
            .in1(N__25136),
            .in2(N__21994),
            .in3(N__26211),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI49V82_13_LC_3_13_7 .C_ON=1'b0;
    defparam \ALU.r5_RNI49V82_13_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI49V82_13_LC_3_13_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r5_RNI49V82_13_LC_3_13_7  (
            .in0(N__26050),
            .in1(N__25419),
            .in2(N__21424),
            .in3(N__21979),
            .lcout(\ALU.r5_RNI49V82Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIPDI91_15_LC_3_14_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIPDI91_15_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIPDI91_15_LC_3_14_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIPDI91_15_LC_3_14_0  (
            .in0(N__22424),
            .in1(N__25600),
            .in2(N__22513),
            .in3(N__25679),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIH8772_15_LC_3_14_1 .C_ON=1'b0;
    defparam \ALU.r6_RNIH8772_15_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIH8772_15_LC_3_14_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNIH8772_15_LC_3_14_1  (
            .in0(N__25601),
            .in1(N__22619),
            .in2(N__21415),
            .in3(N__22529),
            .lcout(\ALU.r6_RNIH8772Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_15_LC_3_14_2 .C_ON=1'b0;
    defparam \ALU.r2_15_LC_3_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_15_LC_3_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_15_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25987),
            .lcout(r2_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56297),
            .ce(N__47706),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNINRNU_15_LC_3_14_3 .C_ON=1'b0;
    defparam \ALU.r6_RNINRNU_15_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNINRNU_15_LC_3_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r6_RNINRNU_15_LC_3_14_3  (
            .in0(N__22620),
            .in1(N__22530),
            .in2(_gnd_net_),
            .in3(N__25067),
            .lcout(\ALU.r6_RNINRNUZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIA0841_0_LC_3_14_4 .C_ON=1'b0;
    defparam \ALU.r6_RNIA0841_0_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIA0841_0_LC_3_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r6_RNIA0841_0_LC_3_14_4  (
            .in0(N__23318),
            .in1(N__23282),
            .in2(_gnd_net_),
            .in3(N__25678),
            .lcout(\ALU.r6_RNIA0841Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_0_LC_3_14_5.C_ON=1'b0;
    defparam TXbuffer_RNO_8_0_LC_3_14_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_0_LC_3_14_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_8_0_LC_3_14_5 (
            .in0(N__29985),
            .in1(N__23578),
            .in2(N__30364),
            .in3(N__28741),
            .lcout(),
            .ltout(TXbuffer_18_6_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_0_LC_3_14_6.C_ON=1'b0;
    defparam TXbuffer_RNO_6_0_LC_3_14_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_0_LC_3_14_6.LUT_INIT=16'b1100101100001011;
    LogicCell40 TXbuffer_RNO_6_0_LC_3_14_6 (
            .in0(N__39205),
            .in1(N__29986),
            .in2(N__21526),
            .in3(N__23283),
            .lcout(TXbuffer_RNO_6Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_7_LC_3_14_7.C_ON=1'b0;
    defparam TXbuffer_RNO_1_7_LC_3_14_7.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_7_LC_3_14_7.LUT_INIT=16'b1110001100100011;
    LogicCell40 TXbuffer_RNO_1_7_LC_3_14_7 (
            .in0(N__22621),
            .in1(N__21511),
            .in2(N__30048),
            .in3(N__27850),
            .lcout(TXbuffer_RNO_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_0_LC_3_15_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_0_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_0_LC_3_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_11_s0_c_RNO_0_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__34549),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\ALU.r0_12_prm_8_11_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s0_c_LC_3_15_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_11_s0_c_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s0_c_LC_3_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_11_s0_c_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__34443),
            .in2(N__31303),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_11_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_11_s0_c_LC_3_15_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_11_s0_c_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_11_s0_c_LC_3_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_11_s0_c_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__21499),
            .in2(N__22792),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_11_s0 ),
            .carryout(\ALU.r0_12_prm_7_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_11_s0_c_LC_3_15_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_11_s0_c_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_11_s0_c_LC_3_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_11_s0_c_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__22798),
            .in2(N__35149),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_11_s0 ),
            .carryout(\ALU.r0_12_prm_6_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_11_s0_c_LC_3_15_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_11_s0_c_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_11_s0_c_LC_3_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_11_s0_c_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__22690),
            .in2(N__21478),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_11_s0 ),
            .carryout(\ALU.r0_12_prm_5_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_11_s0_c_inv_LC_3_15_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_11_s0_c_inv_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_11_s0_c_inv_LC_3_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_4_11_s0_c_inv_LC_3_15_5  (
            .in0(N__40969),
            .in1(N__22696),
            .in2(N__21600),
            .in3(_gnd_net_),
            .lcout(\ALU.a_i_11 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_11_s0 ),
            .carryout(\ALU.r0_12_prm_4_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_11_s0_c_inv_LC_3_15_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_11_s0_c_inv_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_11_s0_c_inv_LC_3_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_11_s0_c_inv_LC_3_15_6  (
            .in0(N__55279),
            .in1(N__21583),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_11_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_11_s0 ),
            .carryout(\ALU.r0_12_prm_3_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_11_s0_c_LC_3_15_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_11_s0_c_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_11_s0_c_LC_3_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_11_s0_c_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__34216),
            .in2(N__35845),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_11_s0 ),
            .carryout(\ALU.r0_12_prm_2_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_11_s0_c_LC_3_16_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_11_s0_c_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_11_s0_c_LC_3_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_11_s0_c_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__35773),
            .in2(N__35731),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\ALU.r0_12_s0_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s0_11_THRU_LUT4_0_LC_3_16_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s0_11_THRU_LUT4_0_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s0_11_THRU_LUT4_0_LC_3_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s0_11_THRU_LUT4_0_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21577),
            .lcout(\ALU.r0_12_s0_11_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_21_LC_4_1_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_21_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_21_LC_4_1_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_g0_21_LC_4_1_0  (
            .in0(N__45188),
            .in1(N__32476),
            .in2(N__36784),
            .in3(N__32375),
            .lcout(\ALU.a4_b_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g1_7_LC_4_1_1 .C_ON=1'b0;
    defparam \ALU.mult_g1_7_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g1_7_LC_4_1_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.mult_g1_7_LC_4_1_1  (
            .in0(N__29220),
            .in1(N__29100),
            .in2(_gnd_net_),
            .in3(N__28978),
            .lcout(),
            .ltout(\ALU.g1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_19_LC_4_1_2 .C_ON=1'b0;
    defparam \ALU.mult_g0_19_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_19_LC_4_1_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \ALU.mult_g0_19_LC_4_1_2  (
            .in0(N__22954),
            .in1(N__44347),
            .in2(N__21562),
            .in3(N__24430),
            .lcout(),
            .ltout(\ALU.N_663_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_16_LC_4_1_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_16_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_16_LC_4_1_3 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_g0_16_LC_4_1_3  (
            .in0(N__24175),
            .in1(N__21559),
            .in2(N__21553),
            .in3(N__21548),
            .lcout(\ALU.N_683_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_76_LC_4_1_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_76_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_76_LC_4_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_76_LC_4_1_4  (
            .in0(N__48291),
            .in1(N__40519),
            .in2(N__45230),
            .in3(N__49348),
            .lcout(),
            .ltout(\ALU.madd_43_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_77_LC_4_1_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_77_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_77_LC_4_1_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_madd_77_LC_4_1_5  (
            .in0(N__44348),
            .in1(N__21715),
            .in2(N__21718),
            .in3(N__42815),
            .lcout(\ALU.madd_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_77_0_tz_LC_4_1_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_77_0_tz_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_77_0_tz_LC_4_1_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_77_0_tz_LC_4_1_6  (
            .in0(N__48290),
            .in1(N__40518),
            .in2(N__45229),
            .in3(N__49349),
            .lcout(\ALU.madd_77_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a6_b_7_LC_4_2_0 .C_ON=1'b0;
    defparam \ALU.mult_a6_b_7_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a6_b_7_LC_4_2_0 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \ALU.mult_a6_b_7_LC_4_2_0  (
            .in0(N__44704),
            .in1(N__36625),
            .in2(N__26515),
            .in3(N__26437),
            .lcout(\ALU.a6_b_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_345_LC_4_2_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_345_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_345_LC_4_2_1 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_345_LC_4_2_1  (
            .in0(N__21709),
            .in1(N__22033),
            .in2(_gnd_net_),
            .in3(N__21687),
            .lcout(\ALU.madd_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_159_N_3L3_LC_4_2_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_159_N_3L3_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_159_N_3L3_LC_4_2_2 .LUT_INIT=16'b0000010101011111;
    LogicCell40 \ALU.mult_madd_159_N_3L3_LC_4_2_2  (
            .in0(N__22905),
            .in1(_gnd_net_),
            .in2(N__22939),
            .in3(N__22923),
            .lcout(\ALU.madd_159_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_108_LC_4_2_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_108_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_108_LC_4_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_108_LC_4_2_3  (
            .in0(N__48922),
            .in1(N__46307),
            .in2(N__44763),
            .in3(N__48512),
            .lcout(\ALU.madd_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_140_0_LC_4_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_140_0_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_140_0_LC_4_2_4 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_140_0_LC_4_2_4  (
            .in0(N__44705),
            .in1(N__48289),
            .in2(N__43643),
            .in3(N__49366),
            .lcout(\ALU.madd_140_0 ),
            .ltout(\ALU.madd_140_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_155_1_LC_4_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_155_1_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_155_1_LC_4_2_5 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \ALU.mult_madd_155_1_LC_4_2_5  (
            .in0(N__22922),
            .in1(N__22935),
            .in2(N__21610),
            .in3(N__22904),
            .lcout(\ALU.madd_155_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_144_0_tz_LC_4_2_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_144_0_tz_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_144_0_tz_LC_4_2_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_144_0_tz_LC_4_2_6  (
            .in0(N__48511),
            .in1(N__44719),
            .in2(N__46348),
            .in3(N__48288),
            .lcout(\ALU.madd_144_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_6_1_LC_4_2_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_6_1_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_6_1_LC_4_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_g0_6_1_LC_4_2_7  (
            .in0(N__22843),
            .in1(N__21873),
            .in2(_gnd_net_),
            .in3(N__31563),
            .lcout(\ALU.g0_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_10_LC_4_3_0 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_10_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_10_LC_4_3_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a0_b_10_LC_4_3_0  (
            .in0(N__21838),
            .in1(N__21817),
            .in2(N__24653),
            .in3(N__48830),
            .lcout(\ALU.a0_b_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_8_LC_4_3_1 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_8_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_8_LC_4_3_1 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \ALU.mult_a5_b_8_LC_4_3_1  (
            .in0(N__28999),
            .in1(N__29096),
            .in2(N__36681),
            .in3(N__46308),
            .lcout(\ALU.a5_b_8 ),
            .ltout(\ALU.a5_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_325_LC_4_3_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_325_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_325_LC_4_3_2 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_325_LC_4_3_2  (
            .in0(N__43589),
            .in1(N__22041),
            .in2(N__21793),
            .in3(N__44544),
            .lcout(\ALU.madd_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI435F3_7_LC_4_3_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI435F3_7_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI435F3_7_LC_4_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNI435F3_7_LC_4_3_3  (
            .in0(N__24711),
            .in1(N__22447),
            .in2(_gnd_net_),
            .in3(N__29533),
            .lcout(\ALU.b_7 ),
            .ltout(\ALU.b_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_7_LC_4_3_4 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_7_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_7_LC_4_3_4 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \ALU.mult_a5_b_7_LC_4_3_4  (
            .in0(N__29095),
            .in1(N__36621),
            .in2(N__21763),
            .in3(N__28998),
            .lcout(\ALU.a5_b_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_5_LC_4_3_5 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_5_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_5_LC_4_3_5 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \ALU.mult_a5_b_5_LC_4_3_5  (
            .in0(N__28997),
            .in1(N__29094),
            .in2(N__36680),
            .in3(N__45181),
            .lcout(\ALU.a5_b_5 ),
            .ltout(\ALU.a5_b_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_176_LC_4_3_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_176_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_176_LC_4_3_6 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_176_LC_4_3_6  (
            .in0(N__43280),
            .in1(N__22972),
            .in2(N__21745),
            .in3(N__40510),
            .lcout(\ALU.madd_176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_321_LC_4_3_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_321_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_321_LC_4_3_7 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_321_LC_4_3_7  (
            .in0(N__44545),
            .in1(N__22051),
            .in2(N__22045),
            .in3(N__43590),
            .lcout(\ALU.madd_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIPVKU_6_LC_4_4_1 .C_ON=1'b0;
    defparam \ALU.r2_RNIPVKU_6_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIPVKU_6_LC_4_4_1 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r2_RNIPVKU_6_LC_4_4_1  (
            .in0(N__29515),
            .in1(N__23463),
            .in2(N__26859),
            .in3(N__23749),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIIH042_6_LC_4_4_2 .C_ON=1'b0;
    defparam \ALU.r6_RNIIH042_6_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIIH042_6_LC_4_4_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNIIH042_6_LC_4_4_2  (
            .in0(N__21993),
            .in1(N__27883),
            .in2(N__22018),
            .in3(N__38793),
            .lcout(),
            .ltout(\ALU.r6_RNIIH042Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI6AI74_6_LC_4_4_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI6AI74_6_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI6AI74_6_LC_4_4_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r4_RNI6AI74_6_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__24642),
            .in2(N__22015),
            .in3(N__21889),
            .lcout(\ALU.b_6 ),
            .ltout(\ALU.b_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2BKQ8_1_6_LC_4_4_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI2BKQ8_1_6_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2BKQ8_1_6_LC_4_4_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \ALU.r4_RNI2BKQ8_1_6_LC_4_4_4  (
            .in0(N__43396),
            .in1(_gnd_net_),
            .in2(N__22012),
            .in3(_gnd_net_),
            .lcout(\ALU.r4_RNI2BKQ8_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_2_N_3L3_LC_4_4_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_2_N_3L3_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_2_N_3L3_LC_4_4_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ALU.mult_g0_2_N_3L3_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(N__37888),
            .in2(_gnd_net_),
            .in3(N__52139),
            .lcout(\ALU.g0_2_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNILJ8Q_6_LC_4_4_6 .C_ON=1'b0;
    defparam \ALU.r0_RNILJ8Q_6_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNILJ8Q_6_LC_4_4_6 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r0_RNILJ8Q_6_LC_4_4_6  (
            .in0(N__23496),
            .in1(N__29514),
            .in2(N__38520),
            .in3(N__26846),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIAP7R1_6_LC_4_4_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIAP7R1_6_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIAP7R1_6_LC_4_4_7 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.r4_RNIAP7R1_6_LC_4_4_7  (
            .in0(N__33783),
            .in1(N__21992),
            .in2(N__21892),
            .in3(N__25360),
            .lcout(\ALU.r4_RNIAP7R1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a9_b_5_LC_4_5_0 .C_ON=1'b0;
    defparam \ALU.mult_a9_b_5_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a9_b_5_LC_4_5_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ALU.mult_a9_b_5_LC_4_5_0  (
            .in0(N__45128),
            .in1(N__30813),
            .in2(N__32265),
            .in3(N__23229),
            .lcout(\ALU.a9_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_14_LC_4_5_1 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_14_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_14_LC_4_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a0_b_14_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__47112),
            .in2(_gnd_net_),
            .in3(N__48915),
            .lcout(\ALU.a0_b_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g2_LC_4_5_2 .C_ON=1'b0;
    defparam \ALU.mult_g2_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g2_LC_4_5_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_g2_LC_4_5_2  (
            .in0(N__48914),
            .in1(N__44489),
            .in2(N__51979),
            .in3(N__23236),
            .lcout(\ALU.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_2_N_4L5_LC_4_5_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_2_N_4L5_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_2_N_4L5_LC_4_5_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ALU.mult_g0_2_N_4L5_LC_4_5_3  (
            .in0(N__44488),
            .in1(N__46009),
            .in2(N__43936),
            .in3(N__46779),
            .lcout(\ALU.g0_2_N_4L5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_134_0_tz_LC_4_5_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_134_0_tz_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_134_0_tz_LC_4_5_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_134_0_tz_LC_4_5_4  (
            .in0(N__46777),
            .in1(N__43899),
            .in2(N__46074),
            .in3(N__44487),
            .lcout(\ALU.madd_134_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_227_LC_4_5_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_227_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_227_LC_4_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_227_LC_4_5_5  (
            .in0(N__51940),
            .in1(N__48913),
            .in2(N__35588),
            .in3(N__48509),
            .lcout(\ALU.madd_130_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_130_LC_4_5_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_130_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_130_LC_4_5_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ALU.mult_madd_130_LC_4_5_6  (
            .in0(N__46776),
            .in1(_gnd_net_),
            .in2(N__46073),
            .in3(N__23113),
            .lcout(\ALU.madd_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_171_sx_LC_4_5_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_171_sx_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_171_sx_LC_4_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_171_sx_LC_4_5_7  (
            .in0(N__43900),
            .in1(N__46778),
            .in2(N__52228),
            .in3(N__46008),
            .lcout(\ALU.madd_171_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_224_0_LC_4_6_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_224_0_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_224_0_LC_4_6_0 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_224_0_LC_4_6_0  (
            .in0(N__51939),
            .in1(N__48342),
            .in2(N__47435),
            .in3(N__48514),
            .lcout(\ALU.madd_224_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_9_s0_c_RNO_LC_4_6_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_9_s0_c_RNO_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_9_s0_c_RNO_LC_4_6_1 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_9_s0_c_RNO_LC_4_6_1  (
            .in0(N__53676),
            .in1(N__52143),
            .in2(N__53232),
            .in3(N__47394),
            .lcout(\ALU.r0_12_prm_6_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_0_l_ofx_LC_4_6_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_0_l_ofx_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_0_l_ofx_LC_4_6_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_madd_axb_0_l_ofx_LC_4_6_2  (
            .in0(N__37828),
            .in1(N__48515),
            .in2(N__46832),
            .in3(N__48921),
            .lcout(\ALU.madd_axb_0_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_0_s1_c_RNO_LC_4_6_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_0_s1_c_RNO_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_0_s1_c_RNO_LC_4_6_4 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_0_s1_c_RNO_LC_4_6_4  (
            .in0(N__37829),
            .in1(N__53675),
            .in2(N__53208),
            .in3(N__48920),
            .lcout(\ALU.r0_12_prm_6_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_213_LC_4_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_213_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_213_LC_4_6_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ALU.mult_madd_213_LC_4_6_5  (
            .in0(N__40932),
            .in1(N__23146),
            .in2(N__23020),
            .in3(N__37827),
            .lcout(\ALU.madd_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a9_b_3_LC_4_6_6 .C_ON=1'b0;
    defparam \ALU.mult_a9_b_3_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a9_b_3_LC_4_6_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ALU.mult_a9_b_3_LC_4_6_6  (
            .in0(N__44342),
            .in1(N__30814),
            .in2(N__36783),
            .in3(N__23228),
            .lcout(\ALU.a9_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_167_0_LC_4_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_167_0_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_167_0_LC_4_6_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_167_0_LC_4_6_7  (
            .in0(N__45988),
            .in1(N__37826),
            .in2(N__51806),
            .in3(N__43920),
            .lcout(\ALU.madd_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNILTKU_5_LC_4_7_0 .C_ON=1'b0;
    defparam \ALU.r2_RNILTKU_5_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNILTKU_5_LC_4_7_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \ALU.r2_RNILTKU_5_LC_4_7_0  (
            .in0(N__23774),
            .in1(N__33140),
            .in2(N__24922),
            .in3(N__24138),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIBP2O1_5_LC_4_7_1 .C_ON=1'b0;
    defparam \ALU.r6_RNIBP2O1_5_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIBP2O1_5_LC_4_7_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.r6_RNIBP2O1_5_LC_4_7_1  (
            .in0(N__24032),
            .in1(N__23964),
            .in2(N__22174),
            .in3(N__26832),
            .lcout(\ALU.r6_RNIBP2O1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIFAMP_5_LC_4_7_2 .C_ON=1'b0;
    defparam \ALU.r0_RNIFAMP_5_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIFAMP_5_LC_4_7_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNIFAMP_5_LC_4_7_2  (
            .in0(N__22316),
            .in1(N__33303),
            .in2(N__37129),
            .in3(N__33203),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI0QNE1_5_LC_4_7_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI0QNE1_5_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI0QNE1_5_LC_4_7_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNI0QNE1_5_LC_4_7_3  (
            .in0(N__33141),
            .in1(N__25927),
            .in2(N__22171),
            .in3(N__25391),
            .lcout(),
            .ltout(\ALU.r4_RNI0QNE1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKI4F3_5_LC_4_7_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIKI4F3_5_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKI4F3_5_LC_4_7_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.r4_RNIKI4F3_5_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__22168),
            .in2(N__22162),
            .in3(N__24710),
            .lcout(\ALU.b_5 ),
            .ltout(\ALU.b_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI8B628_1_5_LC_4_7_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI8B628_1_5_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI8B628_1_5_LC_4_7_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \ALU.r4_RNI8B628_1_5_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22264),
            .in3(N__45512),
            .lcout(\ALU.r4_RNI8B628_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_5_LC_4_7_6 .C_ON=1'b0;
    defparam \ALU.r0_5_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_5_LC_4_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_5_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37209),
            .lcout(r0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56263),
            .ce(N__49739),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIPK3D2_9_LC_4_8_0 .C_ON=1'b0;
    defparam \ALU.r6_RNIPK3D2_9_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIPK3D2_9_LC_4_8_0 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ALU.r6_RNIPK3D2_9_LC_4_8_0  (
            .in0(N__22253),
            .in1(N__30927),
            .in2(N__27799),
            .in3(N__23419),
            .lcout(\ALU.r6_RNIPK3D2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_9_LC_4_8_1 .C_ON=1'b0;
    defparam \ALU.r6_9_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_9_LC_4_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_9_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34032),
            .lcout(r6_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56267),
            .ce(N__45853),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_1_LC_4_8_2.C_ON=1'b0;
    defparam TXbuffer_RNO_7_1_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_1_LC_4_8_2.LUT_INIT=16'b0101010100100111;
    LogicCell40 TXbuffer_RNO_7_1_LC_4_8_2 (
            .in0(N__30386),
            .in1(N__31147),
            .in2(N__35092),
            .in3(N__30038),
            .lcout(),
            .ltout(TXbuffer_18_3_ns_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_1_LC_4_8_3.C_ON=1'b0;
    defparam TXbuffer_RNO_5_1_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_1_LC_4_8_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_5_1_LC_4_8_3 (
            .in0(N__30039),
            .in1(N__34401),
            .in2(N__22261),
            .in3(N__34369),
            .lcout(),
            .ltout(TXbuffer_RNO_5Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_1_LC_4_8_4.C_ON=1'b0;
    defparam TXbuffer_RNO_2_1_LC_4_8_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_1_LC_4_8_4.LUT_INIT=16'b0100010101100111;
    LogicCell40 TXbuffer_RNO_2_1_LC_4_8_4 (
            .in0(N__29675),
            .in1(N__49969),
            .in2(N__22258),
            .in3(N__22237),
            .lcout(TXbuffer_18_15_ns_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_1_LC_4_8_5.C_ON=1'b0;
    defparam TXbuffer_RNO_8_1_LC_4_8_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_1_LC_4_8_5.LUT_INIT=16'b0000101101011011;
    LogicCell40 TXbuffer_RNO_8_1_LC_4_8_5 (
            .in0(N__30036),
            .in1(N__28662),
            .in2(N__30398),
            .in3(N__23706),
            .lcout(),
            .ltout(TXbuffer_18_6_ns_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_1_LC_4_8_6.C_ON=1'b0;
    defparam TXbuffer_RNO_6_1_LC_4_8_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_1_LC_4_8_6.LUT_INIT=16'b1100101100001011;
    LogicCell40 TXbuffer_RNO_6_1_LC_4_8_6 (
            .in0(N__22254),
            .in1(N__30037),
            .in2(N__22240),
            .in3(N__29396),
            .lcout(TXbuffer_RNO_6Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_1_LC_4_8_7 .C_ON=1'b0;
    defparam \ALU.r6_1_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_1_LC_4_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r6_1_LC_4_8_7  (
            .in0(N__42163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56267),
            .ce(N__45853),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIG3U21_5_LC_4_9_0 .C_ON=1'b0;
    defparam \ALU.r0_RNIG3U21_5_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIG3U21_5_LC_4_9_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.r0_RNIG3U21_5_LC_4_9_0  (
            .in0(N__28788),
            .in1(N__22323),
            .in2(N__37124),
            .in3(N__30557),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI24Q22_5_LC_4_9_1 .C_ON=1'b0;
    defparam \ALU.r4_RNI24Q22_5_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI24Q22_5_LC_4_9_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r4_RNI24Q22_5_LC_4_9_1  (
            .in0(N__25926),
            .in1(N__25393),
            .in2(N__22300),
            .in3(N__25597),
            .lcout(\ALU.r4_RNI24Q22Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_0_rep2_LC_4_9_2.C_ON=1'b0;
    defparam a_0_rep2_LC_4_9_2.SEQ_MODE=4'b1000;
    defparam a_0_rep2_LC_4_9_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 a_0_rep2_LC_4_9_2 (
            .in0(N__28791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_0_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56271),
            .ce(N__56044),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNICBU71_10_LC_4_9_3 .C_ON=1'b0;
    defparam \ALU.r2_RNICBU71_10_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNICBU71_10_LC_4_9_3 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.r2_RNICBU71_10_LC_4_9_3  (
            .in0(N__30558),
            .in1(N__22289),
            .in2(N__22389),
            .in3(N__28789),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIP3372_10_LC_4_9_4 .C_ON=1'b0;
    defparam \ALU.r6_RNIP3372_10_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIP3372_10_LC_4_9_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNIP3372_10_LC_4_9_4  (
            .in0(N__30912),
            .in1(N__22679),
            .in2(N__22273),
            .in3(N__22568),
            .lcout(\ALU.r6_RNIP3372Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIEDU71_11_LC_4_9_5 .C_ON=1'b0;
    defparam \ALU.r2_RNIEDU71_11_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIEDU71_11_LC_4_9_5 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.r2_RNIEDU71_11_LC_4_9_5  (
            .in0(N__30559),
            .in1(N__24815),
            .in2(N__22363),
            .in3(N__28790),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIT7372_11_LC_4_9_6 .C_ON=1'b0;
    defparam \ALU.r6_RNIT7372_11_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIT7372_11_LC_4_9_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNIT7372_11_LC_4_9_6  (
            .in0(N__30913),
            .in1(N__22650),
            .in2(N__22270),
            .in3(N__24767),
            .lcout(),
            .ltout(\ALU.r6_RNIT7372Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI8VFH4_11_LC_4_9_7 .C_ON=1'b0;
    defparam \ALU.r5_RNI8VFH4_11_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI8VFH4_11_LC_4_9_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r5_RNI8VFH4_11_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__29202),
            .in2(N__22267),
            .in3(N__23671),
            .lcout(\ALU.a_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINJA71_7_LC_4_10_0 .C_ON=1'b0;
    defparam \ALU.r2_RNINJA71_7_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINJA71_7_LC_4_10_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNINJA71_7_LC_4_10_0  (
            .in0(N__22406),
            .in1(N__30570),
            .in2(N__22482),
            .in3(N__25004),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIGC3D2_7_LC_4_10_1 .C_ON=1'b0;
    defparam \ALU.r6_RNIGC3D2_7_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIGC3D2_7_LC_4_10_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIGC3D2_7_LC_4_10_1  (
            .in0(N__27842),
            .in1(N__38681),
            .in2(N__22453),
            .in3(N__30885),
            .lcout(\ALU.r6_RNIGC3D2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_7_LC_4_10_2 .C_ON=1'b0;
    defparam \ALU.r2_7_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_7_LC_4_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_7_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38754),
            .lcout(r2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56276),
            .ce(N__47690),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIP1LU_7_LC_4_10_3 .C_ON=1'b0;
    defparam \ALU.r2_RNIP1LU_7_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIP1LU_7_LC_4_10_3 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \ALU.r2_RNIP1LU_7_LC_4_10_3  (
            .in0(N__33139),
            .in1(N__24923),
            .in2(N__22481),
            .in3(N__22407),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIJ13O1_7_LC_4_10_4 .C_ON=1'b0;
    defparam \ALU.r6_RNIJ13O1_7_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIJ13O1_7_LC_4_10_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.r6_RNIJ13O1_7_LC_4_10_4  (
            .in0(N__38682),
            .in1(N__27843),
            .in2(N__22450),
            .in3(N__26850),
            .lcout(\ALU.r6_RNIJ13O1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_7_LC_4_10_5.C_ON=1'b0;
    defparam TXbuffer_RNO_8_7_LC_4_10_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_7_LC_4_10_5.LUT_INIT=16'b0001000110101111;
    LogicCell40 TXbuffer_RNO_8_7_LC_4_10_5 (
            .in0(N__30044),
            .in1(N__22435),
            .in2(N__22411),
            .in3(N__30305),
            .lcout(),
            .ltout(TXbuffer_18_6_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_7_LC_4_10_6.C_ON=1'b0;
    defparam TXbuffer_RNO_6_7_LC_4_10_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_7_LC_4_10_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 TXbuffer_RNO_6_7_LC_4_10_6 (
            .in0(N__38683),
            .in1(N__30045),
            .in2(N__22393),
            .in3(N__22534),
            .lcout(TXbuffer_RNO_6Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r3_0_LC_4_11_0 .C_ON=1'b0;
    defparam \ALU.r3_0_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_0_LC_4_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_0_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35018),
            .lcout(r3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_10_LC_4_11_1 .C_ON=1'b0;
    defparam \ALU.r3_10_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_10_LC_4_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_10_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28189),
            .lcout(r3_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_11_LC_4_11_2 .C_ON=1'b0;
    defparam \ALU.r3_11_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_11_LC_4_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_11_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26155),
            .lcout(r3_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_15_LC_4_11_3 .C_ON=1'b0;
    defparam \ALU.r3_15_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_15_LC_4_11_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \ALU.r3_15_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25993),
            .in3(_gnd_net_),
            .lcout(r3_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_7_LC_4_11_4 .C_ON=1'b0;
    defparam \ALU.r3_7_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_7_LC_4_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_7_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38755),
            .lcout(r3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_8_LC_4_11_5 .C_ON=1'b0;
    defparam \ALU.r3_8_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_8_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_8_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39525),
            .lcout(r3_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_9_LC_4_11_6 .C_ON=1'b0;
    defparam \ALU.r3_9_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_9_LC_4_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_9_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34026),
            .lcout(r3_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_1_LC_4_11_7 .C_ON=1'b0;
    defparam \ALU.r3_1_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_1_LC_4_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_1_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42155),
            .lcout(r3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56281),
            .ce(N__47755),
            .sr(_gnd_net_));
    defparam \ALU.r3_6_LC_4_12_0 .C_ON=1'b0;
    defparam \ALU.r3_6_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_6_LC_4_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_6_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38878),
            .lcout(r3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56285),
            .ce(N__47762),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_6_LC_4_12_1.C_ON=1'b0;
    defparam TXbuffer_RNO_4_6_LC_4_12_1.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_6_LC_4_12_1.LUT_INIT=16'b0001000110101111;
    LogicCell40 TXbuffer_RNO_4_6_LC_4_12_1 (
            .in0(N__29968),
            .in1(N__25820),
            .in2(N__23453),
            .in3(N__30303),
            .lcout(),
            .ltout(TXbuffer_18_13_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_6_LC_4_12_2.C_ON=1'b0;
    defparam TXbuffer_RNO_1_6_LC_4_12_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_6_LC_4_12_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_1_6_LC_4_12_2 (
            .in0(N__29974),
            .in1(N__25796),
            .in2(N__22456),
            .in3(N__27882),
            .lcout(TXbuffer_RNO_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r3_14_LC_4_12_3 .C_ON=1'b0;
    defparam \ALU.r3_14_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_14_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_14_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28312),
            .lcout(r3_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56285),
            .ce(N__47762),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_2_LC_4_12_4.C_ON=1'b0;
    defparam TXbuffer_RNO_7_2_LC_4_12_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_2_LC_4_12_4.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_7_2_LC_4_12_4 (
            .in0(N__29972),
            .in1(N__28121),
            .in2(N__30354),
            .in3(N__33418),
            .lcout(),
            .ltout(TXbuffer_18_3_ns_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_2_LC_4_12_5.C_ON=1'b0;
    defparam TXbuffer_RNO_5_2_LC_4_12_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_2_LC_4_12_5.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_5_2_LC_4_12_5 (
            .in0(N__29967),
            .in1(N__25478),
            .in2(N__22606),
            .in3(N__34333),
            .lcout(TXbuffer_RNO_5Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_4_LC_4_12_6.C_ON=1'b0;
    defparam TXbuffer_RNO_7_4_LC_4_12_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_4_LC_4_12_6.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_7_4_LC_4_12_6 (
            .in0(N__29973),
            .in1(N__28374),
            .in2(N__30355),
            .in3(N__33511),
            .lcout(TXbuffer_18_3_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_0_LC_4_13_0 .C_ON=1'b0;
    defparam \ALU.r6_0_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_0_LC_4_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35025),
            .lcout(r6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_10_LC_4_13_1 .C_ON=1'b0;
    defparam \ALU.r6_10_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_10_LC_4_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_10_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28191),
            .lcout(r6_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_11_LC_4_13_2 .C_ON=1'b0;
    defparam \ALU.r6_11_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_11_LC_4_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r6_11_LC_4_13_2  (
            .in0(N__26156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r6_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_12_LC_4_13_3 .C_ON=1'b0;
    defparam \ALU.r6_12_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_12_LC_4_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_12_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28440),
            .lcout(r6_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_13_LC_4_13_4 .C_ON=1'b0;
    defparam \ALU.r6_13_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_13_LC_4_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_13_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26277),
            .lcout(r6_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_14_LC_4_13_5 .C_ON=1'b0;
    defparam \ALU.r6_14_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_14_LC_4_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_14_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28309),
            .lcout(r6_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_15_LC_4_13_6 .C_ON=1'b0;
    defparam \ALU.r6_15_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_15_LC_4_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_15_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25976),
            .lcout(r6_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r6_5_LC_4_13_7 .C_ON=1'b0;
    defparam \ALU.r6_5_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_5_LC_4_13_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ALU.r6_5_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__37211),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56289),
            .ce(N__45842),
            .sr(_gnd_net_));
    defparam \ALU.r7_0_LC_4_14_0 .C_ON=1'b0;
    defparam \ALU.r7_0_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_0_LC_4_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_0_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35026),
            .lcout(r7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_10_LC_4_14_1 .C_ON=1'b0;
    defparam \ALU.r7_10_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_10_LC_4_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_10_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28190),
            .lcout(r7_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_11_LC_4_14_2 .C_ON=1'b0;
    defparam \ALU.r7_11_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_11_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_11_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26176),
            .lcout(r7_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_12_LC_4_14_3 .C_ON=1'b0;
    defparam \ALU.r7_12_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_12_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_12_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28446),
            .lcout(r7_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_13_LC_4_14_4 .C_ON=1'b0;
    defparam \ALU.r7_13_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_13_LC_4_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_13_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26279),
            .lcout(r7_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_14_LC_4_14_5 .C_ON=1'b0;
    defparam \ALU.r7_14_LC_4_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_14_LC_4_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_14_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28311),
            .lcout(r7_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_15_LC_4_14_6 .C_ON=1'b0;
    defparam \ALU.r7_15_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_15_LC_4_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_15_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25972),
            .lcout(r7_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam \ALU.r7_5_LC_4_14_7 .C_ON=1'b0;
    defparam \ALU.r7_5_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_5_LC_4_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r7_5_LC_4_14_7  (
            .in0(N__37212),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56293),
            .ce(N__45895),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_6_LC_4_15_0.C_ON=1'b0;
    defparam TXbuffer_RNO_3_6_LC_4_15_0.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_6_LC_4_15_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_3_6_LC_4_15_0 (
            .in0(N__29932),
            .in1(N__28246),
            .in2(N__30324),
            .in3(N__38524),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_6_LC_4_15_1.C_ON=1'b0;
    defparam TXbuffer_RNO_0_6_LC_4_15_1.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_6_LC_4_15_1.LUT_INIT=16'b1000111110000011;
    LogicCell40 TXbuffer_RNO_0_6_LC_4_15_1 (
            .in0(N__33784),
            .in1(N__29933),
            .in2(N__22756),
            .in3(N__26025),
            .lcout(),
            .ltout(TXbuffer_RNO_0Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_6_LC_4_15_2.C_ON=1'b0;
    defparam TXbuffer_6_LC_4_15_2.SEQ_MODE=4'b1000;
    defparam TXbuffer_6_LC_4_15_2.LUT_INIT=16'b1010000011011101;
    LogicCell40 TXbuffer_6_LC_4_15_2 (
            .in0(N__49889),
            .in1(N__22753),
            .in2(N__22741),
            .in3(N__22726),
            .lcout(TXbufferZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56298),
            .ce(N__56038),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_6_LC_4_15_3.C_ON=1'b0;
    defparam TXbuffer_RNO_6_6_LC_4_15_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_6_LC_4_15_3.LUT_INIT=16'b1110010001010101;
    LogicCell40 TXbuffer_RNO_6_6_LC_4_15_3 (
            .in0(N__22738),
            .in1(N__25764),
            .in2(N__38800),
            .in3(N__29931),
            .lcout(),
            .ltout(TXbuffer_RNO_6Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_6_LC_4_15_4.C_ON=1'b0;
    defparam TXbuffer_RNO_2_6_LC_4_15_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_6_LC_4_15_4.LUT_INIT=16'b0100011001010111;
    LogicCell40 TXbuffer_RNO_2_6_LC_4_15_4 (
            .in0(N__29668),
            .in1(N__49888),
            .in2(N__22729),
            .in3(N__22717),
            .lcout(TXbuffer_18_15_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_6_LC_4_15_5.C_ON=1'b0;
    defparam TXbuffer_RNO_7_6_LC_4_15_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_6_LC_4_15_5.LUT_INIT=16'b0000001111011101;
    LogicCell40 TXbuffer_RNO_7_6_LC_4_15_5 (
            .in0(N__23497),
            .in1(N__29929),
            .in2(N__25723),
            .in3(N__30269),
            .lcout(),
            .ltout(TXbuffer_18_3_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_6_LC_4_15_6.C_ON=1'b0;
    defparam TXbuffer_RNO_5_6_LC_4_15_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_6_LC_4_15_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_5_6_LC_4_15_6 (
            .in0(N__29930),
            .in1(N__25888),
            .in2(N__22720),
            .in3(N__25356),
            .lcout(TXbuffer_RNO_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_11_s1_c_RNO_LC_4_16_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_11_s1_c_RNO_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_11_s1_c_RNO_LC_4_16_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_11_s1_c_RNO_LC_4_16_0  (
            .in0(N__54054),
            .in1(N__53003),
            .in2(N__54779),
            .in3(N__40968),
            .lcout(\ALU.r0_12_prm_4_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIAFVE5_11_LC_4_16_1 .C_ON=1'b0;
    defparam \ALU.r5_RNIAFVE5_11_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIAFVE5_11_LC_4_16_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r5_RNIAFVE5_11_LC_4_16_1  (
            .in0(N__40965),
            .in1(N__54596),
            .in2(N__53166),
            .in3(N__54052),
            .lcout(\ALU.r5_RNIAFVE5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_11_s0_c_RNO_LC_4_16_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_11_s0_c_RNO_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_11_s0_c_RNO_LC_4_16_2 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_11_s0_c_RNO_LC_4_16_2  (
            .in0(N__54595),
            .in1(N__35579),
            .in2(N__53169),
            .in3(N__40966),
            .lcout(\ALU.r0_12_prm_5_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNISP2L9_0_12_LC_4_16_3 .C_ON=1'b0;
    defparam \ALU.r5_RNISP2L9_0_12_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNISP2L9_0_12_LC_4_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.r5_RNISP2L9_0_12_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__39830),
            .in2(_gnd_net_),
            .in3(N__41329),
            .lcout(\ALU.r5_RNISP2L9_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_11_s0_c_RNO_LC_4_16_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_11_s0_c_RNO_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_11_s0_c_RNO_LC_4_16_4 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_11_s0_c_RNO_LC_4_16_4  (
            .in0(N__54051),
            .in1(N__35578),
            .in2(N__53168),
            .in3(N__40964),
            .lcout(\ALU.r0_12_prm_6_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_13_s1_c_RNO_LC_4_16_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_13_s1_c_RNO_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_13_s1_c_RNO_LC_4_16_5 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_13_s1_c_RNO_LC_4_16_5  (
            .in0(N__52996),
            .in1(N__35392),
            .in2(_gnd_net_),
            .in3(N__41464),
            .lcout(\ALU.r0_12_prm_7_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_11_s0_c_RNO_LC_4_16_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_11_s0_c_RNO_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_11_s0_c_RNO_LC_4_16_6 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_11_s0_c_RNO_LC_4_16_6  (
            .in0(N__53004),
            .in1(N__35577),
            .in2(_gnd_net_),
            .in3(N__40963),
            .lcout(\ALU.r0_12_prm_7_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_11_s1_c_RNO_LC_4_16_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_11_s1_c_RNO_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_11_s1_c_RNO_LC_4_16_7 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_11_s1_c_RNO_LC_4_16_7  (
            .in0(N__40967),
            .in1(N__54053),
            .in2(N__53167),
            .in3(N__35580),
            .lcout(\ALU.r0_12_prm_6_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_5_LC_4_17_0.C_ON=1'b0;
    defparam TXbuffer_RNO_5_5_LC_4_17_0.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_5_LC_4_17_0.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_5_5_LC_4_17_0 (
            .in0(N__29989),
            .in1(N__25426),
            .in2(N__22768),
            .in3(N__25392),
            .lcout(TXbuffer_RNO_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_5_LC_4_17_2.C_ON=1'b0;
    defparam TXbuffer_RNO_8_5_LC_4_17_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_5_LC_4_17_2.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_8_5_LC_4_17_2 (
            .in0(N__29988),
            .in1(N__23917),
            .in2(N__30359),
            .in3(N__23776),
            .lcout(TXbuffer_18_6_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_5_LC_4_17_5.C_ON=1'b0;
    defparam TXbuffer_RNO_4_5_LC_4_17_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_5_LC_4_17_5.LUT_INIT=16'b0101010100100111;
    LogicCell40 TXbuffer_RNO_4_5_LC_4_17_5 (
            .in0(N__30317),
            .in1(N__24101),
            .in2(N__24128),
            .in3(N__29990),
            .lcout(TXbuffer_18_13_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_105_LC_5_1_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_105_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_105_LC_5_1_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ALU.mult_madd_105_LC_5_1_1  (
            .in0(N__22993),
            .in1(N__48949),
            .in2(_gnd_net_),
            .in3(N__46363),
            .lcout(\ALU.madd_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a4_b_4_LC_5_1_2 .C_ON=1'b0;
    defparam \ALU.mult_a4_b_4_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a4_b_4_LC_5_1_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a4_b_4_LC_5_1_2  (
            .in0(N__32472),
            .in1(N__32373),
            .in2(N__36782),
            .in3(N__40520),
            .lcout(\ALU.a4_b_4 ),
            .ltout(\ALU.a4_b_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_104_LC_5_1_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_104_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_104_LC_5_1_3 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_104_LC_5_1_3  (
            .in0(N__24183),
            .in1(N__45232),
            .in2(N__22846),
            .in3(N__49350),
            .lcout(\ALU.madd_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_68_LC_5_1_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_68_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_68_LC_5_1_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALU.mult_madd_68_LC_5_1_4  (
            .in0(N__45504),
            .in1(N__24237),
            .in2(_gnd_net_),
            .in3(N__43930),
            .lcout(\ALU.madd_68 ),
            .ltout(\ALU.madd_68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_82_0_LC_5_1_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_82_0_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_82_0_LC_5_1_5 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \ALU.mult_madd_82_0_LC_5_1_5  (
            .in0(N__24166),
            .in1(N__43644),
            .in2(N__22822),
            .in3(N__48513),
            .lcout(\ALU.madd_82_0 ),
            .ltout(\ALU.madd_82_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_119_LC_5_1_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_119_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_119_LC_5_1_6 .LUT_INIT=16'b1111111011001000;
    LogicCell40 \ALU.mult_madd_119_LC_5_1_6  (
            .in0(N__24226),
            .in1(N__24217),
            .in2(N__22819),
            .in3(N__24205),
            .lcout(\ALU.madd_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_100_LC_5_1_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_100_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_100_LC_5_1_7 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_100_LC_5_1_7  (
            .in0(N__24184),
            .in1(N__45233),
            .in2(N__38451),
            .in3(N__49351),
            .lcout(\ALU.madd_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_68_0_LC_5_2_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_68_0_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_68_0_LC_5_2_0 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_68_0_LC_5_2_0  (
            .in0(N__37897),
            .in1(N__44518),
            .in2(N__43355),
            .in3(N__46745),
            .lcout(\ALU.madd_68_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_0_LC_5_2_1 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_0_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_0_LC_5_2_1 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a5_b_0_LC_5_2_1  (
            .in0(N__29079),
            .in1(N__29005),
            .in2(N__32186),
            .in3(N__37898),
            .lcout(\ALU.a5_b_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIS02J4_6_LC_5_2_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIS02J4_6_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIS02J4_6_LC_5_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIS02J4_6_LC_5_2_2  (
            .in0(N__29219),
            .in1(N__26508),
            .in2(_gnd_net_),
            .in3(N__26436),
            .lcout(\ALU.a_6 ),
            .ltout(\ALU.a_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_72_0_tz_LC_5_2_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_72_0_tz_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_72_0_tz_LC_5_2_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_72_0_tz_LC_5_2_3  (
            .in0(N__46744),
            .in1(N__45454),
            .in2(N__22801),
            .in3(N__43886),
            .lcout(\ALU.madd_72_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g3_LC_5_2_4 .C_ON=1'b0;
    defparam \ALU.mult_g3_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g3_LC_5_2_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \ALU.mult_g3_LC_5_2_4  (
            .in0(N__49277),
            .in1(N__45201),
            .in2(N__24469),
            .in3(N__40485),
            .lcout(\ALU.g3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_71_LC_5_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_71_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_71_LC_5_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_71_LC_5_2_5  (
            .in0(N__46746),
            .in1(N__43279),
            .in2(N__45495),
            .in3(N__43887),
            .lcout(),
            .ltout(\ALU.madd_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_72_LC_5_2_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_72_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_72_LC_5_2_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_madd_72_LC_5_2_6  (
            .in0(N__37899),
            .in1(N__22948),
            .in2(N__22942),
            .in3(N__44519),
            .lcout(\ALU.madd_72 ),
            .ltout(\ALU.madd_72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_110_LC_5_2_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_110_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_110_LC_5_2_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_110_LC_5_2_7  (
            .in0(N__22927),
            .in1(_gnd_net_),
            .in2(N__22909),
            .in3(N__22906),
            .lcout(\ALU.madd_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIVA4L3_8_LC_5_3_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIVA4L3_8_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIVA4L3_8_LC_5_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIVA4L3_8_LC_5_3_0  (
            .in0(N__24623),
            .in1(N__23515),
            .in2(_gnd_net_),
            .in3(N__22981),
            .lcout(\ALU.b_8 ),
            .ltout(\ALU.b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_143_LC_5_3_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_143_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_143_LC_5_3_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_143_LC_5_3_1  (
            .in0(N__44675),
            .in1(N__48235),
            .in2(N__22891),
            .in3(N__48472),
            .lcout(\ALU.madd_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_8_s0_c_RNO_LC_5_3_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_8_s0_c_RNO_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_8_s0_c_RNO_LC_5_3_2 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_8_s0_c_RNO_LC_5_3_2  (
            .in0(N__46317),
            .in1(N__53898),
            .in2(N__53068),
            .in3(N__46080),
            .lcout(\ALU.r0_12_prm_6_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_222_LC_5_3_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_222_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_222_LC_5_3_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_222_LC_5_3_3  (
            .in0(N__44678),
            .in1(N__46316),
            .in2(N__42755),
            .in3(N__49236),
            .lcout(),
            .ltout(\ALU.madd_127_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_223_LC_5_3_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_223_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_223_LC_5_3_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_madd_223_LC_5_3_4  (
            .in0(N__45505),
            .in1(N__43520),
            .in2(N__22876),
            .in3(N__22999),
            .lcout(\ALU.madd_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_223_0_tz_LC_5_3_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_223_0_tz_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_223_0_tz_LC_5_3_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_madd_223_0_tz_LC_5_3_5  (
            .in0(N__44677),
            .in1(N__46315),
            .in2(N__42754),
            .in3(N__49237),
            .lcout(\ALU.madd_223_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_105_0_LC_5_3_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_105_0_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_105_0_LC_5_3_6 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_105_0_LC_5_3_6  (
            .in0(N__48473),
            .in1(N__43521),
            .in2(N__48292),
            .in3(N__44676),
            .lcout(\ALU.madd_105_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIU5NK1_8_LC_5_3_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIU5NK1_8_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIU5NK1_8_LC_5_3_7 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.r4_RNIU5NK1_8_LC_5_3_7  (
            .in0(N__26852),
            .in1(N__34069),
            .in2(N__33727),
            .in3(N__23140),
            .lcout(\ALU.r4_RNIU5NK1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2THO8_0_3_LC_5_4_0 .C_ON=1'b0;
    defparam \ALU.r4_RNI2THO8_0_3_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2THO8_0_3_LC_5_4_0 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \ALU.r4_RNI2THO8_0_3_LC_5_4_0  (
            .in0(N__31911),
            .in1(N__44252),
            .in2(N__32264),
            .in3(N__31824),
            .lcout(\ALU.un9_addsub_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIUES39_0_1_LC_5_4_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIUES39_0_1_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIUES39_0_1_LC_5_4_1 .LUT_INIT=16'b0101001110101100;
    LogicCell40 \ALU.r4_RNIUES39_0_1_LC_5_4_1  (
            .in0(N__31631),
            .in1(N__31721),
            .in2(N__32263),
            .in3(N__46672),
            .lcout(),
            .ltout(\ALU.un9_addsub_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI90J9E_1_LC_5_4_2 .C_ON=1'b0;
    defparam \ALU.r4_RNI90J9E_1_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI90J9E_1_LC_5_4_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.r4_RNI90J9E_1_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22975),
            .in3(N__48505),
            .lcout(\ALU.r4_RNI90J9EZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a7_b_3_LC_5_4_3 .C_ON=1'b0;
    defparam \ALU.mult_a7_b_3_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a7_b_3_LC_5_4_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a7_b_3_LC_5_4_3  (
            .in0(N__44251),
            .in1(N__23101),
            .in2(N__36685),
            .in3(N__30715),
            .lcout(\ALU.a7_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJPM55_2_LC_5_4_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIJPM55_2_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJPM55_2_LC_5_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIJPM55_2_LC_5_4_4  (
            .in0(N__27754),
            .in1(N__32656),
            .in2(_gnd_net_),
            .in3(N__32574),
            .lcout(\ALU.a_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIBHM55_1_LC_5_4_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIBHM55_1_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIBHM55_1_LC_5_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r4_RNIBHM55_1_LC_5_4_5  (
            .in0(N__31630),
            .in1(N__31720),
            .in2(_gnd_net_),
            .in3(N__27753),
            .lcout(\ALU.a_1 ),
            .ltout(\ALU.a_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_228_0_tz_LC_5_4_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_228_0_tz_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_228_0_tz_LC_5_4_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_madd_228_0_tz_LC_5_4_6  (
            .in0(N__35581),
            .in1(N__51975),
            .in2(N__22966),
            .in3(N__48759),
            .lcout(\ALU.madd_228_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIUES39_1_LC_5_4_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIUES39_1_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIUES39_1_LC_5_4_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r4_RNIUES39_1_LC_5_4_7  (
            .in0(N__31632),
            .in1(N__31722),
            .in2(N__46775),
            .in3(N__32245),
            .lcout(\ALU.r4_RNIUES39Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIURI55_9_LC_5_5_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIURI55_9_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIURI55_9_LC_5_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r4_RNIURI55_9_LC_5_5_0  (
            .in0(N__27751),
            .in1(N__30812),
            .in2(_gnd_net_),
            .in3(N__23224),
            .lcout(\ALU.a_9 ),
            .ltout(\ALU.a_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_9_LC_5_5_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_9_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_9_LC_5_5_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ALU.mult_g0_9_LC_5_5_1  (
            .in0(N__24403),
            .in1(N__32995),
            .in2(N__23131),
            .in3(N__37831),
            .lcout(\ALU.N_675_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIR1GK3_0_LC_5_5_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIR1GK3_0_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIR1GK3_0_LC_5_5_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r4_RNIR1GK3_0_LC_5_5_2  (
            .in0(N__32744),
            .in1(N__24712),
            .in2(_gnd_net_),
            .in3(N__32708),
            .lcout(\ALU.bZ0Z_0 ),
            .ltout(\ALU.bZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_130_0_LC_5_5_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_130_0_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_130_0_LC_5_5_3 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_130_0_LC_5_5_3  (
            .in0(N__43822),
            .in1(N__52102),
            .in2(N__23116),
            .in3(N__44435),
            .lcout(\ALU.madd_130_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIDBI55_7_LC_5_5_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIDBI55_7_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIDBI55_7_LC_5_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIDBI55_7_LC_5_5_4  (
            .in0(N__27750),
            .in1(N__23100),
            .in2(_gnd_net_),
            .in3(N__30711),
            .lcout(\ALU.a_7 ),
            .ltout(\ALU.a_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_133_LC_5_5_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_133_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_133_LC_5_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_133_LC_5_5_5  (
            .in0(N__46670),
            .in1(N__43837),
            .in2(N__23053),
            .in3(N__46055),
            .lcout(\ALU.madd_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_213_0_tz_LC_5_5_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_213_0_tz_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_213_0_tz_LC_5_5_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \ALU.mult_madd_213_0_tz_LC_5_5_6  (
            .in0(N__52104),
            .in1(N__43823),
            .in2(N__51807),
            .in3(N__46671),
            .lcout(\ALU.madd_213_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_209_0_LC_5_5_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_209_0_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_209_0_LC_5_5_7 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_209_0_LC_5_5_7  (
            .in0(N__43821),
            .in1(N__52103),
            .in2(N__40970),
            .in3(N__37830),
            .lcout(\ALU.madd_209_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a8_b_4_LC_5_6_0 .C_ON=1'b0;
    defparam \ALU.mult_a8_b_4_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a8_b_4_LC_5_6_0 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \ALU.mult_a8_b_4_LC_5_6_0  (
            .in0(N__36697),
            .in1(N__40429),
            .in2(N__30621),
            .in3(N__23406),
            .lcout(\ALU.a8_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_7_x1_LC_5_6_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_7_x1_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_7_x1_LC_5_6_1 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \ALU.mult_g0_7_x1_LC_5_6_1  (
            .in0(N__23405),
            .in1(N__30614),
            .in2(N__46754),
            .in3(N__27741),
            .lcout(),
            .ltout(\ALU.g0_7_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_7_ns_LC_5_6_2 .C_ON=1'b0;
    defparam \ALU.mult_g0_7_ns_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_7_ns_LC_5_6_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.mult_g0_7_ns_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23239),
            .in3(N__43860),
            .lcout(\ALU.madd_76_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a9_b_4_LC_5_6_3 .C_ON=1'b0;
    defparam \ALU.mult_a9_b_4_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a9_b_4_LC_5_6_3 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \ALU.mult_a9_b_4_LC_5_6_3  (
            .in0(N__40428),
            .in1(N__30811),
            .in2(N__23230),
            .in3(N__36698),
            .lcout(\ALU.a9_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNILJI55_8_LC_5_6_4 .C_ON=1'b0;
    defparam \ALU.r4_RNILJI55_8_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNILJI55_8_LC_5_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNILJI55_8_LC_5_6_4  (
            .in0(N__27740),
            .in1(N__23404),
            .in2(_gnd_net_),
            .in3(N__30613),
            .lcout(\ALU.a_8 ),
            .ltout(\ALU.a_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNICTFPA_9_LC_5_6_5 .C_ON=1'b0;
    defparam \ALU.r4_RNICTFPA_9_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNICTFPA_9_LC_5_6_5 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.r4_RNICTFPA_9_LC_5_6_5  (
            .in0(N__54128),
            .in1(N__52122),
            .in2(N__23176),
            .in3(N__53811),
            .lcout(\ALU.lshift_3_ns_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_224_LC_5_6_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_224_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_224_LC_5_6_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALU.mult_madd_224_LC_5_6_6  (
            .in0(N__48870),
            .in1(N__23173),
            .in2(_gnd_net_),
            .in3(N__35562),
            .lcout(\ALU.madd_224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_212_LC_5_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_212_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_212_LC_5_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_212_LC_5_6_7  (
            .in0(N__46693),
            .in1(N__52121),
            .in2(N__43914),
            .in3(N__51732),
            .lcout(\ALU.madd_121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI6GLV_8_LC_5_7_0 .C_ON=1'b0;
    defparam \ALU.r0_RNI6GLV_8_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI6GLV_8_LC_5_7_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r0_RNI6GLV_8_LC_5_7_0  (
            .in0(N__39439),
            .in1(N__24906),
            .in2(N__30663),
            .in3(N__33288),
            .lcout(\ALU.b_3_ns_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_0_rep1_LC_5_7_1.C_ON=1'b0;
    defparam b_0_rep1_LC_5_7_1.SEQ_MODE=4'b1000;
    defparam b_0_rep1_LC_5_7_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 b_0_rep1_LC_5_7_1 (
            .in0(N__24909),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_0_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56259),
            .ce(N__56047),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIUF141_2_LC_5_7_2 .C_ON=1'b0;
    defparam \ALU.r2_RNIUF141_2_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIUF141_2_LC_5_7_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r2_RNIUF141_2_LC_5_7_2  (
            .in0(N__23386),
            .in1(N__24905),
            .in2(N__23362),
            .in3(N__33289),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIE5FT1_2_LC_5_7_3 .C_ON=1'b0;
    defparam \ALU.r6_RNIE5FT1_2_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIE5FT1_2_LC_5_7_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNIE5FT1_2_LC_5_7_3  (
            .in0(N__26797),
            .in1(N__28088),
            .in2(N__23332),
            .in3(N__39169),
            .lcout(\ALU.r6_RNIE5FT1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI0I141_3_LC_5_7_4 .C_ON=1'b0;
    defparam \ALU.r2_RNI0I141_3_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI0I141_3_LC_5_7_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r2_RNI0I141_3_LC_5_7_4  (
            .in0(N__24794),
            .in1(N__24907),
            .in2(N__23665),
            .in3(N__33290),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNII9FT1_3_LC_5_7_5 .C_ON=1'b0;
    defparam \ALU.r6_RNII9FT1_3_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNII9FT1_3_LC_5_7_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNII9FT1_3_LC_5_7_5  (
            .in0(N__26798),
            .in1(N__28059),
            .in2(N__23329),
            .in3(N__39132),
            .lcout(\ALU.r6_RNII9FT1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIQB141_0_LC_5_7_6 .C_ON=1'b0;
    defparam \ALU.r2_RNIQB141_0_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIQB141_0_LC_5_7_6 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r2_RNIQB141_0_LC_5_7_6  (
            .in0(N__28740),
            .in1(N__24908),
            .in2(N__28839),
            .in3(N__33291),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI6TET1_0_LC_5_7_7 .C_ON=1'b0;
    defparam \ALU.r6_RNI6TET1_0_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI6TET1_0_LC_5_7_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNI6TET1_0_LC_5_7_7  (
            .in0(N__26799),
            .in1(N__23325),
            .in2(N__23293),
            .in3(N__23290),
            .lcout(\ALU.r6_RNI6TET1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNII5U21_6_LC_5_8_0 .C_ON=1'b0;
    defparam \ALU.r0_RNII5U21_6_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNII5U21_6_LC_5_8_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r0_RNII5U21_6_LC_5_8_0  (
            .in0(N__28781),
            .in1(N__38519),
            .in2(N__30563),
            .in3(N__23483),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI68Q22_6_LC_5_8_1 .C_ON=1'b0;
    defparam \ALU.r4_RNI68Q22_6_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI68Q22_6_LC_5_8_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNI68Q22_6_LC_5_8_1  (
            .in0(N__25569),
            .in1(N__25352),
            .in2(N__23266),
            .in3(N__33770),
            .lcout(\ALU.r4_RNI68Q22Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_6_LC_5_8_2 .C_ON=1'b0;
    defparam \ALU.r0_6_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_6_LC_5_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r0_6_LC_5_8_2  (
            .in0(N__38871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56264),
            .ce(N__49746),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIKFA71_5_LC_5_8_3 .C_ON=1'b0;
    defparam \ALU.r2_RNIKFA71_5_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIKFA71_5_LC_5_8_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIKFA71_5_LC_5_8_3  (
            .in0(N__23775),
            .in1(N__30543),
            .in2(N__24139),
            .in3(N__28784),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIASIB2_5_LC_5_8_4 .C_ON=1'b0;
    defparam \ALU.r6_RNIASIB2_5_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIASIB2_5_LC_5_8_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIASIB2_5_LC_5_8_4  (
            .in0(N__23957),
            .in1(N__24037),
            .in2(N__23467),
            .in3(N__25571),
            .lcout(\ALU.r6_RNIASIB2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIMHA71_6_LC_5_8_5 .C_ON=1'b0;
    defparam \ALU.r2_RNIMHA71_6_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIMHA71_6_LC_5_8_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIMHA71_6_LC_5_8_5  (
            .in0(N__23741),
            .in1(N__30541),
            .in2(N__23464),
            .in3(N__28782),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIE0JB2_6_LC_5_8_6 .C_ON=1'b0;
    defparam \ALU.r6_RNIE0JB2_6_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIE0JB2_6_LC_5_8_6 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIE0JB2_6_LC_5_8_6  (
            .in0(N__27878),
            .in1(N__38786),
            .in2(N__23422),
            .in3(N__25570),
            .lcout(\ALU.r6_RNIE0JB2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNISNA71_9_LC_5_8_7 .C_ON=1'b0;
    defparam \ALU.r2_RNISNA71_9_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNISNA71_9_LC_5_8_7 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNISNA71_9_LC_5_8_7  (
            .in0(N__23705),
            .in1(N__30542),
            .in2(N__27588),
            .in3(N__28783),
            .lcout(\ALU.a_6_ns_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIPLA71_8_LC_5_9_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIPLA71_8_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIPLA71_8_LC_5_9_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIPLA71_8_LC_5_9_0  (
            .in0(N__23564),
            .in1(N__30567),
            .in2(N__23548),
            .in3(N__25003),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIKG3D2_8_LC_5_9_1 .C_ON=1'b0;
    defparam \ALU.r6_RNIKG3D2_8_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIKG3D2_8_LC_5_9_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIKG3D2_8_LC_5_9_1  (
            .in0(N__27824),
            .in1(N__39200),
            .in2(N__23413),
            .in3(N__30915),
            .lcout(\ALU.r6_RNIKG3D2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_8_LC_5_9_2 .C_ON=1'b0;
    defparam \ALU.r2_8_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_8_LC_5_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_8_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39526),
            .lcout(r2_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56268),
            .ce(N__47708),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIR3LU_8_LC_5_9_3 .C_ON=1'b0;
    defparam \ALU.r2_RNIR3LU_8_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIR3LU_8_LC_5_9_3 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.r2_RNIR3LU_8_LC_5_9_3  (
            .in0(N__24924),
            .in1(N__33112),
            .in2(N__23571),
            .in3(N__23546),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIN53O1_8_LC_5_9_4 .C_ON=1'b0;
    defparam \ALU.r6_RNIN53O1_8_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIN53O1_8_LC_5_9_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.r6_RNIN53O1_8_LC_5_9_4  (
            .in0(N__39201),
            .in1(N__27825),
            .in2(N__23518),
            .in3(N__26851),
            .lcout(\ALU.r6_RNIN53O1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIQUF71_1_LC_5_9_5 .C_ON=1'b0;
    defparam \ALU.r2_RNIQUF71_1_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIQUF71_1_LC_5_9_5 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.r2_RNIQUF71_1_LC_5_9_5  (
            .in0(N__25002),
            .in1(N__28652),
            .in2(N__28700),
            .in3(N__31062),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI7B8D2_1_LC_5_9_6 .C_ON=1'b0;
    defparam \ALU.r6_RNI7B8D2_1_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI7B8D2_1_LC_5_9_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNI7B8D2_1_LC_5_9_6  (
            .in0(N__30914),
            .in1(N__29439),
            .in2(N__23506),
            .in3(N__29406),
            .lcout(\ALU.r6_RNI7B8D2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_1_LC_5_9_7 .C_ON=1'b0;
    defparam \ALU.r2_1_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_1_LC_5_9_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ALU.r2_1_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__42156),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56268),
            .ce(N__47708),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIMIB71_10_LC_5_10_0 .C_ON=1'b0;
    defparam \ALU.r1_RNIMIB71_10_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIMIB71_10_LC_5_10_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r1_RNIMIB71_10_LC_5_10_0  (
            .in0(N__28122),
            .in1(N__25000),
            .in2(N__27962),
            .in3(N__31061),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIVQN52_10_LC_5_10_1 .C_ON=1'b0;
    defparam \ALU.r5_RNIVQN52_10_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIVQN52_10_LC_5_10_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r5_RNIVQN52_10_LC_5_10_1  (
            .in0(N__27932),
            .in1(N__25479),
            .in2(N__23503),
            .in3(N__30888),
            .lcout(\ALU.r5_RNIVQN52Z0Z_10 ),
            .ltout(\ALU.r5_RNIVQN52Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI0NFH4_10_LC_5_10_2 .C_ON=1'b0;
    defparam \ALU.r5_RNI0NFH4_10_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI0NFH4_10_LC_5_10_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.r5_RNI0NFH4_10_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__29156),
            .in2(N__23500),
            .in3(N__36795),
            .lcout(\ALU.a_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_0_rep1_LC_5_10_3.C_ON=1'b0;
    defparam a_0_rep1_LC_5_10_3.SEQ_MODE=4'b1000;
    defparam a_0_rep1_LC_5_10_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 a_0_rep1_LC_5_10_3 (
            .in0(N__25001),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_0_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56272),
            .ce(N__56045),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIOKB71_11_LC_5_10_4 .C_ON=1'b0;
    defparam \ALU.r1_RNIOKB71_11_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIOKB71_11_LC_5_10_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.r1_RNIOKB71_11_LC_5_10_4  (
            .in0(N__24543),
            .in1(N__24998),
            .in2(N__25196),
            .in3(N__31060),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI3VN52_11_LC_5_10_5 .C_ON=1'b0;
    defparam \ALU.r5_RNI3VN52_11_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI3VN52_11_LC_5_10_5 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.r5_RNI3VN52_11_LC_5_10_5  (
            .in0(N__24734),
            .in1(N__26111),
            .in2(N__23674),
            .in3(N__30886),
            .lcout(\ALU.r5_RNI3VN52Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIU2G71_3_LC_5_10_6 .C_ON=1'b0;
    defparam \ALU.r2_RNIU2G71_3_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIU2G71_3_LC_5_10_6 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \ALU.r2_RNIU2G71_3_LC_5_10_6  (
            .in0(N__24795),
            .in1(N__24999),
            .in2(N__31084),
            .in3(N__23657),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIFJ8D2_3_LC_5_10_7 .C_ON=1'b0;
    defparam \ALU.r6_RNIFJ8D2_3_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIFJ8D2_3_LC_5_10_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNIFJ8D2_3_LC_5_10_7  (
            .in0(N__28046),
            .in1(N__39128),
            .in2(N__23629),
            .in3(N__30887),
            .lcout(\ALU.r6_RNIFJ8D2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIEV9A1_12_LC_5_11_0 .C_ON=1'b0;
    defparam \ALU.r1_RNIEV9A1_12_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIEV9A1_12_LC_5_11_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r1_RNIEV9A1_12_LC_5_11_0  (
            .in0(N__28375),
            .in1(N__30889),
            .in2(N__25163),
            .in3(N__25647),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIS3672_12_LC_5_11_1 .C_ON=1'b0;
    defparam \ALU.r5_RNIS3672_12_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIS3672_12_LC_5_11_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r5_RNIS3672_12_LC_5_11_1  (
            .in0(N__25563),
            .in1(N__26078),
            .in2(N__23626),
            .in3(N__25448),
            .lcout(\ALU.r5_RNIS3672Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIJ7I91_12_LC_5_11_2 .C_ON=1'b0;
    defparam \ALU.r2_RNIJ7I91_12_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIJ7I91_12_LC_5_11_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIJ7I91_12_LC_5_11_2  (
            .in0(N__25304),
            .in1(N__25564),
            .in2(N__23870),
            .in3(N__25648),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI5S672_12_LC_5_11_3 .C_ON=1'b0;
    defparam \ALU.r6_RNI5S672_12_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI5S672_12_LC_5_11_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNI5S672_12_LC_5_11_3  (
            .in0(N__25565),
            .in1(N__23621),
            .in2(N__23590),
            .in3(N__25253),
            .lcout(),
            .ltout(\ALU.r6_RNI5S672Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI9O1J4_12_LC_5_11_4 .C_ON=1'b0;
    defparam \ALU.r5_RNI9O1J4_12_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI9O1J4_12_LC_5_11_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r5_RNI9O1J4_12_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__29207),
            .in2(N__23587),
            .in3(N__23584),
            .lcout(\ALU.a_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_2_LC_5_11_5.C_ON=1'b0;
    defparam a_2_LC_5_11_5.SEQ_MODE=4'b1000;
    defparam a_2_LC_5_11_5.LUT_INIT=16'b0101101011110000;
    LogicCell40 a_2_LC_5_11_5 (
            .in0(N__25650),
            .in1(_gnd_net_),
            .in2(N__25596),
            .in3(N__32161),
            .lcout(aZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56277),
            .ce(N__56042),
            .sr(_gnd_net_));
    defparam a_2_rep2_LC_5_11_6.C_ON=1'b0;
    defparam a_2_rep2_LC_5_11_6.SEQ_MODE=4'b1000;
    defparam a_2_rep2_LC_5_11_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 a_2_rep2_LC_5_11_6 (
            .in0(N__32162),
            .in1(N__30890),
            .in2(_gnd_net_),
            .in3(N__25651),
            .lcout(a_2_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56277),
            .ce(N__56042),
            .sr(_gnd_net_));
    defparam a_0_LC_5_11_7.C_ON=1'b0;
    defparam a_0_LC_5_11_7.SEQ_MODE=4'b1000;
    defparam a_0_LC_5_11_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 a_0_LC_5_11_7 (
            .in0(N__25649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56277),
            .ce(N__56042),
            .sr(_gnd_net_));
    defparam \ALU.r2_12_LC_5_12_0 .C_ON=1'b0;
    defparam \ALU.r2_12_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_12_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_12_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28441),
            .lcout(r2_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56282),
            .ce(N__47686),
            .sr(_gnd_net_));
    defparam \ALU.r2_14_LC_5_12_1 .C_ON=1'b0;
    defparam \ALU.r2_14_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_14_LC_5_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r2_14_LC_5_12_1  (
            .in0(N__28310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r2_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56282),
            .ce(N__47686),
            .sr(_gnd_net_));
    defparam \ALU.r2_5_LC_5_12_2 .C_ON=1'b0;
    defparam \ALU.r2_5_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_5_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_5_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37210),
            .lcout(r2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56282),
            .ce(N__47686),
            .sr(_gnd_net_));
    defparam \ALU.r2_6_LC_5_12_3 .C_ON=1'b0;
    defparam \ALU.r2_6_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_6_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_6_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38873),
            .lcout(r2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56282),
            .ce(N__47686),
            .sr(_gnd_net_));
    defparam \ALU.r2_9_LC_5_12_4 .C_ON=1'b0;
    defparam \ALU.r2_9_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_9_LC_5_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_9_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34033),
            .lcout(r2_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56282),
            .ce(N__47686),
            .sr(_gnd_net_));
    defparam \ALU.r2_3_LC_5_12_5 .C_ON=1'b0;
    defparam \ALU.r2_3_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_3_LC_5_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r2_3_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50200),
            .lcout(r2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56282),
            .ce(N__47686),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_0_LC_5_13_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_0_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_0_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_15_s1_c_RNO_0_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__37519),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\ALU.r0_12_prm_8_15_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s1_c_LC_5_13_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_15_s1_c_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s1_c_LC_5_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_15_s1_c_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__36031),
            .in2(N__31201),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_15_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_15_s1_c_LC_5_13_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_15_s1_c_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_15_s1_c_LC_5_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_15_s1_c_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__35986),
            .in2(N__23836),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_15_s1 ),
            .carryout(\ALU.r0_12_prm_7_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_15_s1_c_LC_5_13_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_15_s1_c_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_15_s1_c_LC_5_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_15_s1_c_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__35949),
            .in2(N__23821),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_15_s1 ),
            .carryout(\ALU.r0_12_prm_6_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_15_s1_c_LC_5_13_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_15_s1_c_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_15_s1_c_LC_5_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_15_s1_c_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__35911),
            .in2(N__37540),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_15_s1 ),
            .carryout(\ALU.r0_12_prm_5_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_15_s1_c_LC_5_13_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_15_s1_c_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_15_s1_c_LC_5_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_15_s1_c_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__35881),
            .in2(N__23806),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_15_s1 ),
            .carryout(\ALU.r0_12_prm_4_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_15_s1_c_LC_5_13_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_15_s1_c_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_15_s1_c_LC_5_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_15_s1_c_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__55216),
            .in2(N__56413),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_15_s1 ),
            .carryout(\ALU.r0_12_prm_3_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_15_s1_c_LC_5_13_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_15_s1_c_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_15_s1_c_LC_5_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_15_s1_c_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__36259),
            .in2(N__31249),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_15_s1 ),
            .carryout(\ALU.r0_12_prm_2_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_15_s1_c_LC_5_14_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_15_s1_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_15_s1_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_15_s1_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__37297),
            .in2(N__37252),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\ALU.r0_12_s1_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_15_s0_c_RNI2DJ0GB2_LC_5_14_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_15_s0_c_RNI2DJ0GB2_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_15_s0_c_RNI2DJ0GB2_LC_5_14_1 .LUT_INIT=16'b1011111010000010;
    LogicCell40 \ALU.r0_12_prm_1_15_s0_c_RNI2DJ0GB2_LC_5_14_1  (
            .in0(N__36190),
            .in1(N__23791),
            .in2(N__27358),
            .in3(N__23779),
            .lcout(\ALU.r0_12_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_15_LC_5_14_2 .C_ON=1'b0;
    defparam \ALU.r0_15_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_15_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_15_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25968),
            .lcout(r0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56290),
            .ce(N__49717),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIHPP81_13_LC_5_15_0 .C_ON=1'b0;
    defparam \ALU.r1_RNIHPP81_13_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIHPP81_13_LC_5_15_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r1_RNIHPP81_13_LC_5_15_0  (
            .in0(N__26198),
            .in1(N__25598),
            .in2(N__25137),
            .in3(N__25680),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI10M52_13_LC_5_15_1 .C_ON=1'b0;
    defparam \ALU.r5_RNI10M52_13_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI10M52_13_LC_5_15_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r5_RNI10M52_13_LC_5_15_1  (
            .in0(N__26045),
            .in1(N__25412),
            .in2(N__23920),
            .in3(N__25602),
            .lcout(\ALU.r5_RNI10M52Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIL9I91_13_LC_5_15_2 .C_ON=1'b0;
    defparam \ALU.r2_RNIL9I91_13_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIL9I91_13_LC_5_15_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIL9I91_13_LC_5_15_2  (
            .in0(N__23916),
            .in1(N__25599),
            .in2(N__24102),
            .in3(N__25681),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI90772_13_LC_5_15_3 .C_ON=1'b0;
    defparam \ALU.r6_RNI90772_13_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI90772_13_LC_5_15_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNI90772_13_LC_5_15_3  (
            .in0(N__23981),
            .in1(N__24071),
            .in2(N__23887),
            .in3(N__25603),
            .lcout(),
            .ltout(\ALU.r6_RNI90772Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIIOHH4_13_LC_5_15_4 .C_ON=1'b0;
    defparam \ALU.r5_RNIIOHH4_13_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIIOHH4_13_LC_5_15_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r5_RNIIOHH4_13_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__29206),
            .in2(N__23884),
            .in3(N__23881),
            .lcout(\ALU.a_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIPV8A9_13_LC_5_15_6 .C_ON=1'b0;
    defparam \ALU.r5_RNIPV8A9_13_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIPV8A9_13_LC_5_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r5_RNIPV8A9_13_LC_5_15_6  (
            .in0(N__53900),
            .in1(N__47003),
            .in2(_gnd_net_),
            .in3(N__41445),
            .lcout(),
            .ltout(\ALU.r5_RNIPV8A9Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNILM5AE_15_LC_5_15_7 .C_ON=1'b0;
    defparam \ALU.r5_RNILM5AE_15_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNILM5AE_15_LC_5_15_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ALU.r5_RNILM5AE_15_LC_5_15_7  (
            .in0(N__53955),
            .in1(N__54383),
            .in2(N__23875),
            .in3(N__40142),
            .lcout(\ALU.r5_RNILM5AEZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r3_4_LC_5_16_2 .C_ON=1'b0;
    defparam \ALU.r3_4_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_4_LC_5_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_4_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39091),
            .lcout(r3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56299),
            .ce(N__47764),
            .sr(_gnd_net_));
    defparam \ALU.r3_12_LC_5_16_3 .C_ON=1'b0;
    defparam \ALU.r3_12_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_12_LC_5_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_12_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28423),
            .lcout(r3_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56299),
            .ce(N__47764),
            .sr(_gnd_net_));
    defparam \ALU.r3_5_LC_5_16_6 .C_ON=1'b0;
    defparam \ALU.r3_5_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_5_LC_5_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_5_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37216),
            .lcout(r3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56299),
            .ce(N__47764),
            .sr(_gnd_net_));
    defparam \ALU.r3_13_LC_5_16_7 .C_ON=1'b0;
    defparam \ALU.r3_13_LC_5_16_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r3_13_LC_5_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r3_13_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26242),
            .lcout(r3_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56299),
            .ce(N__47764),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_5_LC_5_17_2.C_ON=1'b0;
    defparam TXbuffer_RNO_6_5_LC_5_17_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_5_LC_5_17_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_6_5_LC_5_17_2 (
            .in0(N__30049),
            .in1(N__24079),
            .in2(N__24049),
            .in3(N__24036),
            .lcout(),
            .ltout(TXbuffer_RNO_6Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_5_LC_5_17_3.C_ON=1'b0;
    defparam TXbuffer_RNO_2_5_LC_5_17_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_5_LC_5_17_3.LUT_INIT=16'b0101010100011011;
    LogicCell40 TXbuffer_RNO_2_5_LC_5_17_3 (
            .in0(N__29669),
            .in1(N__23998),
            .in2(N__23992),
            .in3(N__49925),
            .lcout(TXbuffer_18_15_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_5_LC_5_17_4.C_ON=1'b0;
    defparam TXbuffer_RNO_1_5_LC_5_17_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_5_LC_5_17_4.LUT_INIT=16'b1010000011011101;
    LogicCell40 TXbuffer_RNO_1_5_LC_5_17_4 (
            .in0(N__30050),
            .in1(N__23989),
            .in2(N__23965),
            .in3(N__23932),
            .lcout(TXbuffer_RNO_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_5_LC_5_17_6.C_ON=1'b0;
    defparam TXbuffer_RNO_0_5_LC_5_17_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_5_LC_5_17_6.LUT_INIT=16'b1110001100100011;
    LogicCell40 TXbuffer_RNO_0_5_LC_5_17_6 (
            .in0(N__26049),
            .in1(N__23926),
            .in2(N__30080),
            .in3(N__25922),
            .lcout(TXbuffer_RNO_0Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_5_LC_5_18_3.C_ON=1'b0;
    defparam TXbuffer_RNO_3_5_LC_5_18_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_5_LC_5_18_3.LUT_INIT=16'b0000110100111101;
    LogicCell40 TXbuffer_RNO_3_5_LC_5_18_3 (
            .in0(N__37125),
            .in1(N__29987),
            .in2(N__30394),
            .in3(N__25138),
            .lcout(TXbuffer_18_10_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_4_c_RNO_LC_6_1_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_4_c_RNO_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_4_c_RNO_LC_6_1_0 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_4_c_RNO_LC_6_1_0  (
            .in0(N__40487),
            .in1(N__53212),
            .in2(N__53812),
            .in3(N__42788),
            .lcout(\ALU.r0_12_prm_6_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_6_s1_c_RNO_LC_6_1_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_6_s1_c_RNO_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_6_s1_c_RNO_LC_6_1_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_6_s1_c_RNO_LC_6_1_1  (
            .in0(N__54555),
            .in1(N__53590),
            .in2(N__53250),
            .in3(N__43283),
            .lcout(\ALU.r0_12_prm_4_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_81_LC_6_1_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_81_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_81_LC_6_1_2 .LUT_INIT=16'b0110000011000000;
    LogicCell40 \ALU.mult_madd_81_LC_6_1_2  (
            .in0(N__45500),
            .in1(N__24238),
            .in2(N__24165),
            .in3(N__43929),
            .lcout(\ALU.madd_46_0 ),
            .ltout(\ALU.madd_46_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_115_LC_6_1_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_115_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_115_LC_6_1_3 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ALU.mult_madd_115_LC_6_1_3  (
            .in0(N__24216),
            .in1(N__24204),
            .in2(N__24193),
            .in3(N__24190),
            .lcout(\ALU.madd_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_3_LC_6_1_4 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_3_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_3_LC_6_1_4 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a5_b_3_LC_6_1_4  (
            .in0(N__29078),
            .in1(N__29009),
            .in2(N__36753),
            .in3(N__44308),
            .lcout(\ALU.a5_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2BKQ8_6_LC_6_1_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI2BKQ8_6_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2BKQ8_6_LC_6_1_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r4_RNI2BKQ8_6_LC_6_1_5  (
            .in0(_gnd_net_),
            .in1(N__43648),
            .in2(_gnd_net_),
            .in3(N__43282),
            .lcout(\ALU.un14_log_0_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g2_0_LC_6_1_7 .C_ON=1'b0;
    defparam \ALU.mult_g2_0_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g2_0_LC_6_1_7 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_g2_0_LC_6_1_7  (
            .in0(N__44309),
            .in1(N__43281),
            .in2(N__45513),
            .in3(N__40486),
            .lcout(\ALU.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_7_LC_6_2_0 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_7_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_7_LC_6_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a0_b_7_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__48760),
            .in2(_gnd_net_),
            .in3(N__44765),
            .lcout(\ALU.a0_b_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_34_LC_6_2_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_34_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_34_LC_6_2_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \ALU.mult_madd_34_LC_6_2_1  (
            .in0(N__48762),
            .in1(N__26590),
            .in2(N__45257),
            .in3(N__26689),
            .lcout(\ALU.madd_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_33_LC_6_2_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_33_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_33_LC_6_2_2 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_33_LC_6_2_2  (
            .in0(N__24289),
            .in1(N__49288),
            .in2(N__24148),
            .in3(N__43896),
            .lcout(\ALU.madd_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_38_LC_6_2_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_38_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_38_LC_6_2_3 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \ALU.mult_madd_38_LC_6_2_3  (
            .in0(N__48763),
            .in1(N__26589),
            .in2(N__45258),
            .in3(N__26688),
            .lcout(\ALU.madd_38 ),
            .ltout(\ALU.madd_38_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_60_LC_6_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_60_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_60_LC_6_2_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_60_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__26643),
            .in2(N__24280),
            .in3(N__26661),
            .lcout(\ALU.madd_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_87_LC_6_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_87_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_87_LC_6_2_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_87_LC_6_2_5  (
            .in0(N__27163),
            .in1(N__27154),
            .in2(_gnd_net_),
            .in3(N__27139),
            .lcout(\ALU.madd_87 ),
            .ltout(\ALU.madd_87_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_120_LC_6_2_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_120_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_120_LC_6_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_120_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(N__26568),
            .in2(N__24277),
            .in3(N__26556),
            .lcout(\ALU.madd_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_6_LC_6_2_7 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_6_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_6_LC_6_2_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_a0_b_6_LC_6_2_7  (
            .in0(N__48761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43606),
            .lcout(\ALU.a0_b_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_92_LC_6_3_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_92_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_92_LC_6_3_0 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \ALU.mult_madd_92_LC_6_3_0  (
            .in0(N__24250),
            .in1(N__24265),
            .in2(N__27127),
            .in3(N__24271),
            .lcout(\ALU.madd_92 ),
            .ltout(\ALU.madd_92_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_7_LC_6_3_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_7_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_7_LC_6_3_1 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_axb_7_LC_6_3_1  (
            .in0(N__24352),
            .in1(N__26680),
            .in2(N__24274),
            .in3(N__26599),
            .lcout(\ALU.madd_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_78_0_LC_6_3_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_78_0_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_78_0_LC_6_3_2 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_78_0_LC_6_3_2  (
            .in0(N__48793),
            .in1(N__44790),
            .in2(N__43665),
            .in3(N__48510),
            .lcout(\ALU.madd_78_0 ),
            .ltout(\ALU.madd_78_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_88_LC_6_3_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_88_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_88_LC_6_3_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_88_LC_6_3_3  (
            .in0(N__24264),
            .in1(N__27123),
            .in2(N__24253),
            .in3(N__24249),
            .lcout(\ALU.madd_332 ),
            .ltout(\ALU.madd_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_6_l_ofx_LC_6_3_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_6_l_ofx_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_6_l_ofx_LC_6_3_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ALU.mult_madd_axb_6_l_ofx_LC_6_3_4  (
            .in0(N__26598),
            .in1(N__28892),
            .in2(N__24241),
            .in3(N__28876),
            .lcout(\ALU.madd_axb_6_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNII0MP4_0_LC_6_3_5 .C_ON=1'b0;
    defparam \ALU.r2_RNII0MP4_0_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNII0MP4_0_LC_6_3_5 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.r2_RNII0MP4_0_LC_6_3_5  (
            .in0(N__24376),
            .in1(N__28753),
            .in2(N__29208),
            .in3(N__27700),
            .lcout(\ALU.aZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI6N1R4_4_LC_6_3_6 .C_ON=1'b0;
    defparam \ALU.r4_RNI6N1R4_4_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI6N1R4_4_LC_6_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.r4_RNI6N1R4_4_LC_6_3_6  (
            .in0(N__32361),
            .in1(N__32453),
            .in2(_gnd_net_),
            .in3(N__29183),
            .lcout(\ALU.a_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_8_l_fx_LC_6_3_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_8_l_fx_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_8_l_fx_LC_6_3_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_axb_8_l_fx_LC_6_3_7  (
            .in0(N__26668),
            .in1(N__24358),
            .in2(N__27223),
            .in3(N__24351),
            .lcout(\ALU.madd_axb_8_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_0_ma_LC_6_4_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_0_ma_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_0_ma_LC_6_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_cry_0_ma_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__48792),
            .in2(_gnd_net_),
            .in3(N__46680),
            .lcout(\ALU.madd_cry_0_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_4_LC_6_4_1 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_4_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_4_LC_6_4_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.mult_a2_b_4_LC_6_4_1  (
            .in0(N__32675),
            .in1(N__40433),
            .in2(N__32173),
            .in3(N__32589),
            .lcout(\ALU.a2_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJQGK3_3_LC_6_4_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIJQGK3_3_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJQGK3_3_LC_6_4_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r4_RNIJQGK3_3_LC_6_4_2  (
            .in0(N__24329),
            .in1(N__24706),
            .in2(_gnd_net_),
            .in3(N__33030),
            .lcout(\ALU.b_3 ),
            .ltout(\ALU.b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2THO8_3_LC_6_4_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI2THO8_3_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2THO8_3_LC_6_4_3 .LUT_INIT=16'b1100001110100101;
    LogicCell40 \ALU.r4_RNI2THO8_3_LC_6_4_3  (
            .in0(N__31797),
            .in1(N__31902),
            .in2(N__24310),
            .in3(N__32129),
            .lcout(\ALU.un2_addsub_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI0TRV3_1_LC_6_4_4 .C_ON=1'b0;
    defparam \ALU.r2_RNI0TRV3_1_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI0TRV3_1_LC_6_4_4 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \ALU.r2_RNI0TRV3_1_LC_6_4_4  (
            .in0(N__29374),
            .in1(N__26731),
            .in2(N__28636),
            .in3(N__24705),
            .lcout(\ALU.b_1 ),
            .ltout(\ALU.b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a4_b_1_LC_6_4_5 .C_ON=1'b0;
    defparam \ALU.mult_a4_b_1_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a4_b_1_LC_6_4_5 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \ALU.mult_a4_b_1_LC_6_4_5  (
            .in0(N__32102),
            .in1(N__32460),
            .in2(N__24292),
            .in3(N__32362),
            .lcout(\ALU.a4_b_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIS1N55_3_LC_6_4_6 .C_ON=1'b0;
    defparam \ALU.r4_RNIS1N55_3_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIS1N55_3_LC_6_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIS1N55_3_LC_6_4_6  (
            .in0(N__27752),
            .in1(N__31901),
            .in2(_gnd_net_),
            .in3(N__31796),
            .lcout(\ALU.a_3 ),
            .ltout(\ALU.a_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g1_1_LC_6_4_7 .C_ON=1'b0;
    defparam \ALU.mult_g1_1_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g1_1_LC_6_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_g1_1_LC_6_4_7  (
            .in0(N__24462),
            .in1(N__40432),
            .in2(N__24433),
            .in3(N__45218),
            .lcout(\ALU.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNICA4F3_4_LC_6_5_0 .C_ON=1'b0;
    defparam \ALU.r4_RNICA4F3_4_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNICA4F3_4_LC_6_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.r4_RNICA4F3_4_LC_6_5_0  (
            .in0(N__33438),
            .in1(N__24701),
            .in2(_gnd_net_),
            .in3(N__24862),
            .lcout(\ALU.b_4 ),
            .ltout(\ALU.b_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_214_0_LC_6_5_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_214_0_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_214_0_LC_6_5_1 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_214_0_LC_6_5_1  (
            .in0(N__44248),
            .in1(N__45989),
            .in2(N__24418),
            .in3(N__44446),
            .lcout(\ALU.madd_214_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_373_0_LC_6_5_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_373_0_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_373_0_LC_6_5_2 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.mult_madd_373_0_LC_6_5_2  (
            .in0(N__40431),
            .in1(N__44250),
            .in2(N__51839),
            .in3(N__40986),
            .lcout(\ALU.madd_373_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIBIGK3_2_LC_6_5_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIBIGK3_2_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIBIGK3_2_LC_6_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIBIGK3_2_LC_6_5_3  (
            .in0(N__24700),
            .in1(N__29360),
            .in2(_gnd_net_),
            .in3(N__33347),
            .lcout(\ALU.b_2 ),
            .ltout(\ALU.b_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_11_LC_6_5_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_11_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_11_LC_6_5_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ALU.mult_g0_11_LC_6_5_4  (
            .in0(N__44449),
            .in1(N__46182),
            .in2(N__24406),
            .in3(N__46678),
            .lcout(\ALU.madd_134_0_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2QU6A_6_LC_6_5_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI2QU6A_6_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2QU6A_6_LC_6_5_5 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r4_RNI2QU6A_6_LC_6_5_5  (
            .in0(N__53421),
            .in1(N__43408),
            .in2(N__54215),
            .in3(N__44447),
            .lcout(\ALU.lshift_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIC5NE1_0_LC_6_5_6 .C_ON=1'b0;
    defparam \ALU.r4_RNIC5NE1_0_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIC5NE1_0_LC_6_5_6 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ALU.r4_RNIC5NE1_0_LC_6_5_6  (
            .in0(N__27685),
            .in1(N__33142),
            .in2(N__27637),
            .in3(N__33523),
            .lcout(\ALU.r4_RNIC5NE1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_172_0_LC_6_5_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_172_0_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_172_0_LC_6_5_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_172_0_LC_6_5_7  (
            .in0(N__44249),
            .in1(N__40430),
            .in2(N__43431),
            .in3(N__44448),
            .lcout(\ALU.madd_172_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_368_LC_6_6_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_368_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_368_LC_6_6_0 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_368_LC_6_6_0  (
            .in0(N__37886),
            .in1(N__27341),
            .in2(N__24496),
            .in3(N__47001),
            .lcout(\ALU.madd_368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a12_b_2_LC_6_6_1 .C_ON=1'b0;
    defparam \ALU.mult_a12_b_2_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a12_b_2_LC_6_6_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \ALU.mult_a12_b_2_LC_6_6_1  (
            .in0(N__41315),
            .in1(N__29359),
            .in2(N__32841),
            .in3(N__33349),
            .lcout(\ALU.a12_b_2 ),
            .ltout(\ALU.a12_b_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_372_LC_6_6_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_372_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_372_LC_6_6_2 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_372_LC_6_6_2  (
            .in0(N__37887),
            .in1(N__27342),
            .in2(N__24487),
            .in3(N__47002),
            .lcout(\ALU.madd_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a13_b_1_LC_6_6_3 .C_ON=1'b0;
    defparam \ALU.mult_a13_b_1_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a13_b_1_LC_6_6_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_a13_b_1_LC_6_6_3  (
            .in0(N__41548),
            .in1(N__46710),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.a13_b_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_6_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_6_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_368_0_LC_6_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_368_0_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_368_0_LC_6_6_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_368_0_LC_6_6_5  (
            .in0(N__41314),
            .in1(N__37885),
            .in2(N__47041),
            .in3(N__43862),
            .lcout(\ALU.madd_368_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g1_2_LC_6_6_6 .C_ON=1'b0;
    defparam \ALU.mult_g1_2_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g1_2_LC_6_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.mult_g1_2_LC_6_6_6  (
            .in0(N__29215),
            .in1(N__32447),
            .in2(_gnd_net_),
            .in3(N__32350),
            .lcout(\ALU.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_311_0_LC_6_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_311_0_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_311_0_LC_6_6_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_311_0_LC_6_6_7  (
            .in0(N__40931),
            .in1(N__37884),
            .in2(N__41565),
            .in3(N__43861),
            .lcout(\ALU.madd_311_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_2_rep2_LC_6_7_0.C_ON=1'b0;
    defparam b_2_rep2_LC_6_7_0.SEQ_MODE=4'b1000;
    defparam b_2_rep2_LC_6_7_0.LUT_INIT=16'b0111011110001000;
    LogicCell40 b_2_rep2_LC_6_7_0 (
            .in0(N__32816),
            .in1(N__25097),
            .in2(_gnd_net_),
            .in3(N__26827),
            .lcout(b_2_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam b_1_LC_6_7_1.C_ON=1'b0;
    defparam b_1_LC_6_7_1.SEQ_MODE=4'b1000;
    defparam b_1_LC_6_7_1.LUT_INIT=16'b0101010110101010;
    LogicCell40 b_1_LC_6_7_1 (
            .in0(N__25100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32815),
            .lcout(bZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam b_fast_2_LC_6_7_2.C_ON=1'b0;
    defparam b_fast_2_LC_6_7_2.SEQ_MODE=4'b1000;
    defparam b_fast_2_LC_6_7_2.LUT_INIT=16'b0111011110001000;
    LogicCell40 b_fast_2_LC_6_7_2 (
            .in0(N__32817),
            .in1(N__25098),
            .in2(_gnd_net_),
            .in3(N__33295),
            .lcout(b_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam b_fast_1_LC_6_7_3.C_ON=1'b0;
    defparam b_fast_1_LC_6_7_3.SEQ_MODE=4'b1000;
    defparam b_fast_1_LC_6_7_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 b_fast_1_LC_6_7_3 (
            .in0(N__25099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26874),
            .lcout(b_fastZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam b_1_rep1_LC_6_7_4.C_ON=1'b0;
    defparam b_1_rep1_LC_6_7_4.SEQ_MODE=4'b1000;
    defparam b_1_rep1_LC_6_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 b_1_rep1_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(N__25096),
            .in2(_gnd_net_),
            .in3(N__24699),
            .lcout(b_1_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam b_1_rep2_LC_6_7_5.C_ON=1'b0;
    defparam b_1_rep2_LC_6_7_5.SEQ_MODE=4'b1000;
    defparam b_1_rep2_LC_6_7_5.LUT_INIT=16'b0110011001100110;
    LogicCell40 b_1_rep2_LC_6_7_5 (
            .in0(N__25101),
            .in1(N__24581),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b_1_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam params_1_LC_6_7_6.C_ON=1'b0;
    defparam params_1_LC_6_7_6.SEQ_MODE=4'b1000;
    defparam params_1_LC_6_7_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 params_1_LC_6_7_6 (
            .in0(_gnd_net_),
            .in1(N__53356),
            .in2(_gnd_net_),
            .in3(N__54129),
            .lcout(paramsZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam params_0_LC_6_7_7.C_ON=1'b0;
    defparam params_0_LC_6_7_7.SEQ_MODE=4'b1000;
    defparam params_0_LC_6_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 params_0_LC_6_7_7 (
            .in0(N__53357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(paramsZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(N__56049),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIMQ992_3_LC_6_8_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIMQ992_3_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIMQ992_3_LC_6_8_0 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ALU.r4_RNIMQ992_3_LC_6_8_0  (
            .in0(N__33056),
            .in1(N__30924),
            .in2(N__33603),
            .in3(N__30583),
            .lcout(\ALU.r4_RNIMQ992Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_3_LC_6_8_1 .C_ON=1'b0;
    defparam \ALU.r4_3_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_3_LC_6_8_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r4_3_LC_6_8_1  (
            .in0(N__50192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56260),
            .ce(N__47809),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_3_LC_6_8_2.C_ON=1'b0;
    defparam TXbuffer_RNO_7_3_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_3_LC_6_8_2.LUT_INIT=16'b0000111100110101;
    LogicCell40 TXbuffer_RNO_7_3_LC_6_8_2 (
            .in0(N__35053),
            .in1(N__24547),
            .in2(N__30414),
            .in3(N__30064),
            .lcout(),
            .ltout(TXbuffer_18_3_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_3_LC_6_8_3.C_ON=1'b0;
    defparam TXbuffer_RNO_5_3_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_3_LC_6_8_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_5_3_LC_6_8_3 (
            .in0(N__30065),
            .in1(N__24735),
            .in2(N__24850),
            .in3(N__33057),
            .lcout(),
            .ltout(TXbuffer_RNO_5Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_3_LC_6_8_4.C_ON=1'b0;
    defparam TXbuffer_RNO_2_3_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_3_LC_6_8_4.LUT_INIT=16'b0100010101100111;
    LogicCell40 TXbuffer_RNO_2_3_LC_6_8_4 (
            .in0(N__29676),
            .in1(N__49968),
            .in2(N__24847),
            .in3(N__24742),
            .lcout(TXbuffer_18_15_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_3_LC_6_8_5.C_ON=1'b0;
    defparam TXbuffer_RNO_8_3_LC_6_8_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_3_LC_6_8_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_8_3_LC_6_8_5 (
            .in0(N__30062),
            .in1(N__24823),
            .in2(N__30395),
            .in3(N__24799),
            .lcout(),
            .ltout(TXbuffer_18_6_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_3_LC_6_8_6.C_ON=1'b0;
    defparam TXbuffer_RNO_6_3_LC_6_8_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_3_LC_6_8_6.LUT_INIT=16'b1100101000001111;
    LogicCell40 TXbuffer_RNO_6_3_LC_6_8_6 (
            .in0(N__24772),
            .in1(N__39139),
            .in2(N__24745),
            .in3(N__30063),
            .lcout(TXbuffer_RNO_6Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_11_LC_6_8_7 .C_ON=1'b0;
    defparam \ALU.r4_11_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_11_LC_6_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_11_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26183),
            .lcout(r4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56260),
            .ce(N__47809),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIUF9K8_1_10_LC_6_9_0 .C_ON=1'b0;
    defparam \ALU.r5_RNIUF9K8_1_10_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIUF9K8_1_10_LC_6_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r5_RNIUF9K8_1_10_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__52000),
            .in2(_gnd_net_),
            .in3(N__51652),
            .lcout(\ALU.r5_RNIUF9K8_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_2_rep1_LC_6_9_1.C_ON=1'b0;
    defparam a_2_rep1_LC_6_9_1.SEQ_MODE=4'b1000;
    defparam a_2_rep1_LC_6_9_1.LUT_INIT=16'b0101111110100000;
    LogicCell40 a_2_rep1_LC_6_9_1 (
            .in0(N__32043),
            .in1(_gnd_net_),
            .in2(N__25692),
            .in3(N__30568),
            .lcout(a_2_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam a_1_LC_6_9_2.C_ON=1'b0;
    defparam a_1_LC_6_9_2.SEQ_MODE=4'b1000;
    defparam a_1_LC_6_9_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 a_1_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(N__25682),
            .in2(_gnd_net_),
            .in3(N__32042),
            .lcout(aZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam a_fast_2_LC_6_9_3.C_ON=1'b0;
    defparam a_fast_2_LC_6_9_3.SEQ_MODE=4'b1000;
    defparam a_fast_2_LC_6_9_3.LUT_INIT=16'b0101111110100000;
    LogicCell40 a_fast_2_LC_6_9_3 (
            .in0(N__32044),
            .in1(_gnd_net_),
            .in2(N__25693),
            .in3(N__31066),
            .lcout(a_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam a_fast_1_LC_6_9_4.C_ON=1'b0;
    defparam a_fast_1_LC_6_9_4.SEQ_MODE=4'b1000;
    defparam a_fast_1_LC_6_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 a_fast_1_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__25684),
            .in2(_gnd_net_),
            .in3(N__27734),
            .lcout(a_fastZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam a_1_rep1_LC_6_9_5.C_ON=1'b0;
    defparam a_1_rep1_LC_6_9_5.SEQ_MODE=4'b1000;
    defparam a_1_rep1_LC_6_9_5.LUT_INIT=16'b0110011001100110;
    LogicCell40 a_1_rep1_LC_6_9_5 (
            .in0(N__25691),
            .in1(N__29160),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_1_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam a_1_rep2_LC_6_9_6.C_ON=1'b0;
    defparam a_1_rep2_LC_6_9_6.SEQ_MODE=4'b1000;
    defparam a_1_rep2_LC_6_9_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 a_1_rep2_LC_6_9_6 (
            .in0(_gnd_net_),
            .in1(N__25683),
            .in2(_gnd_net_),
            .in3(N__36563),
            .lcout(a_1_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam b_2_rep1_LC_6_9_7.C_ON=1'b0;
    defparam b_2_rep1_LC_6_9_7.SEQ_MODE=4'b1000;
    defparam b_2_rep1_LC_6_9_7.LUT_INIT=16'b0110011010101010;
    LogicCell40 b_2_rep1_LC_6_9_7 (
            .in0(N__33113),
            .in1(N__25102),
            .in2(_gnd_net_),
            .in3(N__32834),
            .lcout(b_2_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56265),
            .ce(N__56046),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIHDA71_4_LC_6_10_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIHDA71_4_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIHDA71_4_LC_6_10_0 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.r2_RNIHDA71_4_LC_6_10_0  (
            .in0(N__25011),
            .in1(N__30553),
            .in2(N__25287),
            .in3(N__24953),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI403D2_4_LC_6_10_1 .C_ON=1'b0;
    defparam \ALU.r6_RNI403D2_4_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI403D2_4_LC_6_10_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.r6_RNI403D2_4_LC_6_10_1  (
            .in0(N__39000),
            .in1(N__28017),
            .in2(N__24961),
            .in3(N__30925),
            .lcout(\ALU.r6_RNI403D2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_4_LC_6_10_2 .C_ON=1'b0;
    defparam \ALU.r2_4_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_4_LC_6_10_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r2_4_LC_6_10_2  (
            .in0(N__39090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56269),
            .ce(N__47664),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIJRKU_4_LC_6_10_3 .C_ON=1'b0;
    defparam \ALU.r2_RNIJRKU_4_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIJRKU_4_LC_6_10_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNIJRKU_4_LC_6_10_3  (
            .in0(N__25275),
            .in1(N__33111),
            .in2(N__24957),
            .in3(N__24925),
            .lcout(),
            .ltout(\ALU.b_6_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNI7L2O1_4_LC_6_10_4 .C_ON=1'b0;
    defparam \ALU.r6_RNI7L2O1_4_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNI7L2O1_4_LC_6_10_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r6_RNI7L2O1_4_LC_6_10_4  (
            .in0(N__28016),
            .in1(N__38999),
            .in2(N__24865),
            .in3(N__26828),
            .lcout(\ALU.r6_RNI7L2O1Z0Z_4 ),
            .ltout(\ALU.r6_RNI7L2O1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIE2CL3_4_LC_6_10_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIE2CL3_4_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIE2CL3_4_LC_6_10_5 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \ALU.r4_RNIE2CL3_4_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__32830),
            .in2(N__25321),
            .in3(N__33439),
            .lcout(\ALU.b_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_8_4_LC_6_10_6.C_ON=1'b0;
    defparam TXbuffer_RNO_8_4_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_8_4_LC_6_10_6.LUT_INIT=16'b0001000110101111;
    LogicCell40 TXbuffer_RNO_8_4_LC_6_10_6 (
            .in0(N__30046),
            .in1(N__25318),
            .in2(N__25288),
            .in3(N__30309),
            .lcout(),
            .ltout(TXbuffer_18_6_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_6_4_LC_6_10_7.C_ON=1'b0;
    defparam TXbuffer_RNO_6_4_LC_6_10_7.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_6_4_LC_6_10_7.LUT_INIT=16'b1000111110000011;
    LogicCell40 TXbuffer_RNO_6_4_LC_6_10_7 (
            .in0(N__39001),
            .in1(N__30047),
            .in2(N__25264),
            .in3(N__25261),
            .lcout(TXbuffer_RNO_6Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_10_LC_6_11_0 .C_ON=1'b0;
    defparam \ALU.r1_10_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_10_LC_6_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_10_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28160),
            .lcout(r1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r1_11_LC_6_11_1 .C_ON=1'b0;
    defparam \ALU.r1_11_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_11_LC_6_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_11_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26184),
            .lcout(r1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r1_12_LC_6_11_2 .C_ON=1'b0;
    defparam \ALU.r1_12_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_12_LC_6_11_2 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \ALU.r1_12_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28447),
            .in3(_gnd_net_),
            .lcout(r1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r1_13_LC_6_11_3 .C_ON=1'b0;
    defparam \ALU.r1_13_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_13_LC_6_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_13_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26280),
            .lcout(r1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r1_15_LC_6_11_4 .C_ON=1'b0;
    defparam \ALU.r1_15_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_15_LC_6_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_15_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25989),
            .lcout(r1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r1_8_LC_6_11_5 .C_ON=1'b0;
    defparam \ALU.r1_8_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_8_LC_6_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_8_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39523),
            .lcout(r1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r1_9_LC_6_11_6 .C_ON=1'b0;
    defparam \ALU.r1_9_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_9_LC_6_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_9_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34031),
            .lcout(r1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56273),
            .ce(N__47560),
            .sr(_gnd_net_));
    defparam \ALU.r4_0_LC_6_12_0 .C_ON=1'b0;
    defparam \ALU.r4_0_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_0_LC_6_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_0_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35000),
            .lcout(r4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_10_LC_6_12_1 .C_ON=1'b0;
    defparam \ALU.r4_10_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_10_LC_6_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_10_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28159),
            .lcout(r4_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_12_LC_6_12_2 .C_ON=1'b0;
    defparam \ALU.r4_12_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_12_LC_6_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_12_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28442),
            .lcout(r4_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_13_LC_6_12_3 .C_ON=1'b0;
    defparam \ALU.r4_13_LC_6_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_13_LC_6_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_13_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26278),
            .lcout(r4_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_14_LC_6_12_4 .C_ON=1'b0;
    defparam \ALU.r4_14_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_14_LC_6_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_14_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28308),
            .lcout(r4_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_15_LC_6_12_5 .C_ON=1'b0;
    defparam \ALU.r4_15_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_15_LC_6_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_15_LC_6_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25988),
            .lcout(r4_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_5_LC_6_12_6 .C_ON=1'b0;
    defparam \ALU.r4_5_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_5_LC_6_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r4_5_LC_6_12_6  (
            .in0(N__37189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r4_6_LC_6_12_7 .C_ON=1'b0;
    defparam \ALU.r4_6_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_6_LC_6_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_6_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38872),
            .lcout(r4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56278),
            .ce(N__47802),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNIJRP81_14_LC_6_13_0 .C_ON=1'b0;
    defparam \ALU.r1_RNIJRP81_14_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNIJRP81_14_LC_6_13_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r1_RNIJRP81_14_LC_6_13_0  (
            .in0(N__25706),
            .in1(N__25575),
            .in2(N__28238),
            .in3(N__25662),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI54M52_14_LC_6_13_1 .C_ON=1'b0;
    defparam \ALU.r5_RNI54M52_14_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI54M52_14_LC_6_13_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r5_RNI54M52_14_LC_6_13_1  (
            .in0(N__25576),
            .in1(N__26021),
            .in2(N__25891),
            .in3(N__25880),
            .lcout(\ALU.r5_RNI54M52Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINBI91_14_LC_6_13_2 .C_ON=1'b0;
    defparam \ALU.r2_RNINBI91_14_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINBI91_14_LC_6_13_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r2_RNINBI91_14_LC_6_13_2  (
            .in0(N__25844),
            .in1(N__25578),
            .in2(N__25831),
            .in3(N__25664),
            .lcout(),
            .ltout(\ALU.a_6_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNID4772_14_LC_6_13_3 .C_ON=1'b0;
    defparam \ALU.r6_RNID4772_14_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNID4772_14_LC_6_13_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r6_RNID4772_14_LC_6_13_3  (
            .in0(N__25580),
            .in1(N__25797),
            .in2(N__25768),
            .in3(N__25765),
            .lcout(),
            .ltout(\ALU.r6_RNID4772Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIR0IH4_14_LC_6_13_4 .C_ON=1'b0;
    defparam \ALU.r5_RNIR0IH4_14_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIR0IH4_14_LC_6_13_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r5_RNIR0IH4_14_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(N__36664),
            .in2(N__25735),
            .in3(N__25732),
            .lcout(\ALU.a_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_14_LC_6_13_5 .C_ON=1'b0;
    defparam \ALU.r0_14_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_14_LC_6_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r0_14_LC_6_13_5  (
            .in0(N__28295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56283),
            .ce(N__49730),
            .sr(_gnd_net_));
    defparam \ALU.r1_RNILTP81_15_LC_6_13_6 .C_ON=1'b0;
    defparam \ALU.r1_RNILTP81_15_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r1_RNILTP81_15_LC_6_13_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r1_RNILTP81_15_LC_6_13_6  (
            .in0(N__30107),
            .in1(N__25577),
            .in2(N__30479),
            .in3(N__25663),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI98M52_15_LC_6_13_7 .C_ON=1'b0;
    defparam \ALU.r5_RNI98M52_15_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI98M52_15_LC_6_13_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r5_RNI98M52_15_LC_6_13_7  (
            .in0(N__25579),
            .in1(N__30434),
            .in2(N__25495),
            .in3(N__29708),
            .lcout(\ALU.r5_RNI98M52Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_0_LC_6_14_0 .C_ON=1'b0;
    defparam \ALU.r5_0_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_0_LC_6_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_0_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35009),
            .lcout(r5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_10_LC_6_14_1 .C_ON=1'b0;
    defparam \ALU.r5_10_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_10_LC_6_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_10_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28176),
            .lcout(r5_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_11_LC_6_14_2 .C_ON=1'b0;
    defparam \ALU.r5_11_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_11_LC_6_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_11_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26185),
            .lcout(r5_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_12_LC_6_14_3 .C_ON=1'b0;
    defparam \ALU.r5_12_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_12_LC_6_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_12_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28427),
            .lcout(r5_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_13_LC_6_14_4 .C_ON=1'b0;
    defparam \ALU.r5_13_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_13_LC_6_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_13_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26261),
            .lcout(r5_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_14_LC_6_14_5 .C_ON=1'b0;
    defparam \ALU.r5_14_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_14_LC_6_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_14_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28294),
            .lcout(r5_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_15_LC_6_14_6 .C_ON=1'b0;
    defparam \ALU.r5_15_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_15_LC_6_14_6 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \ALU.r5_15_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25986),
            .in3(_gnd_net_),
            .lcout(r5_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r5_5_LC_6_14_7 .C_ON=1'b0;
    defparam \ALU.r5_5_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_5_LC_6_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_5_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37208),
            .lcout(r5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56286),
            .ce(N__45805),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_0_LC_6_15_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_0_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_0_LC_6_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_13_s0_c_RNO_0_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__39658),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\ALU.r0_12_prm_8_13_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s0_c_LC_6_15_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_13_s0_c_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s0_c_LC_6_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_13_s0_c_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__36160),
            .in2(N__35713),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_13_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_13_s0_c_LC_6_15_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_13_s0_c_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_13_s0_c_LC_6_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_13_s0_c_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__31476),
            .in2(N__26335),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_13_s0 ),
            .carryout(\ALU.r0_12_prm_7_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_13_s0_c_LC_6_15_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_13_s0_c_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_13_s0_c_LC_6_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_13_s0_c_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__31432),
            .in2(N__26350),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_13_s0 ),
            .carryout(\ALU.r0_12_prm_6_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_13_s0_c_LC_6_15_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_13_s0_c_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_13_s0_c_LC_6_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_13_s0_c_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__26359),
            .in2(N__31398),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_13_s0 ),
            .carryout(\ALU.r0_12_prm_5_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_13_s0_c_inv_LC_6_15_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_13_s0_c_inv_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_13_s0_c_inv_LC_6_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_13_s0_c_inv_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(N__31359),
            .in2(N__26371),
            .in3(N__41468),
            .lcout(\ALU.a_i_13 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_13_s0 ),
            .carryout(\ALU.r0_12_prm_4_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_13_s0_c_inv_LC_6_15_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_13_s0_c_inv_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_13_s0_c_inv_LC_6_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_3_13_s0_c_inv_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(N__26290),
            .in2(_gnd_net_),
            .in3(N__55220),
            .lcout(\ALU.r0_12_prm_3_13_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_13_s0 ),
            .carryout(\ALU.r0_12_prm_3_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_13_s0_c_LC_6_15_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_13_s0_c_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_13_s0_c_LC_6_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_13_s0_c_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(N__34597),
            .in2(N__31234),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_13_s0 ),
            .carryout(\ALU.r0_12_prm_2_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_13_s0_c_LC_6_16_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_13_s0_c_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_13_s0_c_LC_6_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_13_s0_c_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__35302),
            .in2(N__34624),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_16_0_),
            .carryout(\ALU.r0_12_s0_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_13_s0_c_RNIMPTBGM2_LC_6_16_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_13_s0_c_RNIMPTBGM2_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_13_s0_c_RNIMPTBGM2_LC_6_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r0_12_prm_1_13_s0_c_RNIMPTBGM2_LC_6_16_1  (
            .in0(N__27412),
            .in1(N__31513),
            .in2(_gnd_net_),
            .in3(N__26284),
            .lcout(\ALU.r0_12_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_13_LC_6_16_2 .C_ON=1'b0;
    defparam \ALU.r0_13_LC_6_16_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_13_LC_6_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_13_LC_6_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26241),
            .lcout(r0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56294),
            .ce(N__49726),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_13_s1_c_RNO_LC_6_17_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_13_s1_c_RNO_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_13_s1_c_RNO_LC_6_17_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r0_12_prm_4_13_s1_c_RNO_LC_6_17_0  (
            .in0(N__41500),
            .in1(N__54592),
            .in2(N__54061),
            .in3(N__52982),
            .lcout(\ALU.r0_12_prm_4_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIK81F5_13_LC_6_17_1 .C_ON=1'b0;
    defparam \ALU.r5_RNIK81F5_13_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIK81F5_13_LC_6_17_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r5_RNIK81F5_13_LC_6_17_1  (
            .in0(N__54028),
            .in1(N__54594),
            .in2(N__53163),
            .in3(N__41504),
            .lcout(\ALU.r5_RNIK81F5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_13_s0_c_RNO_LC_6_17_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_13_s0_c_RNO_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_13_s0_c_RNO_LC_6_17_2 .LUT_INIT=16'b0110100110100101;
    LogicCell40 \ALU.r0_12_prm_5_13_s0_c_RNO_LC_6_17_2  (
            .in0(N__41503),
            .in1(N__52985),
            .in2(N__35427),
            .in3(N__54593),
            .lcout(\ALU.r0_12_prm_5_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_12_s1_c_RNO_LC_6_17_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_12_s1_c_RNO_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_12_s1_c_RNO_LC_6_17_3 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_12_s1_c_RNO_LC_6_17_3  (
            .in0(N__54590),
            .in1(N__39859),
            .in2(N__53160),
            .in3(N__41316),
            .lcout(\ALU.r0_12_prm_5_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_13_s0_c_RNO_LC_6_17_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_13_s0_c_RNO_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_13_s0_c_RNO_LC_6_17_4 .LUT_INIT=16'b1100100100000101;
    LogicCell40 \ALU.r0_12_prm_6_13_s0_c_RNO_LC_6_17_4  (
            .in0(N__41502),
            .in1(N__52983),
            .in2(N__35426),
            .in3(N__54027),
            .lcout(\ALU.r0_12_prm_6_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_13_s1_c_RNO_LC_6_17_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_13_s1_c_RNO_LC_6_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_13_s1_c_RNO_LC_6_17_5 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_13_s1_c_RNO_LC_6_17_5  (
            .in0(N__54026),
            .in1(N__35410),
            .in2(N__53161),
            .in3(N__41498),
            .lcout(\ALU.r0_12_prm_6_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_13_s0_c_RNO_LC_6_17_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_13_s0_c_RNO_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_13_s0_c_RNO_LC_6_17_6 .LUT_INIT=16'b1010000001011111;
    LogicCell40 \ALU.r0_12_prm_7_13_s0_c_RNO_LC_6_17_6  (
            .in0(N__41501),
            .in1(_gnd_net_),
            .in2(N__35425),
            .in3(N__52984),
            .lcout(\ALU.r0_12_prm_7_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_13_s1_c_RNO_LC_6_17_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_13_s1_c_RNO_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_13_s1_c_RNO_LC_6_17_7 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_13_s1_c_RNO_LC_6_17_7  (
            .in0(N__54591),
            .in1(N__35411),
            .in2(N__53162),
            .in3(N__41499),
            .lcout(\ALU.r0_12_prm_5_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_9_l_ofx_LC_7_1_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_9_l_ofx_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_9_l_ofx_LC_7_1_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_axb_9_l_ofx_LC_7_1_0  (
            .in0(N__26545),
            .in1(N__26533),
            .in2(N__26323),
            .in3(N__26305),
            .lcout(\ALU.madd_axb_9_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_9_ma_LC_7_1_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_9_ma_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_9_ma_LC_7_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_cry_9_ma_LC_7_1_1  (
            .in0(_gnd_net_),
            .in1(N__26544),
            .in2(_gnd_net_),
            .in3(N__26532),
            .lcout(\ALU.madd_cry_9_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_124_LC_7_1_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_124_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_124_LC_7_1_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_124_LC_7_1_2  (
            .in0(N__26581),
            .in1(N__26575),
            .in2(_gnd_net_),
            .in3(N__26557),
            .lcout(\ALU.madd_124 ),
            .ltout(\ALU.madd_124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_165_LC_7_1_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_165_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_165_LC_7_1_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_165_LC_7_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26536),
            .in3(N__26531),
            .lcout(\ALU.madd_165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_0_s1_c_RNO_LC_7_1_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_0_s1_c_RNO_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_0_s1_c_RNO_LC_7_1_4 .LUT_INIT=16'b1001110001100011;
    LogicCell40 \ALU.r0_12_prm_1_0_s1_c_RNO_LC_7_1_4  (
            .in0(N__53946),
            .in1(N__48910),
            .in2(N__55955),
            .in3(N__38007),
            .lcout(\ALU.r0_12_prm_1_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a6_b_6_LC_7_1_5 .C_ON=1'b0;
    defparam \ALU.mult_a6_b_6_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a6_b_6_LC_7_1_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.mult_a6_b_6_LC_7_1_5  (
            .in0(N__26514),
            .in1(N__43607),
            .in2(N__32261),
            .in3(N__26447),
            .lcout(\ALU.a6_b_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_0_s0_c_RNO_LC_7_1_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_0_s0_c_RNO_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_0_s0_c_RNO_LC_7_1_6 .LUT_INIT=16'b1001110001100011;
    LogicCell40 \ALU.r0_12_prm_1_0_s0_c_RNO_LC_7_1_6  (
            .in0(N__53948),
            .in1(N__48912),
            .in2(N__55956),
            .in3(N__38008),
            .lcout(\ALU.r0_12_prm_1_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIKG5N5_0_LC_7_1_7 .C_ON=1'b0;
    defparam \ALU.r2_RNIKG5N5_0_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIKG5N5_0_LC_7_1_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r2_RNIKG5N5_0_LC_7_1_7  (
            .in0(N__48911),
            .in1(N__53947),
            .in2(N__53257),
            .in3(N__54556),
            .lcout(\ALU.r2_RNIKG5N5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_29_0_LC_7_2_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_29_0_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_29_0_LC_7_2_0 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_29_0_LC_7_2_0  (
            .in0(N__42723),
            .in1(N__37967),
            .in2(N__45496),
            .in3(N__46748),
            .lcout(\ALU.madd_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_14_LC_7_2_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_14_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_14_LC_7_2_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_14_LC_7_2_1  (
            .in0(N__37969),
            .in1(N__40731),
            .in2(N__26383),
            .in3(N__42725),
            .lcout(\ALU.madd_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_1_LC_7_2_2 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_1_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_1_LC_7_2_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a3_b_1_LC_7_2_2  (
            .in0(N__31935),
            .in1(N__31828),
            .in2(N__36771),
            .in3(N__46747),
            .lcout(\ALU.a3_b_1 ),
            .ltout(\ALU.a3_b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_18_LC_7_2_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_18_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_18_LC_7_2_3 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_18_LC_7_2_3  (
            .in0(N__37968),
            .in1(N__40730),
            .in2(N__26374),
            .in3(N__42724),
            .lcout(\ALU.madd_18 ),
            .ltout(\ALU.madd_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_43_LC_7_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_43_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_43_LC_7_2_4 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \ALU.mult_madd_43_LC_7_2_4  (
            .in0(N__29562),
            .in1(N__28593),
            .in2(N__26695),
            .in3(N__28617),
            .lcout(\ALU.madd_43 ),
            .ltout(\ALU.madd_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_5_l_fx_LC_7_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_5_l_fx_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_5_l_fx_LC_7_2_5 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \ALU.mult_madd_axb_5_l_fx_LC_7_2_5  (
            .in0(N__26725),
            .in1(N__26628),
            .in2(N__26692),
            .in3(N__29266),
            .lcout(\ALU.madd_axb_5_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_3_LC_7_2_6 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_3_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_3_LC_7_2_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a2_b_3_LC_7_2_6  (
            .in0(N__32685),
            .in1(N__32593),
            .in2(N__36770),
            .in3(N__44313),
            .lcout(\ALU.a2_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_94_LC_7_2_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_94_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_94_LC_7_2_7 .LUT_INIT=16'b1110100000000000;
    LogicCell40 \ALU.mult_madd_94_LC_7_2_7  (
            .in0(N__26724),
            .in1(N__26611),
            .in2(N__26632),
            .in3(N__26679),
            .lcout(\ALU.madd_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_56_LC_7_3_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_56_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_56_LC_7_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_56_LC_7_3_0  (
            .in0(N__26662),
            .in1(N__26650),
            .in2(_gnd_net_),
            .in3(N__26644),
            .lcout(\ALU.madd_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_51_LC_7_3_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_51_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_51_LC_7_3_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_51_LC_7_3_1  (
            .in0(N__44276),
            .in1(N__26902),
            .in2(N__26893),
            .in3(N__49254),
            .lcout(\ALU.madd_51 ),
            .ltout(\ALU.madd_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_65_LC_7_3_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_65_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_65_LC_7_3_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_65_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__26718),
            .in2(N__26614),
            .in3(N__26610),
            .lcout(\ALU.madd_331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a1_b_4_LC_7_3_3 .C_ON=1'b0;
    defparam \ALU.mult_a1_b_4_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a1_b_4_LC_7_3_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a1_b_4_LC_7_3_3  (
            .in0(N__31647),
            .in1(N__31738),
            .in2(N__36765),
            .in3(N__40531),
            .lcout(\ALU.a1_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_73_0_LC_7_3_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_73_0_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_73_0_LC_7_3_4 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_73_0_LC_7_3_4  (
            .in0(N__40532),
            .in1(N__49238),
            .in2(N__42787),
            .in3(N__44274),
            .lcout(),
            .ltout(\ALU.madd_73_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_73_LC_7_3_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_73_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_73_LC_7_3_5 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ALU.mult_madd_73_LC_7_3_5  (
            .in0(N__45190),
            .in1(_gnd_net_),
            .in2(N__26905),
            .in3(N__48361),
            .lcout(\ALU.madd_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a1_b_5_LC_7_3_6 .C_ON=1'b0;
    defparam \ALU.mult_a1_b_5_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a1_b_5_LC_7_3_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ALU.mult_a1_b_5_LC_7_3_6  (
            .in0(N__31739),
            .in1(N__45189),
            .in2(N__32185),
            .in3(N__31648),
            .lcout(\ALU.a1_b_5 ),
            .ltout(\ALU.a1_b_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_55_LC_7_3_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_55_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_55_LC_7_3_7 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_55_LC_7_3_7  (
            .in0(N__44275),
            .in1(N__26889),
            .in2(N__26878),
            .in3(N__49253),
            .lcout(\ALU.madd_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_2_LC_7_4_0 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_2_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_2_LC_7_4_0 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \ALU.mult_a2_b_2_LC_7_4_0  (
            .in0(N__43818),
            .in1(N__36734),
            .in2(N__32591),
            .in3(N__32677),
            .lcout(\ALU.a2_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIMTDQ_1_LC_7_4_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIMTDQ_1_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIMTDQ_1_LC_7_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.r4_RNIMTDQ_1_LC_7_4_1  (
            .in0(N__34368),
            .in1(N__33202),
            .in2(_gnd_net_),
            .in3(N__33663),
            .lcout(),
            .ltout(\ALU.r4_RNIMTDQZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI73OM1_1_LC_7_4_2 .C_ON=1'b0;
    defparam \ALU.r0_RNI73OM1_1_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI73OM1_1_LC_7_4_2 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \ALU.r0_RNI73OM1_1_LC_7_4_2  (
            .in0(N__26875),
            .in1(N__26833),
            .in2(N__26734),
            .in3(N__32935),
            .lcout(\ALU.b_7_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_46_LC_7_4_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_46_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_46_LC_7_4_3 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_46_LC_7_4_3  (
            .in0(N__42727),
            .in1(N__35116),
            .in2(N__26707),
            .in3(N__43820),
            .lcout(\ALU.madd_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a5_b_1_LC_7_4_4 .C_ON=1'b0;
    defparam \ALU.mult_a5_b_1_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a5_b_1_LC_7_4_4 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \ALU.mult_a5_b_1_LC_7_4_4  (
            .in0(N__29080),
            .in1(N__32106),
            .in2(N__29014),
            .in3(N__46679),
            .lcout(\ALU.a5_b_1 ),
            .ltout(\ALU.a5_b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_50_LC_7_4_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_50_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_50_LC_7_4_5 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_50_LC_7_4_5  (
            .in0(N__42726),
            .in1(N__35115),
            .in2(N__27166),
            .in3(N__43819),
            .lcout(\ALU.madd_50 ),
            .ltout(\ALU.madd_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_83_LC_7_4_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_83_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_83_LC_7_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_83_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(N__27153),
            .in2(N__27142),
            .in3(N__27138),
            .lcout(\ALU.madd_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIHCHO8_2_LC_7_4_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIHCHO8_2_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIHCHO8_2_LC_7_4_7 .LUT_INIT=16'b1010110001010011;
    LogicCell40 \ALU.r4_RNIHCHO8_2_LC_7_4_7  (
            .in0(N__32676),
            .in1(N__32579),
            .in2(N__32174),
            .in3(N__43817),
            .lcout(\ALU.un2_addsub_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_2_LC_7_5_0.C_ON=1'b0;
    defparam TXbuffer_2_LC_7_5_0.SEQ_MODE=4'b1000;
    defparam TXbuffer_2_LC_7_5_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 TXbuffer_2_LC_7_5_0 (
            .in0(N__27115),
            .in1(N__27895),
            .in2(N__49978),
            .in3(N__27097),
            .lcout(TXbufferZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56253),
            .ce(N__56051),
            .sr(_gnd_net_));
    defparam clkdiv_RNIQAHO1_0_LC_7_5_3.C_ON=1'b0;
    defparam clkdiv_RNIQAHO1_0_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam clkdiv_RNIQAHO1_0_LC_7_5_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 clkdiv_RNIQAHO1_0_LC_7_5_3 (
            .in0(N__27082),
            .in1(N__27055),
            .in2(N__27031),
            .in3(N__26989),
            .lcout(params5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_3_LC_7_5_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_3_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_3_LC_7_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_axb_3_LC_7_5_4  (
            .in0(N__26937),
            .in1(N__28524),
            .in2(_gnd_net_),
            .in3(N__29331),
            .lcout(\ALU.madd_axb_3 ),
            .ltout(\ALU.madd_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_3_s_LC_7_5_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_3_s_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_3_s_LC_7_5_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_cry_3_s_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26941),
            .in3(N__38544),
            .lcout(\ALU.mult_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_28_LC_7_5_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_28_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_28_LC_7_5_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_28_LC_7_5_6  (
            .in0(N__26938),
            .in1(N__28525),
            .in2(_gnd_net_),
            .in3(N__29332),
            .lcout(\ALU.madd_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_0_0_c_LC_7_6_0 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_0_0_c_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_0_0_c_LC_7_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_madd_cry_0_0_c_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__26926),
            .in2(N__26917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\ALU.madd_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_0_THRU_LUT4_0_LC_7_6_1 .C_ON=1'b1;
    defparam \ALU.madd_cry_0_THRU_LUT4_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_0_THRU_LUT4_0_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_0_THRU_LUT4_0_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__42898),
            .in2(_gnd_net_),
            .in3(N__27268),
            .lcout(\ALU.madd_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_0 ),
            .carryout(\ALU.madd_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_1_THRU_LUT4_0_LC_7_6_2 .C_ON=1'b1;
    defparam \ALU.madd_cry_1_THRU_LUT4_0_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_1_THRU_LUT4_0_LC_7_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_1_THRU_LUT4_0_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__50052),
            .in2(_gnd_net_),
            .in3(N__27265),
            .lcout(\ALU.madd_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_1 ),
            .carryout(\ALU.madd_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_2_THRU_LUT4_0_LC_7_6_3 .C_ON=1'b1;
    defparam \ALU.madd_cry_2_THRU_LUT4_0_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_2_THRU_LUT4_0_LC_7_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_2_THRU_LUT4_0_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__38559),
            .in2(_gnd_net_),
            .in3(N__27262),
            .lcout(\ALU.madd_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_2 ),
            .carryout(\ALU.madd_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_4_s_LC_7_6_4 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_4_s_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_4_s_LC_7_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_4_s_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__28563),
            .in2(N__28552),
            .in3(N__27259),
            .lcout(\ALU.mult_5 ),
            .ltout(),
            .carryin(\ALU.madd_cry_3 ),
            .carryout(\ALU.madd_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_5_s_LC_7_6_5 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_5_s_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_5_s_LC_7_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_5_s_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__29262),
            .in2(N__27256),
            .in3(N__27244),
            .lcout(\ALU.mult_6 ),
            .ltout(),
            .carryin(\ALU.madd_cry_4 ),
            .carryout(\ALU.madd_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_6_0_s_LC_7_6_6 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_6_0_s_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_6_0_s_LC_7_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_6_0_s_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__27241),
            .in2(N__28855),
            .in3(N__27229),
            .lcout(\ALU.mult_7 ),
            .ltout(),
            .carryin(\ALU.madd_cry_5 ),
            .carryout(\ALU.madd_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_6_THRU_LUT4_0_LC_7_6_7 .C_ON=1'b1;
    defparam \ALU.madd_cry_6_THRU_LUT4_0_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_6_THRU_LUT4_0_LC_7_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_6_THRU_LUT4_0_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__39561),
            .in2(_gnd_net_),
            .in3(N__27226),
            .lcout(\ALU.madd_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_6 ),
            .carryout(\ALU.madd_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_8_s_LC_7_7_0 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_8_s_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_8_s_LC_7_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_8_s_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__27219),
            .in2(N__27196),
            .in3(N__27181),
            .lcout(\ALU.mult_9 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\ALU.madd_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_9_0_s_LC_7_7_1 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_9_0_s_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_9_0_s_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_9_0_s_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__27178),
            .in2(N__27550),
            .in3(N__27538),
            .lcout(\ALU.mult_10 ),
            .ltout(),
            .carryin(\ALU.madd_cry_8 ),
            .carryout(\ALU.madd_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_9_THRU_LUT4_0_LC_7_7_2 .C_ON=1'b1;
    defparam \ALU.madd_cry_9_THRU_LUT4_0_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_9_THRU_LUT4_0_LC_7_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_9_THRU_LUT4_0_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27535),
            .in3(N__27490),
            .lcout(\ALU.madd_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_9 ),
            .carryout(\ALU.madd_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_11_s_LC_7_7_3 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_11_s_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_11_s_LC_7_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_11_s_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__27487),
            .in2(N__27460),
            .in3(N__27445),
            .lcout(\ALU.mult_12 ),
            .ltout(),
            .carryin(\ALU.madd_cry_10 ),
            .carryout(\ALU.madd_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_12_0_s_LC_7_7_4 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_12_0_s_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_12_0_s_LC_7_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_12_0_s_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__27442),
            .in2(N__27430),
            .in3(N__27397),
            .lcout(\ALU.mult_13 ),
            .ltout(),
            .carryin(\ALU.madd_cry_11 ),
            .carryout(\ALU.madd_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_13_0_s_LC_7_7_5 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_13_0_s_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_13_0_s_LC_7_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_13_0_s_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__27394),
            .in2(N__27379),
            .in3(N__27364),
            .lcout(\ALU.mult_14 ),
            .ltout(),
            .carryin(\ALU.madd_cry_12 ),
            .carryout(\ALU.madd_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_13_THRU_LUT4_0_LC_7_7_6 .C_ON=1'b0;
    defparam \ALU.madd_cry_13_THRU_LUT4_0_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_13_THRU_LUT4_0_LC_7_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_13_THRU_LUT4_0_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27361),
            .lcout(\ALU.madd_cry_13_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_398_0_LC_7_7_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_398_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_398_0_LC_7_7_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_398_0_LC_7_7_7  (
            .in0(N__27343),
            .in1(N__27328),
            .in2(N__27316),
            .in3(N__27307),
            .lcout(\ALU.madd_398_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJJH11_0_LC_7_8_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIJJH11_0_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJJH11_0_LC_7_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r4_RNIJJH11_0_LC_7_8_0  (
            .in0(N__27629),
            .in1(N__27680),
            .in2(_gnd_net_),
            .in3(N__30978),
            .lcout(\ALU.r4_RNIJJH11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIBROO_0_LC_7_8_1 .C_ON=1'b0;
    defparam \ALU.r0_RNIBROO_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIBROO_0_LC_7_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r0_RNIBROO_0_LC_7_8_1  (
            .in0(N__30979),
            .in1(N__34854),
            .in2(_gnd_net_),
            .in3(N__34941),
            .lcout(),
            .ltout(\ALU.r0_RNIBROOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIVVDO2_0_LC_7_8_2 .C_ON=1'b0;
    defparam \ALU.r0_RNIVVDO2_0_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIVVDO2_0_LC_7_8_2 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \ALU.r0_RNIVVDO2_0_LC_7_8_2  (
            .in0(N__27763),
            .in1(N__30928),
            .in2(N__27757),
            .in3(N__27720),
            .lcout(\ALU.a_7_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_0_LC_7_8_4.C_ON=1'b0;
    defparam TXbuffer_RNO_7_0_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_0_LC_7_8_4.LUT_INIT=16'b0000110100111101;
    LogicCell40 TXbuffer_RNO_7_0_LC_7_8_4 (
            .in0(N__34942),
            .in1(N__30067),
            .in2(N__30416),
            .in3(N__39438),
            .lcout(),
            .ltout(TXbuffer_18_3_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_0_LC_7_8_5.C_ON=1'b0;
    defparam TXbuffer_RNO_5_0_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_0_LC_7_8_5.LUT_INIT=16'b1000111110000011;
    LogicCell40 TXbuffer_RNO_5_0_LC_7_8_5 (
            .in0(N__27681),
            .in1(N__30079),
            .in2(N__27658),
            .in3(N__34065),
            .lcout(TXbuffer_RNO_5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_0_LC_7_8_6.C_ON=1'b0;
    defparam TXbuffer_RNO_3_0_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_0_LC_7_8_6.LUT_INIT=16'b0000110100111101;
    LogicCell40 TXbuffer_RNO_3_0_LC_7_8_6 (
            .in0(N__34855),
            .in1(N__30066),
            .in2(N__30415),
            .in3(N__30656),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_0_LC_7_8_7.C_ON=1'b0;
    defparam TXbuffer_RNO_0_0_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_0_LC_7_8_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_0_0_LC_7_8_7 (
            .in0(N__30068),
            .in1(N__33717),
            .in2(N__27640),
            .in3(N__27630),
            .lcout(TXbuffer_RNO_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_1_1_LC_7_9_0.C_ON=1'b0;
    defparam TXbuffer_RNO_1_1_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_1_1_LC_7_9_0.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_1_1_LC_7_9_0 (
            .in0(N__30060),
            .in1(N__27785),
            .in2(N__27559),
            .in3(N__29429),
            .lcout(TXbuffer_RNO_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_4_1_LC_7_9_1.C_ON=1'b0;
    defparam TXbuffer_RNO_4_1_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_4_1_LC_7_9_1.LUT_INIT=16'b0011010000110111;
    LogicCell40 TXbuffer_RNO_4_1_LC_7_9_1 (
            .in0(N__27589),
            .in1(N__30371),
            .in2(N__30081),
            .in3(N__28701),
            .lcout(TXbuffer_18_13_ns_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_1_LC_7_9_2.C_ON=1'b0;
    defparam TXbuffer_RNO_3_1_LC_7_9_2.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_1_LC_7_9_2.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_3_1_LC_7_9_2 (
            .in0(N__30061),
            .in1(N__31010),
            .in2(N__30397),
            .in3(N__32959),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_1_LC_7_9_3.C_ON=1'b0;
    defparam TXbuffer_RNO_0_1_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_1_LC_7_9_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_0_1_LC_7_9_3 (
            .in0(N__30058),
            .in1(N__33691),
            .in2(N__28000),
            .in3(N__33664),
            .lcout(),
            .ltout(TXbuffer_RNO_0Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_1_LC_7_9_4.C_ON=1'b0;
    defparam TXbuffer_1_LC_7_9_4.SEQ_MODE=4'b1000;
    defparam TXbuffer_1_LC_7_9_4.LUT_INIT=16'b1101010110010001;
    LogicCell40 TXbuffer_1_LC_7_9_4 (
            .in0(N__27997),
            .in1(N__49970),
            .in2(N__27982),
            .in3(N__27979),
            .lcout(TXbufferZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56261),
            .ce(N__56048),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_2_LC_7_9_5.C_ON=1'b0;
    defparam TXbuffer_RNO_3_2_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_2_LC_7_9_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_3_2_LC_7_9_5 (
            .in0(N__30054),
            .in1(N__27972),
            .in2(N__30396),
            .in3(N__33388),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_2_LC_7_9_6.C_ON=1'b0;
    defparam TXbuffer_RNO_0_2_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_2_LC_7_9_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_0_2_LC_7_9_6 (
            .in0(N__30059),
            .in1(N__27936),
            .in2(N__27898),
            .in3(N__33634),
            .lcout(TXbuffer_RNO_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r7_6_LC_7_10_0 .C_ON=1'b0;
    defparam \ALU.r7_6_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_6_LC_7_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_6_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38874),
            .lcout(r7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_7_LC_7_10_1 .C_ON=1'b0;
    defparam \ALU.r7_7_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_7_LC_7_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_7_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38740),
            .lcout(r7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_8_LC_7_10_2 .C_ON=1'b0;
    defparam \ALU.r7_8_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_8_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_8_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39524),
            .lcout(r7_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_9_LC_7_10_3 .C_ON=1'b0;
    defparam \ALU.r7_9_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_9_LC_7_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r7_9_LC_7_10_3  (
            .in0(N__34027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r7_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_1_LC_7_10_4 .C_ON=1'b0;
    defparam \ALU.r7_1_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_1_LC_7_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_1_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42147),
            .lcout(r7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_2_LC_7_10_5 .C_ON=1'b0;
    defparam \ALU.r7_2_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_2_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_2_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40287),
            .lcout(r7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_3_LC_7_10_6 .C_ON=1'b0;
    defparam \ALU.r7_3_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_3_LC_7_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_3_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50188),
            .lcout(r7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r7_4_LC_7_10_7 .C_ON=1'b0;
    defparam \ALU.r7_4_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r7_4_LC_7_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r7_4_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39083),
            .lcout(r7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56266),
            .ce(N__45888),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_0_LC_7_11_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_0_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_10_s0_c_RNO_0_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__33010),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\ALU.r0_12_prm_8_10_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s0_c_LC_7_11_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_10_s0_c_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s0_c_LC_7_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_10_s0_c_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__42342),
            .in2(N__41998),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_10_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_10_s0_c_LC_7_11_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_10_s0_c_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_10_s0_c_LC_7_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_10_s0_c_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__34513),
            .in2(N__51562),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_10_s0 ),
            .carryout(\ALU.r0_12_prm_7_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_10_s0_c_LC_7_11_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_10_s0_c_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_10_s0_c_LC_7_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_10_s0_c_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__34737),
            .in2(N__35257),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_10_s0 ),
            .carryout(\ALU.r0_12_prm_6_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_10_s0_c_LC_7_11_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_10_s0_c_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_10_s0_c_LC_7_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_10_s0_c_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__34698),
            .in2(N__45565),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_10_s0 ),
            .carryout(\ALU.r0_12_prm_5_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_10_s0_c_inv_LC_7_11_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_10_s0_c_inv_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_10_s0_c_inv_LC_7_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_10_s0_c_inv_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__34665),
            .in2(N__34612),
            .in3(N__51794),
            .lcout(\ALU.a_i_10 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_10_s0 ),
            .carryout(\ALU.r0_12_prm_4_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_10_s0_c_inv_LC_7_11_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_10_s0_c_inv_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_10_s0_c_inv_LC_7_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_10_s0_c_inv_LC_7_11_6  (
            .in0(N__55167),
            .in1(N__28213),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_10_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_10_s0 ),
            .carryout(\ALU.r0_12_prm_3_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_10_s0_c_LC_7_11_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_10_s0_c_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_10_s0_c_LC_7_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_10_s0_c_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__35641),
            .in2(N__35857),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_10_s0 ),
            .carryout(\ALU.r0_12_prm_2_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_10_s0_c_LC_7_12_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_10_s0_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_10_s0_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_10_s0_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__36109),
            .in2(N__34201),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\ALU.r0_12_s0_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_10_s0_c_RNI4UV4363_LC_7_12_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_10_s0_c_RNI4UV4363_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_10_s0_c_RNI4UV4363_LC_7_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r0_12_prm_1_10_s0_c_RNI4UV4363_LC_7_12_1  (
            .in0(N__28207),
            .in1(N__34639),
            .in2(_gnd_net_),
            .in3(N__28195),
            .lcout(\ALU.r0_12_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_10_LC_7_12_2 .C_ON=1'b0;
    defparam \ALU.r0_10_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_10_LC_7_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_10_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28158),
            .lcout(r0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56274),
            .ce(N__49719),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_0_LC_7_13_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_0_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_0_LC_7_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_14_s0_c_RNO_0_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__46525),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\ALU.r0_12_prm_8_14_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s0_c_LC_7_13_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_14_s0_c_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s0_c_LC_7_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_14_s0_c_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__47980),
            .in2(N__39634),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_14_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_14_s0_c_LC_7_13_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_14_s0_c_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_14_s0_c_LC_7_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_14_s0_c_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__47928),
            .in2(N__42955),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_14_s0 ),
            .carryout(\ALU.r0_12_prm_7_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_14_s0_c_LC_7_13_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_14_s0_c_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_14_s0_c_LC_7_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_14_s0_c_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__47895),
            .in2(N__39646),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_14_s0 ),
            .carryout(\ALU.r0_12_prm_6_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_14_s0_c_LC_7_13_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_14_s0_c_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_14_s0_c_LC_7_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_14_s0_c_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__39667),
            .in2(N__47866),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_14_s0 ),
            .carryout(\ALU.r0_12_prm_5_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_14_s0_c_inv_LC_7_13_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_14_s0_c_inv_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_14_s0_c_inv_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_14_s0_c_inv_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__47823),
            .in2(N__39685),
            .in3(N__46959),
            .lcout(\ALU.a_i_14 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_14_s0 ),
            .carryout(\ALU.r0_12_prm_4_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_14_s0_c_inv_LC_7_13_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_14_s0_c_inv_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_14_s0_c_inv_LC_7_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_14_s0_c_inv_LC_7_13_6  (
            .in0(N__55168),
            .in1(_gnd_net_),
            .in2(N__28336),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_14_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_14_s0 ),
            .carryout(\ALU.r0_12_prm_3_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_14_s0_c_LC_7_13_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_14_s0_c_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_14_s0_c_LC_7_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_14_s0_c_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__49140),
            .in2(N__36052),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_14_s0 ),
            .carryout(\ALU.r0_12_prm_2_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_14_s0_c_LC_7_14_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_14_s0_c_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_14_s0_c_LC_7_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_14_s0_c_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__49083),
            .in2(N__31216),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\ALU.r0_12_s0_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_14_s0_c_RNI357RUG3_LC_7_14_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_14_s0_c_RNI357RUG3_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_14_s0_c_RNI357RUG3_LC_7_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r0_12_prm_1_14_s0_c_RNI357RUG3_LC_7_14_1  (
            .in0(N__28327),
            .in1(N__49033),
            .in2(_gnd_net_),
            .in3(N__28315),
            .lcout(\ALU.r0_12_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_14_LC_7_14_2 .C_ON=1'b0;
    defparam \ALU.r1_14_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_14_LC_7_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_14_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28293),
            .lcout(r1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56284),
            .ce(N__47569),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_0_LC_7_15_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_0_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_0_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_12_s0_c_RNO_0_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__35656),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\ALU.r0_12_prm_8_12_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s0_c_LC_7_15_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_12_s0_c_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s0_c_LC_7_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_12_s0_c_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__37468),
            .in2(N__34480),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_12_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_12_s0_c_LC_7_15_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_12_s0_c_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_12_s0_c_LC_7_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_12_s0_c_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__37437),
            .in2(N__31285),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_12_s0 ),
            .carryout(\ALU.r0_12_prm_7_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_12_s0_c_LC_7_15_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_12_s0_c_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_12_s0_c_LC_7_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_12_s0_c_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__37410),
            .in2(N__31270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_12_s0 ),
            .carryout(\ALU.r0_12_prm_6_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_12_s0_c_LC_7_15_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_12_s0_c_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_12_s0_c_LC_7_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_12_s0_c_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__37369),
            .in2(N__31318),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_12_s0 ),
            .carryout(\ALU.r0_12_prm_5_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_12_s0_c_inv_LC_7_15_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_12_s0_c_inv_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_12_s0_c_inv_LC_7_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_12_s0_c_inv_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__37323),
            .in2(N__36175),
            .in3(N__41350),
            .lcout(\ALU.a_i_12 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_12_s0 ),
            .carryout(\ALU.r0_12_prm_4_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_12_s0_c_inv_LC_7_15_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_12_s0_c_inv_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_12_s0_c_inv_LC_7_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_12_s0_c_inv_LC_7_15_6  (
            .in0(N__55166),
            .in1(N__28465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_12_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_12_s0 ),
            .carryout(\ALU.r0_12_prm_3_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_12_s0_c_LC_7_15_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_12_s0_c_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_12_s0_c_LC_7_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_12_s0_c_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__37654),
            .in2(N__35695),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_12_s0 ),
            .carryout(\ALU.r0_12_prm_2_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_12_s0_c_LC_7_16_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_12_s0_c_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_12_s0_c_LC_7_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_12_s0_c_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__37594),
            .in2(N__36064),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\ALU.r0_12_s0_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_12_s0_c_RNIS2VGA6_LC_7_16_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_12_s0_c_RNIS2VGA6_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_12_s0_c_RNIS2VGA6_LC_7_16_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r0_12_prm_1_12_s0_c_RNIS2VGA6_LC_7_16_1  (
            .in0(N__37552),
            .in1(N__28459),
            .in2(_gnd_net_),
            .in3(N__28450),
            .lcout(\ALU.r0_12_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_LC_7_16_2 .C_ON=1'b0;
    defparam \ALU.r0_12_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_12_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28402),
            .lcout(r0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56291),
            .ce(N__49718),
            .sr(_gnd_net_));
    defparam TXbuffer_5_LC_7_17_2.C_ON=1'b0;
    defparam TXbuffer_5_LC_7_17_2.SEQ_MODE=4'b1000;
    defparam TXbuffer_5_LC_7_17_2.LUT_INIT=16'b1100000010101111;
    LogicCell40 TXbuffer_5_LC_7_17_2 (
            .in0(N__28510),
            .in1(N__28501),
            .in2(N__49967),
            .in3(N__28492),
            .lcout(TXbufferZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56295),
            .ce(N__56039),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_1_LC_9_1_0 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_1_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_1_LC_9_1_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \ALU.mult_a2_b_1_LC_9_1_0  (
            .in0(N__32548),
            .in1(N__32692),
            .in2(N__32277),
            .in3(N__46797),
            .lcout(\ALU.a2_b_1 ),
            .ltout(\ALU.a2_b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_8_LC_9_1_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_8_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_8_LC_9_1_1 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_8_LC_9_1_1  (
            .in0(N__28480),
            .in1(N__49353),
            .in2(N__28483),
            .in3(N__37994),
            .lcout(\ALU.madd_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a1_b_2_LC_9_1_2 .C_ON=1'b0;
    defparam \ALU.mult_a1_b_2_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a1_b_2_LC_9_1_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a1_b_2_LC_9_1_2  (
            .in0(N__31666),
            .in1(N__31719),
            .in2(N__32276),
            .in3(N__43931),
            .lcout(\ALU.a1_b_2 ),
            .ltout(\ALU.a1_b_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_4_LC_9_1_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_4_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_4_LC_9_1_3 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_4_LC_9_1_3  (
            .in0(N__28474),
            .in1(N__49352),
            .in2(N__28468),
            .in3(N__37993),
            .lcout(\ALU.madd_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_3_c_RNO_LC_9_1_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_3_c_RNO_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_3_c_RNO_LC_9_1_4 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_3_c_RNO_LC_9_1_4  (
            .in0(N__44359),
            .in1(N__53951),
            .in2(N__53216),
            .in3(N__49360),
            .lcout(\ALU.r0_12_prm_6_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a2_b_0_LC_9_1_5 .C_ON=1'b0;
    defparam \ALU.mult_a2_b_0_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a2_b_0_LC_9_1_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a2_b_0_LC_9_1_5  (
            .in0(N__32691),
            .in1(N__32549),
            .in2(N__32236),
            .in3(N__37992),
            .lcout(\ALU.a2_b_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_2_c_RNO_LC_9_1_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_2_c_RNO_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_2_c_RNO_LC_9_1_6 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_2_c_RNO_LC_9_1_6  (
            .in0(N__54553),
            .in1(N__48402),
            .in2(N__53217),
            .in3(N__43932),
            .lcout(\ALU.r0_12_prm_5_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIL9636_2_LC_9_1_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIL9636_2_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIL9636_2_LC_9_1_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r4_RNIL9636_2_LC_9_1_7  (
            .in0(N__48403),
            .in1(N__53090),
            .in2(N__54047),
            .in3(N__54554),
            .lcout(\ALU.r4_RNIL9636Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_39_LC_9_2_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_39_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_39_LC_9_2_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_39_LC_9_2_0  (
            .in0(N__28621),
            .in1(N__28606),
            .in2(N__29563),
            .in3(N__28597),
            .lcout(\ALU.madd_39 ),
            .ltout(\ALU.madd_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_45_LC_9_2_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_45_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_45_LC_9_2_1 .LUT_INIT=16'b1110000010000000;
    LogicCell40 \ALU.mult_madd_45_LC_9_2_1  (
            .in0(N__31591),
            .in1(N__28918),
            .in2(N__28582),
            .in3(N__28537),
            .lcout(\ALU.madd_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI97EK9_5_LC_9_2_2 .C_ON=1'b0;
    defparam \ALU.r4_RNI97EK9_5_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI97EK9_5_LC_9_2_2 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r4_RNI97EK9_5_LC_9_2_2  (
            .in0(N__53949),
            .in1(N__45360),
            .in2(N__54787),
            .in3(N__43365),
            .lcout(\ALU.lshift_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_23_LC_9_2_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_23_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_23_LC_9_2_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_23_LC_9_2_3  (
            .in0(N__31590),
            .in1(N__28917),
            .in2(_gnd_net_),
            .in3(N__28536),
            .lcout(),
            .ltout(\ALU.madd_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_4_l_fx_LC_9_2_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_4_l_fx_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_4_l_fx_LC_9_2_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ALU.mult_madd_axb_4_l_fx_LC_9_2_4  (
            .in0(_gnd_net_),
            .in1(N__28579),
            .in2(N__28573),
            .in3(N__28570),
            .lcout(\ALU.madd_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_19_LC_9_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_19_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_19_LC_9_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_19_LC_9_2_5  (
            .in0(N__31589),
            .in1(N__28916),
            .in2(_gnd_net_),
            .in3(N__28535),
            .lcout(\ALU.madd_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIM8HG5_5_LC_9_2_6 .C_ON=1'b0;
    defparam \ALU.r4_RNIM8HG5_5_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIM8HG5_5_LC_9_2_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r4_RNIM8HG5_5_LC_9_2_6  (
            .in0(N__53950),
            .in1(N__53159),
            .in2(N__54788),
            .in3(N__45361),
            .lcout(\ALU.r4_RNIM8HG5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_1_LC_9_2_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_1_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_1_LC_9_2_7 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_axb_1_LC_9_2_7  (
            .in0(N__41942),
            .in1(N__48955),
            .in2(N__29319),
            .in3(N__43947),
            .lcout(\ALU.madd_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_0_s1_c_RNO_LC_9_3_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_3_0_s1_c_RNO_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_0_s1_c_RNO_LC_9_3_0 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \ALU.r0_12_prm_3_0_s1_c_RNO_LC_9_3_0  (
            .in0(N__48944),
            .in1(N__38028),
            .in2(_gnd_net_),
            .in3(N__55230),
            .lcout(\ALU.r0_12_prm_3_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_66_LC_9_3_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_66_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_66_LC_9_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.mult_madd_66_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(N__28893),
            .in2(_gnd_net_),
            .in3(N__28868),
            .lcout(\ALU.madd_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKO1J4_5_LC_9_3_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIKO1J4_5_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKO1J4_5_LC_9_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIKO1J4_5_LC_9_3_2  (
            .in0(N__29237),
            .in1(N__29076),
            .in2(_gnd_net_),
            .in3(N__29004),
            .lcout(\ALU.a_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_4_LC_9_3_3 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_4_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_4_LC_9_3_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a0_b_4_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(N__48943),
            .in2(_gnd_net_),
            .in3(N__40523),
            .lcout(\ALU.a0_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIUM9JC_2_LC_9_3_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIUM9JC_2_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIUM9JC_2_LC_9_3_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNIUM9JC_2_LC_9_3_4  (
            .in0(_gnd_net_),
            .in1(N__33936),
            .in2(_gnd_net_),
            .in3(N__28906),
            .lcout(\ALU.r4_RNIUM9JCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_6_ma_LC_9_3_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_6_ma_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_6_ma_LC_9_3_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_cry_6_ma_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(N__28894),
            .in2(_gnd_net_),
            .in3(N__28869),
            .lcout(\ALU.madd_cry_6_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_0_s0_c_RNO_LC_9_3_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_0_s0_c_RNO_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_0_s0_c_RNO_LC_9_3_6 .LUT_INIT=16'b1110000100010001;
    LogicCell40 \ALU.r0_12_prm_6_0_s0_c_RNO_LC_9_3_6  (
            .in0(N__48945),
            .in1(N__38029),
            .in2(N__53213),
            .in3(N__53804),
            .lcout(\ALU.r0_12_prm_6_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI18BO_0_LC_9_4_0 .C_ON=1'b0;
    defparam \ALU.r2_RNI18BO_0_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI18BO_0_LC_9_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r2_RNI18BO_0_LC_9_4_0  (
            .in0(N__28840),
            .in1(N__28724),
            .in2(_gnd_net_),
            .in3(N__28798),
            .lcout(\ALU.r2_RNI18BOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_0_LC_9_4_1 .C_ON=1'b0;
    defparam \ALU.r2_0_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r2_0_LC_9_4_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ALU.r2_0_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__34987),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56245),
            .ce(N__47671),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI4H0S_1_LC_9_4_2 .C_ON=1'b0;
    defparam \ALU.r2_RNI4H0S_1_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI4H0S_1_LC_9_4_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r2_RNI4H0S_1_LC_9_4_2  (
            .in0(N__28705),
            .in1(N__28663),
            .in2(_gnd_net_),
            .in3(N__29518),
            .lcout(\ALU.r2_RNI4H0SZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_RNIC9P41_1_LC_9_4_3 .C_ON=1'b0;
    defparam \ALU.r6_RNIC9P41_1_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r6_RNIC9P41_1_LC_9_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r6_RNIC9P41_1_LC_9_4_3  (
            .in0(N__29517),
            .in1(N__29440),
            .in2(_gnd_net_),
            .in3(N__29407),
            .lcout(\ALU.r6_RNIC9P41Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIDAOQ3_2_LC_9_4_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIDAOQ3_2_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIDAOQ3_2_LC_9_4_4 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \ALU.r4_RNIDAOQ3_2_LC_9_4_4  (
            .in0(N__33340),
            .in1(N__32862),
            .in2(_gnd_net_),
            .in3(N__29365),
            .lcout(\ALU.b_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIHU8AD1_15_LC_9_4_5 .C_ON=1'b0;
    defparam \ALU.r5_RNIHU8AD1_15_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIHU8AD1_15_LC_9_4_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r5_RNIHU8AD1_15_LC_9_4_5  (
            .in0(N__37498),
            .in1(N__51509),
            .in2(_gnd_net_),
            .in3(N__31333),
            .lcout(\ALU.rshift_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_3_LC_9_4_6 .C_ON=1'b0;
    defparam \ALU.mult_a0_b_3_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_3_LC_9_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_a0_b_3_LC_9_4_6  (
            .in0(N__44335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48998),
            .lcout(\ALU.a0_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNID26E8_0_LC_9_4_7 .C_ON=1'b0;
    defparam \ALU.r4_RNID26E8_0_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNID26E8_0_LC_9_4_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ALU.r4_RNID26E8_0_LC_9_4_7  (
            .in0(N__48999),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37988),
            .lcout(\ALU.un14_log_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_13_LC_9_5_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_13_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_13_LC_9_5_0 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_13_LC_9_5_0  (
            .in0(N__29290),
            .in1(_gnd_net_),
            .in2(N__29299),
            .in3(N__29275),
            .lcout(\ALU.madd_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_3_LC_9_5_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_3_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_3_LC_9_5_1 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_3_LC_9_5_1  (
            .in0(N__41951),
            .in1(N__48983),
            .in2(N__29320),
            .in3(N__43916),
            .lcout(\ALU.madd_3 ),
            .ltout(\ALU.madd_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_2_LC_9_5_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_2_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_2_LC_9_5_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_axb_2_LC_9_5_2  (
            .in0(N__29289),
            .in1(_gnd_net_),
            .in2(N__29278),
            .in3(N__29274),
            .lcout(\ALU.madd_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI7AQC9_15_LC_9_5_3 .C_ON=1'b0;
    defparam \ALU.r2_RNI7AQC9_15_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI7AQC9_15_LC_9_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r2_RNI7AQC9_15_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__40175),
            .in2(_gnd_net_),
            .in3(N__40009),
            .lcout(\ALU.un14_log_0_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_1_c_RNO_LC_9_5_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_1_c_RNO_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_1_c_RNO_LC_9_5_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_7_1_c_RNO_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__53098),
            .in2(_gnd_net_),
            .in3(N__41952),
            .lcout(\ALU.r0_12_prm_7_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_2_LC_9_5_5 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_2_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_2_LC_9_5_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a3_b_2_LC_9_5_5  (
            .in0(N__31934),
            .in1(N__31829),
            .in2(N__32272),
            .in3(N__43915),
            .lcout(\ALU.a3_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIRCFPA_0_7_LC_9_5_6 .C_ON=1'b0;
    defparam \ALU.r4_RNIRCFPA_0_7_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIRCFPA_0_7_LC_9_5_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r4_RNIRCFPA_0_7_LC_9_5_6  (
            .in0(N__53742),
            .in1(N__46151),
            .in2(N__54697),
            .in3(N__44552),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI67NNK_10_LC_9_5_7 .C_ON=1'b0;
    defparam \ALU.r5_RNI67NNK_10_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI67NNK_10_LC_9_5_7 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r5_RNI67NNK_10_LC_9_5_7  (
            .in0(N__54520),
            .in1(N__52151),
            .in2(N__29539),
            .in3(N__51805),
            .lcout(\ALU.r5_RNI67NNKZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_2_LC_9_6_0 .C_ON=1'b0;
    defparam \ALU.r1_2_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_2_LC_9_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_2_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40274),
            .lcout(r1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56250),
            .ce(N__47581),
            .sr(_gnd_net_));
    defparam \ALU.r1_3_LC_9_6_1 .C_ON=1'b0;
    defparam \ALU.r1_3_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_3_LC_9_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_3_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50171),
            .lcout(r1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56250),
            .ce(N__47581),
            .sr(_gnd_net_));
    defparam \ALU.r1_4_LC_9_6_2 .C_ON=1'b0;
    defparam \ALU.r1_4_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_4_LC_9_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_4_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39052),
            .lcout(r1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56250),
            .ce(N__47581),
            .sr(_gnd_net_));
    defparam \ALU.r1_1_LC_9_6_5 .C_ON=1'b0;
    defparam \ALU.r1_1_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_1_LC_9_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_1_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42129),
            .lcout(r1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56250),
            .ce(N__47581),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIJEMP_7_LC_9_7_0 .C_ON=1'b0;
    defparam \ALU.r0_RNIJEMP_7_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIJEMP_7_LC_9_7_0 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \ALU.r0_RNIJEMP_7_LC_9_7_0  (
            .in0(N__36917),
            .in1(N__30740),
            .in2(N__33304),
            .in3(N__33184),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI82OE1_7_LC_9_7_1 .C_ON=1'b0;
    defparam \ALU.r4_RNI82OE1_7_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI82OE1_7_LC_9_7_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r4_RNI82OE1_7_LC_9_7_1  (
            .in0(N__33744),
            .in1(N__34089),
            .in2(N__29536),
            .in3(N__33138),
            .lcout(\ALU.r4_RNI82OE1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_7_LC_9_7_2 .C_ON=1'b0;
    defparam \ALU.r0_7_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_7_LC_9_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_7_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38727),
            .lcout(r0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56254),
            .ce(N__49756),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_3_7_LC_9_7_3.C_ON=1'b0;
    defparam TXbuffer_RNO_3_7_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_3_7_LC_9_7_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 TXbuffer_RNO_3_7_LC_9_7_3 (
            .in0(N__30084),
            .in1(N__30487),
            .in2(N__30418),
            .in3(N__36918),
            .lcout(),
            .ltout(TXbuffer_18_10_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_0_7_LC_9_7_4.C_ON=1'b0;
    defparam TXbuffer_RNO_0_7_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_0_7_LC_9_7_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 TXbuffer_RNO_0_7_LC_9_7_4 (
            .in0(N__30083),
            .in1(N__30451),
            .in2(N__30421),
            .in3(N__33745),
            .lcout(TXbuffer_RNO_0Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_7_7_LC_9_7_5.C_ON=1'b0;
    defparam TXbuffer_RNO_7_7_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_7_7_LC_9_7_5.LUT_INIT=16'b0000110100111101;
    LogicCell40 TXbuffer_RNO_7_7_LC_9_7_5 (
            .in0(N__30741),
            .in1(N__30082),
            .in2(N__30417),
            .in3(N__30118),
            .lcout(),
            .ltout(TXbuffer_18_3_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_5_7_LC_9_7_6.C_ON=1'b0;
    defparam TXbuffer_RNO_5_7_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_5_7_LC_9_7_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 TXbuffer_RNO_5_7_LC_9_7_6 (
            .in0(N__34090),
            .in1(N__30085),
            .in2(N__29728),
            .in3(N__29725),
            .lcout(),
            .ltout(TXbuffer_RNO_5Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_RNO_2_7_LC_9_7_7.C_ON=1'b0;
    defparam TXbuffer_RNO_2_7_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam TXbuffer_RNO_2_7_LC_9_7_7.LUT_INIT=16'b0100010101100111;
    LogicCell40 TXbuffer_RNO_2_7_LC_9_7_7 (
            .in0(N__29683),
            .in1(N__49940),
            .in2(N__29587),
            .in3(N__29584),
            .lcout(TXbuffer_18_15_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI5IT71_1_LC_9_8_0 .C_ON=1'b0;
    defparam \ALU.r0_RNI5IT71_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI5IT71_1_LC_9_8_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r0_RNI5IT71_1_LC_9_8_0  (
            .in0(N__30971),
            .in1(N__32955),
            .in2(N__31095),
            .in3(N__35082),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIDI992_1_LC_9_8_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIDI992_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIDI992_1_LC_9_8_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNIDI992_1_LC_9_8_1  (
            .in0(N__30571),
            .in1(N__33653),
            .in2(N__29566),
            .in3(N__34361),
            .lcout(\ALU.r4_RNIDI992Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam a_fast_0_LC_9_8_2.C_ON=1'b0;
    defparam a_fast_0_LC_9_8_2.SEQ_MODE=4'b1000;
    defparam a_fast_0_LC_9_8_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 a_fast_0_LC_9_8_2 (
            .in0(N__30974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(a_fastZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56255),
            .ce(N__56050),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIHUT71_7_LC_9_8_3 .C_ON=1'b0;
    defparam \ALU.r0_RNIHUT71_7_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIHUT71_7_LC_9_8_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNIHUT71_7_LC_9_8_3  (
            .in0(N__30751),
            .in1(N__31086),
            .in2(N__36922),
            .in3(N__30973),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI6BA92_7_LC_9_8_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI6BA92_7_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI6BA92_7_LC_9_8_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNI6BA92_7_LC_9_8_4  (
            .in0(N__30936),
            .in1(N__34083),
            .in2(N__30727),
            .in3(N__33738),
            .lcout(\ALU.r4_RNI6BA92Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIJ0U71_8_LC_9_8_5 .C_ON=1'b0;
    defparam \ALU.r0_RNIJ0U71_8_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIJ0U71_8_LC_9_8_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNIJ0U71_8_LC_9_8_5  (
            .in0(N__39431),
            .in1(N__31088),
            .in2(N__30664),
            .in3(N__30972),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIAFA92_8_LC_9_8_6 .C_ON=1'b0;
    defparam \ALU.r4_RNIAFA92_8_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIAFA92_8_LC_9_8_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNIAFA92_8_LC_9_8_6  (
            .in0(N__30937),
            .in1(N__34055),
            .in2(N__30625),
            .in3(N__33716),
            .lcout(\ALU.r4_RNIAFA92Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI9MT71_3_LC_9_8_7 .C_ON=1'b0;
    defparam \ALU.r0_RNI9MT71_3_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI9MT71_3_LC_9_8_7 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNI9MT71_3_LC_9_8_7  (
            .in0(N__35049),
            .in1(N__31087),
            .in2(N__33237),
            .in3(N__30970),
            .lcout(\ALU.a_3_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI7KT71_2_LC_9_9_0 .C_ON=1'b0;
    defparam \ALU.r0_RNI7KT71_2_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI7KT71_2_LC_9_9_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNI7KT71_2_LC_9_9_0  (
            .in0(N__33407),
            .in1(N__31068),
            .in2(N__33384),
            .in3(N__30975),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIHM992_2_LC_9_9_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIHM992_2_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIHM992_2_LC_9_9_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.r4_RNIHM992_2_LC_9_9_1  (
            .in0(N__33627),
            .in1(N__34325),
            .in2(N__30574),
            .in3(N__30569),
            .lcout(\ALU.r4_RNIHM992Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_2_LC_9_9_2 .C_ON=1'b0;
    defparam \ALU.r0_2_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_2_LC_9_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_2_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40288),
            .lcout(r0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56256),
            .ce(N__49731),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIBOT71_4_LC_9_9_3 .C_ON=1'b0;
    defparam \ALU.r0_RNIBOT71_4_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIBOT71_4_LC_9_9_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r0_RNIBOT71_4_LC_9_9_3  (
            .in0(N__30977),
            .in1(N__33467),
            .in2(N__31085),
            .in3(N__33497),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIQU992_4_LC_9_9_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIQU992_4_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIQU992_4_LC_9_9_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNIQU992_4_LC_9_9_4  (
            .in0(N__30930),
            .in1(N__33561),
            .in2(N__31099),
            .in3(N__34290),
            .lcout(\ALU.r4_RNIQU992Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_4_LC_9_9_5 .C_ON=1'b0;
    defparam \ALU.r0_4_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_4_LC_9_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r0_4_LC_9_9_5  (
            .in0(N__39078),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56256),
            .ce(N__49731),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIL2U71_9_LC_9_9_6 .C_ON=1'b0;
    defparam \ALU.r0_RNIL2U71_9_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIL2U71_9_LC_9_9_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNIL2U71_9_LC_9_9_6  (
            .in0(N__31134),
            .in1(N__31067),
            .in2(N__31012),
            .in3(N__30976),
            .lcout(),
            .ltout(\ALU.a_3_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIEJA92_9_LC_9_9_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIEJA92_9_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIEJA92_9_LC_9_9_7 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.r4_RNIEJA92_9_LC_9_9_7  (
            .in0(N__34391),
            .in1(N__30929),
            .in2(N__30817),
            .in3(N__33680),
            .lcout(\ALU.r4_RNIEJA92Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_0_LC_9_10_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_0_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_0_LC_9_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_9_s0_c_RNO_0_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__43033),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\ALU.r0_12_prm_8_9_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s0_c_LC_9_10_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_9_s0_c_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s0_c_LC_9_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_9_s0_c_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__42586),
            .in2(N__36853),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_9_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_9_s0_c_LC_9_10_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_9_s0_c_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_9_s0_c_LC_9_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_9_s0_c_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__42541),
            .in2(N__45910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_9_s0 ),
            .carryout(\ALU.r0_12_prm_7_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_9_s0_c_LC_9_10_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_9_s0_c_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_9_s0_c_LC_9_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_9_s0_c_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__45544),
            .in2(N__30769),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_9_s0 ),
            .carryout(\ALU.r0_12_prm_6_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_9_s0_c_LC_9_10_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_9_s0_c_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_9_s0_c_LC_9_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_9_s0_c_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__42507),
            .in2(N__42037),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_9_s0 ),
            .carryout(\ALU.r0_12_prm_5_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_9_s0_c_inv_LC_9_10_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_9_s0_c_inv_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_9_s0_c_inv_LC_9_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_4_9_s0_c_inv_LC_9_10_5  (
            .in0(N__52302),
            .in1(N__42468),
            .in2(N__48100),
            .in3(_gnd_net_),
            .lcout(\ALU.a_i_9 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_9_s0 ),
            .carryout(\ALU.r0_12_prm_4_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_9_s0_c_inv_LC_9_10_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_9_s0_c_inv_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_9_s0_c_inv_LC_9_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_3_9_s0_c_inv_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__31186),
            .in2(_gnd_net_),
            .in3(N__55262),
            .lcout(\ALU.r0_12_prm_3_9_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_9_s0 ),
            .carryout(\ALU.r0_12_prm_3_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_9_s0_c_LC_9_10_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_9_s0_c_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_9_s0_c_LC_9_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_9_s0_c_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__42430),
            .in2(N__31180),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_9_s0 ),
            .carryout(\ALU.r0_12_prm_2_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_9_s0_c_LC_9_11_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_9_s0_c_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_9_s0_c_LC_9_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_9_s0_c_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__42399),
            .in2(N__35677),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\ALU.r0_12_s0_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_9_s0_c_RNI39QBSO_LC_9_11_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_9_s0_c_RNI39QBSO_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_9_s0_c_RNI39QBSO_LC_9_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r0_12_prm_1_9_s0_c_RNI39QBSO_LC_9_11_1  (
            .in0(N__31162),
            .in1(N__42970),
            .in2(_gnd_net_),
            .in3(N__31150),
            .lcout(\ALU.r0_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_9_LC_9_11_2 .C_ON=1'b0;
    defparam \ALU.r0_9_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_9_LC_9_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_9_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34015),
            .lcout(r0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56262),
            .ce(N__49732),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNISU5D9_1_9_LC_9_12_0 .C_ON=1'b0;
    defparam \ALU.r4_RNISU5D9_1_9_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNISU5D9_1_9_LC_9_12_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.r4_RNISU5D9_1_9_LC_9_12_0  (
            .in0(N__52309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47476),
            .lcout(\ALU.r4_RNISU5D9_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_LC_9_12_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_LC_9_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_11_s1_c_RNO_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__55528),
            .in2(_gnd_net_),
            .in3(N__34424),
            .lcout(\ALU.r0_12_prm_8_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIA5SI9_12_LC_9_12_2 .C_ON=1'b0;
    defparam \ALU.r5_RNIA5SI9_12_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIA5SI9_12_LC_9_12_2 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r5_RNIA5SI9_12_LC_9_12_2  (
            .in0(N__53753),
            .in1(N__41293),
            .in2(N__54557),
            .in3(N__40981),
            .lcout(\ALU.rshift_10_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_5_s0_c_RNO_LC_9_12_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_5_s0_c_RNO_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_5_s0_c_RNO_LC_9_12_3 .LUT_INIT=16'b1010100100000011;
    LogicCell40 \ALU.r0_12_prm_6_5_s0_c_RNO_LC_9_12_3  (
            .in0(N__53856),
            .in1(N__45453),
            .in2(N__45262),
            .in3(N__53196),
            .lcout(\ALU.r0_12_prm_6_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_12_s0_c_RNO_LC_9_12_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_12_s0_c_RNO_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_12_s0_c_RNO_LC_9_12_4 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_12_s0_c_RNO_LC_9_12_4  (
            .in0(N__39861),
            .in1(N__53857),
            .in2(N__53243),
            .in3(N__41294),
            .lcout(\ALU.r0_12_prm_6_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIUF9K8_0_10_LC_9_12_5 .C_ON=1'b0;
    defparam \ALU.r5_RNIUF9K8_0_10_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIUF9K8_0_10_LC_9_12_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.r5_RNIUF9K8_0_10_LC_9_12_5  (
            .in0(N__51827),
            .in1(_gnd_net_),
            .in2(N__52035),
            .in3(_gnd_net_),
            .lcout(\ALU.r5_RNIUF9K8_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_10_s1_c_RNO_LC_9_12_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_10_s1_c_RNO_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_10_s1_c_RNO_LC_9_12_6 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_10_s1_c_RNO_LC_9_12_6  (
            .in0(N__53195),
            .in1(N__52024),
            .in2(_gnd_net_),
            .in3(N__51826),
            .lcout(\ALU.r0_12_prm_7_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_15_s1_c_RNO_LC_9_12_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_15_s1_c_RNO_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_15_s1_c_RNO_LC_9_12_7 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \ALU.r0_12_prm_2_15_s1_c_RNO_LC_9_12_7  (
            .in0(N__36248),
            .in1(N__55927),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_2_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_13_s0_c_RNO_LC_9_13_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_13_s0_c_RNO_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_13_s0_c_RNO_LC_9_13_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_13_s0_c_RNO_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__55950),
            .in2(_gnd_net_),
            .in3(N__34589),
            .lcout(\ALU.r0_12_prm_2_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_14_s0_c_RNO_LC_9_13_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_14_s0_c_RNO_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_14_s0_c_RNO_LC_9_13_1 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_14_s0_c_RNO_LC_9_13_1  (
            .in0(N__55951),
            .in1(N__53758),
            .in2(_gnd_net_),
            .in3(N__49073),
            .lcout(\ALU.r0_12_prm_1_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIUF9K8_10_LC_9_13_2 .C_ON=1'b0;
    defparam \ALU.r5_RNIUF9K8_10_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIUF9K8_10_LC_9_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r5_RNIUF9K8_10_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__52028),
            .in2(_gnd_net_),
            .in3(N__51831),
            .lcout(\ALU.un14_log_0_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_LC_9_13_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_LC_9_13_4 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \ALU.r0_12_prm_8_15_s1_c_RNO_LC_9_13_4  (
            .in0(N__55529),
            .in1(N__36014),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_8_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNISMSV4_15_LC_9_13_5 .C_ON=1'b0;
    defparam \ALU.r5_RNISMSV4_15_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNISMSV4_15_LC_9_13_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.r5_RNISMSV4_15_LC_9_13_5  (
            .in0(N__54603),
            .in1(N__53757),
            .in2(_gnd_net_),
            .in3(N__40097),
            .lcout(\ALU.r5_RNISMSV4Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI465TI_13_LC_9_13_6 .C_ON=1'b0;
    defparam \ALU.r5_RNI465TI_13_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI465TI_13_LC_9_13_6 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.r5_RNI465TI_13_LC_9_13_6  (
            .in0(N__31342),
            .in1(N__46988),
            .in2(N__54777),
            .in3(N__41556),
            .lcout(\ALU.r5_RNI465TIZ0Z_13 ),
            .ltout(\ALU.r5_RNI465TIZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIOL1S71_10_LC_9_13_7 .C_ON=1'b0;
    defparam \ALU.r5_RNIOL1S71_10_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIOL1S71_10_LC_9_13_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r5_RNIOL1S71_10_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__51033),
            .in2(N__31336),
            .in3(N__32917),
            .lcout(\ALU.r5_RNIOL1S71Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNID2JJ9_13_LC_9_14_0 .C_ON=1'b0;
    defparam \ALU.r5_RNID2JJ9_13_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNID2JJ9_13_LC_9_14_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r5_RNID2JJ9_13_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__35428),
            .in2(_gnd_net_),
            .in3(N__41557),
            .lcout(\ALU.un14_log_0_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_15_s0_c_RNO_LC_9_14_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_15_s0_c_RNO_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_15_s0_c_RNO_LC_9_14_1 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_15_s0_c_RNO_LC_9_14_1  (
            .in0(N__53759),
            .in1(N__40160),
            .in2(N__53241),
            .in3(N__39992),
            .lcout(\ALU.r0_12_prm_6_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_12_s0_c_RNO_LC_9_14_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_12_s0_c_RNO_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_12_s0_c_RNO_LC_9_14_2 .LUT_INIT=16'b0110100111000011;
    LogicCell40 \ALU.r0_12_prm_5_12_s0_c_RNO_LC_9_14_2  (
            .in0(N__54582),
            .in1(N__39874),
            .in2(N__41368),
            .in3(N__53194),
            .lcout(\ALU.r0_12_prm_5_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_10_s1_c_RNO_LC_9_14_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_10_s1_c_RNO_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_10_s1_c_RNO_LC_9_14_3 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_10_s1_c_RNO_LC_9_14_3  (
            .in0(N__51832),
            .in1(N__54581),
            .in2(N__53242),
            .in3(N__52002),
            .lcout(\ALU.r0_12_prm_5_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI7AQC9_1_15_LC_9_14_4 .C_ON=1'b0;
    defparam \ALU.r2_RNI7AQC9_1_15_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI7AQC9_1_15_LC_9_14_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ALU.r2_RNI7AQC9_1_15_LC_9_14_4  (
            .in0(N__39994),
            .in1(_gnd_net_),
            .in2(N__40174),
            .in3(_gnd_net_),
            .lcout(\ALU.r2_RNI7AQC9_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_LC_9_14_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_LC_9_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_11_s0_c_RNO_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__55527),
            .in2(_gnd_net_),
            .in3(N__34423),
            .lcout(\ALU.r0_12_prm_8_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_12_s0_c_RNO_LC_9_14_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_12_s0_c_RNO_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_12_s0_c_RNO_LC_9_14_6 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \ALU.r0_12_prm_7_12_s0_c_RNO_LC_9_14_6  (
            .in0(N__41358),
            .in1(N__39873),
            .in2(_gnd_net_),
            .in3(N__53193),
            .lcout(\ALU.r0_12_prm_7_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_15_s0_c_RNO_LC_9_14_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_15_s0_c_RNO_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_15_s0_c_RNO_LC_9_14_7 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_15_s0_c_RNO_LC_9_14_7  (
            .in0(N__54606),
            .in1(N__40159),
            .in2(N__53240),
            .in3(N__39993),
            .lcout(\ALU.r0_12_prm_5_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_0_LC_9_15_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_0_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_0_LC_9_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_13_s1_c_RNO_0_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__39889),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\ALU.r0_12_prm_8_13_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s1_c_LC_9_15_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_13_s1_c_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s1_c_LC_9_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_13_s1_c_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__36118),
            .in2(N__36159),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_13_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_13_s1_c_LC_9_15_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_13_s1_c_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_13_s1_c_LC_9_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_13_s1_c_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__31492),
            .in2(N__31477),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_13_s1 ),
            .carryout(\ALU.r0_12_prm_7_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_13_s1_c_LC_9_15_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_13_s1_c_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_13_s1_c_LC_9_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_13_s1_c_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__31444),
            .in2(N__31428),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_13_s1 ),
            .carryout(\ALU.r0_12_prm_6_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_13_s1_c_LC_9_15_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_13_s1_c_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_13_s1_c_LC_9_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_13_s1_c_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__31411),
            .in2(N__31399),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_13_s1 ),
            .carryout(\ALU.r0_12_prm_5_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_13_s1_c_LC_9_15_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_13_s1_c_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_13_s1_c_LC_9_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_13_s1_c_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__31372),
            .in2(N__31360),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_13_s1 ),
            .carryout(\ALU.r0_12_prm_4_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_13_s1_c_LC_9_15_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_13_s1_c_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_13_s1_c_LC_9_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_13_s1_c_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__55263),
            .in2(N__56476),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_13_s1 ),
            .carryout(\ALU.r0_12_prm_3_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_13_s1_c_LC_9_15_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_13_s1_c_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_13_s1_c_LC_9_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_13_s1_c_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__34555),
            .in2(N__34596),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_13_s1 ),
            .carryout(\ALU.r0_12_prm_2_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_13_s1_c_LC_9_16_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_13_s1_c_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_13_s1_c_LC_9_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_13_s1_c_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__35301),
            .in2(N__31504),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\ALU.r0_12_s1_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_13_THRU_LUT4_0_LC_9_16_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_13_THRU_LUT4_0_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_13_THRU_LUT4_0_LC_9_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_13_THRU_LUT4_0_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31516),
            .lcout(\ALU.r0_12_s1_13_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_13_s1_c_RNO_LC_9_16_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_13_s1_c_RNO_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_13_s1_c_RNO_LC_9_16_6 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_13_s1_c_RNO_LC_9_16_6  (
            .in0(N__55957),
            .in1(N__53985),
            .in2(_gnd_net_),
            .in3(N__35300),
            .lcout(\ALU.r0_12_prm_1_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_6_s1_c_RNO_LC_10_1_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_6_s1_c_RNO_LC_10_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_6_s1_c_RNO_LC_10_1_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_6_s1_c_RNO_LC_10_1_0  (
            .in0(_gnd_net_),
            .in1(N__55840),
            .in2(_gnd_net_),
            .in3(N__38257),
            .lcout(\ALU.r0_12_prm_2_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_0_s0_c_RNO_LC_10_1_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_3_0_s0_c_RNO_LC_10_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_0_s0_c_RNO_LC_10_1_1 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_3_0_s0_c_RNO_LC_10_1_1  (
            .in0(N__55221),
            .in1(N__49002),
            .in2(_gnd_net_),
            .in3(N__38031),
            .lcout(\ALU.r0_12_prm_3_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_6_s1_c_RNO_LC_10_1_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_6_s1_c_RNO_LC_10_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_6_s1_c_RNO_LC_10_1_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_7_6_s1_c_RNO_LC_10_1_2  (
            .in0(_gnd_net_),
            .in1(N__53080),
            .in2(_gnd_net_),
            .in3(N__41629),
            .lcout(\ALU.r0_12_prm_7_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_6_s1_c_RNO_LC_10_1_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_6_s1_c_RNO_LC_10_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_6_s1_c_RNO_LC_10_1_5 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_6_s1_c_RNO_LC_10_1_5  (
            .in0(N__43656),
            .in1(N__54894),
            .in2(N__53214),
            .in3(N__43416),
            .lcout(\ALU.r0_12_prm_5_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_RNO_4_LC_10_1_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_2_c_RNO_4_LC_10_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_RNO_4_LC_10_1_6 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r0_12_prm_8_2_c_RNO_4_LC_10_1_6  (
            .in0(N__54032),
            .in1(N__48399),
            .in2(N__54920),
            .in3(N__49398),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_RNO_3_LC_10_1_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_2_c_RNO_3_LC_10_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_RNO_3_LC_10_1_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r0_12_prm_8_2_c_RNO_3_LC_10_1_7  (
            .in0(N__54552),
            .in1(N__45452),
            .in2(N__31495),
            .in3(N__42849),
            .lcout(\ALU.r0_12_prm_8_2_c_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a3_b_3_LC_10_2_1 .C_ON=1'b0;
    defparam \ALU.mult_a3_b_3_LC_10_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a3_b_3_LC_10_2_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.mult_a3_b_3_LC_10_2_1  (
            .in0(N__31936),
            .in1(N__44352),
            .in2(N__32229),
            .in3(N__31839),
            .lcout(\ALU.a3_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a1_b_1_LC_10_2_3 .C_ON=1'b0;
    defparam \ALU.mult_a1_b_1_LC_10_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a1_b_1_LC_10_2_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \ALU.mult_a1_b_1_LC_10_2_3  (
            .in0(N__31664),
            .in1(N__31731),
            .in2(N__32228),
            .in3(N__46798),
            .lcout(\ALU.a1_b_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a1_b_3_LC_10_2_4 .C_ON=1'b0;
    defparam \ALU.mult_a1_b_3_LC_10_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a1_b_3_LC_10_2_4 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \ALU.mult_a1_b_3_LC_10_2_4  (
            .in0(N__44351),
            .in1(N__32178),
            .in2(N__31740),
            .in3(N__31665),
            .lcout(\ALU.a1_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_135_0_LC_10_2_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_135_0_LC_10_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_135_0_LC_10_2_5 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.mult_madd_135_0_LC_10_2_5  (
            .in0(N__40504),
            .in1(N__44350),
            .in2(N__45418),
            .in3(N__43308),
            .lcout(\ALU.madd_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_6_s1_c_RNO_LC_10_2_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_6_s1_c_RNO_LC_10_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_6_s1_c_RNO_LC_10_2_7 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_6_s1_c_RNO_LC_10_2_7  (
            .in0(N__54056),
            .in1(N__43655),
            .in2(N__53215),
            .in3(N__43309),
            .lcout(\ALU.r0_12_prm_6_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_4_c_RNO_0_LC_10_3_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_4_c_RNO_0_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_4_c_RNO_0_LC_10_3_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r0_12_prm_6_4_c_RNO_0_LC_10_3_0  (
            .in0(_gnd_net_),
            .in1(N__42818),
            .in2(_gnd_net_),
            .in3(N__40533),
            .lcout(\ALU.un14_log_0_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIO7CSJ_4_LC_10_3_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIO7CSJ_4_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIO7CSJ_4_LC_10_3_1 .LUT_INIT=16'b1011001110000011;
    LogicCell40 \ALU.r4_RNIO7CSJ_4_LC_10_3_1  (
            .in0(N__42816),
            .in1(N__31540),
            .in2(N__54790),
            .in3(N__49397),
            .lcout(\ALU.r4_RNIO7CSJZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI9H7SJ_5_LC_10_3_2 .C_ON=1'b0;
    defparam \ALU.r4_RNI9H7SJ_5_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI9H7SJ_5_LC_10_3_2 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \ALU.r4_RNI9H7SJ_5_LC_10_3_2  (
            .in0(N__31531),
            .in1(N__45383),
            .in2(N__54800),
            .in3(N__42817),
            .lcout(\ALU.r4_RNI9H7SJZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI8B628_0_5_LC_10_3_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI8B628_0_5_LC_10_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI8B628_0_5_LC_10_3_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.r4_RNI8B628_0_5_LC_10_3_3  (
            .in0(N__45384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45231),
            .lcout(\ALU.r4_RNI8B628_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_0_s0_c_RNO_LC_10_3_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_0_s0_c_RNO_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_0_s0_c_RNO_LC_10_3_4 .LUT_INIT=16'b1010010100001111;
    LogicCell40 \ALU.r0_12_prm_7_0_s0_c_RNO_LC_10_3_4  (
            .in0(N__38026),
            .in1(_gnd_net_),
            .in2(N__53218),
            .in3(N__48935),
            .lcout(\ALU.r0_12_prm_7_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIMVMDA_0_1_LC_10_3_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIMVMDA_0_1_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIMVMDA_0_1_LC_10_3_5 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ALU.r4_RNIMVMDA_0_1_LC_10_3_5  (
            .in0(N__48933),
            .in1(N__53782),
            .in2(N__54791),
            .in3(N__48639),
            .lcout(\ALU.N_622_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_0_s0_c_RNO_LC_10_3_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_0_s0_c_RNO_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_0_s0_c_RNO_LC_10_3_6 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_0_s0_c_RNO_LC_10_3_6  (
            .in0(N__38027),
            .in1(N__54658),
            .in2(N__53219),
            .in3(N__48936),
            .lcout(\ALU.r0_12_prm_5_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_0_s1_c_RNO_LC_10_3_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_0_s1_c_RNO_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_0_s1_c_RNO_LC_10_3_7 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \ALU.r0_12_prm_7_0_s1_c_RNO_LC_10_3_7  (
            .in0(N__48934),
            .in1(N__53091),
            .in2(_gnd_net_),
            .in3(N__38025),
            .lcout(\ALU.r0_12_prm_7_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIUU8UD_3_LC_10_4_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIUU8UD_3_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIUU8UD_3_LC_10_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNIUU8UD_3_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(N__31963),
            .in2(_gnd_net_),
            .in3(N__49324),
            .lcout(\ALU.r4_RNIUU8UDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNINNEH9_0_15_LC_10_4_1 .C_ON=1'b0;
    defparam \ALU.r5_RNINNEH9_0_15_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNINNEH9_0_15_LC_10_4_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ALU.r5_RNINNEH9_0_15_LC_10_4_1  (
            .in0(N__54062),
            .in1(N__40176),
            .in2(N__47070),
            .in3(N__54617),
            .lcout(\ALU.N_845_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKUMQ8_1_8_LC_10_4_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIKUMQ8_1_8_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKUMQ8_1_8_LC_10_4_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \ALU.r4_RNIKUMQ8_1_8_LC_10_4_2  (
            .in0(N__46192),
            .in1(_gnd_net_),
            .in2(N__46446),
            .in3(_gnd_net_),
            .lcout(\ALU.r4_RNIKUMQ8_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a8_b_8_LC_10_4_3 .C_ON=1'b0;
    defparam \ALU.mult_a8_b_8_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a8_b_8_LC_10_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a8_b_8_LC_10_4_3  (
            .in0(_gnd_net_),
            .in1(N__46422),
            .in2(_gnd_net_),
            .in3(N__46191),
            .lcout(\ALU.a8_b_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_490_5_LC_10_4_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_490_5_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_490_5_LC_10_4_4 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_490_5_LC_10_4_4  (
            .in0(N__35594),
            .in1(N__42844),
            .in2(N__45451),
            .in3(N__52003),
            .lcout(\ALU.madd_490_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_RNO_4_LC_10_4_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_3_c_RNO_4_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_RNO_4_LC_10_4_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_12_prm_8_3_c_RNO_4_LC_10_4_5  (
            .in0(N__49325),
            .in1(N__54616),
            .in2(N__42862),
            .in3(N__54055),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_RNO_3_LC_10_4_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_3_c_RNO_3_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_RNO_3_LC_10_4_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r0_12_prm_8_3_c_RNO_3_LC_10_4_6  (
            .in0(N__54618),
            .in1(N__45391),
            .in2(N__32923),
            .in3(N__43415),
            .lcout(),
            .ltout(\ALU.r0_12_prm_8_3_c_RNOZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_RNO_2_LC_10_4_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_3_c_RNO_2_LC_10_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_RNO_2_LC_10_4_7 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.r0_12_prm_8_3_c_RNO_2_LC_10_4_7  (
            .in0(N__50995),
            .in1(N__51442),
            .in2(N__32920),
            .in3(N__32910),
            .lcout(\ALU.rshift_15_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_1_LC_10_5_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_1_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_1_LC_10_5_0 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \ALU.r0_12_prm_8_10_s1_c_RNO_1_LC_10_5_0  (
            .in0(N__38050),
            .in1(N__38075),
            .in2(N__51527),
            .in3(N__50992),
            .lcout(\ALU.r0_12_prm_8_10_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKTVI8_0_4_LC_10_5_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIKTVI8_0_4_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKTVI8_0_4_LC_10_5_1 .LUT_INIT=16'b0101011010011010;
    LogicCell40 \ALU.r4_RNIKTVI8_0_4_LC_10_5_1  (
            .in0(N__40511),
            .in1(N__32224),
            .in2(N__32374),
            .in3(N__32469),
            .lcout(\ALU.un9_addsub_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNITPNQ3_0_LC_10_5_2 .C_ON=1'b0;
    defparam \ALU.r4_RNITPNQ3_0_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNITPNQ3_0_LC_10_5_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.r4_RNITPNQ3_0_LC_10_5_2  (
            .in0(N__32861),
            .in1(N__32752),
            .in2(_gnd_net_),
            .in3(N__32718),
            .lcout(\ALU.b_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIHCHO8_0_2_LC_10_5_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIHCHO8_0_2_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIHCHO8_0_2_LC_10_5_3 .LUT_INIT=16'b0100011110111000;
    LogicCell40 \ALU.r4_RNIHCHO8_0_2_LC_10_5_3  (
            .in0(N__32684),
            .in1(N__32223),
            .in2(N__32592),
            .in3(N__43897),
            .lcout(\ALU.un9_addsub_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKTVI8_4_LC_10_5_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIKTVI8_4_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKTVI8_4_LC_10_5_4 .LUT_INIT=16'b1010110001010011;
    LogicCell40 \ALU.r4_RNIKTVI8_4_LC_10_5_4  (
            .in0(N__32468),
            .in1(N__32360),
            .in2(N__32257),
            .in3(N__40512),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI20C8C_4_LC_10_5_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI20C8C_4_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI20C8C_4_LC_10_5_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.r4_RNI20C8C_4_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31966),
            .in3(N__33882),
            .lcout(\ALU.r4_RNI20C8CZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_1_LC_10_5_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_1_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_1_LC_10_5_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \ALU.r0_12_prm_8_10_s0_c_RNO_1_LC_10_5_6  (
            .in0(N__38051),
            .in1(N__38076),
            .in2(N__51528),
            .in3(N__50993),
            .lcout(\ALU.rshift_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_12_LC_10_5_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_12_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_12_LC_10_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_g0_12_LC_10_5_7  (
            .in0(N__43898),
            .in1(N__44529),
            .in2(N__46217),
            .in3(N__46822),
            .lcout(\ALU.madd_76_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKUMQ8_8_LC_10_6_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIKUMQ8_8_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKUMQ8_8_LC_10_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r4_RNIKUMQ8_8_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__46161),
            .in2(_gnd_net_),
            .in3(N__46412),
            .lcout(\ALU.un14_log_0_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI14AH9_11_LC_10_6_1 .C_ON=1'b0;
    defparam \ALU.r5_RNI14AH9_11_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI14AH9_11_LC_10_6_1 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.r5_RNI14AH9_11_LC_10_6_1  (
            .in0(N__53911),
            .in1(N__51804),
            .in2(N__40989),
            .in3(N__54835),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI1RK3K_9_LC_10_6_2 .C_ON=1'b0;
    defparam \ALU.r4_RNI1RK3K_9_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI1RK3K_9_LC_10_6_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNI1RK3K_9_LC_10_6_2  (
            .in0(N__54836),
            .in1(N__46160),
            .in2(N__32983),
            .in3(N__52255),
            .lcout(\ALU.r4_RNI1RK3KZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIQK1ED_4_LC_10_6_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIQK1ED_4_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIQK1ED_4_LC_10_6_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.r4_RNIQK1ED_4_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32980),
            .in3(N__42838),
            .lcout(\ALU.r4_RNIQK1EDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIVLAIA_9_LC_10_6_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIVLAIA_9_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIVLAIA_9_LC_10_6_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.r4_RNIVLAIA_9_LC_10_6_4  (
            .in0(N__46162),
            .in1(N__53912),
            .in2(_gnd_net_),
            .in3(N__52256),
            .lcout(\ALU.r4_RNIVLAIAZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2H9PK_6_LC_10_6_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI2H9PK_6_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2H9PK_6_LC_10_6_5 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \ALU.r4_RNI2H9PK_6_LC_10_6_5  (
            .in0(N__44588),
            .in1(N__32971),
            .in2(N__43437),
            .in3(N__54837),
            .lcout(\ALU.r4_RNI2H9PKZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_7_s0_c_RNO_LC_10_6_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_7_s0_c_RNO_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_7_s0_c_RNO_LC_10_6_6 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_7_s0_c_RNO_LC_10_6_6  (
            .in0(N__44797),
            .in1(N__53913),
            .in2(N__53220),
            .in3(N__44589),
            .lcout(\ALU.r0_12_prm_6_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIE5LH_1_LC_10_6_7 .C_ON=1'b0;
    defparam \ALU.r0_RNIE5LH_1_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIE5LH_1_LC_10_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.r0_RNIE5LH_1_LC_10_6_7  (
            .in0(N__32954),
            .in1(N__35069),
            .in2(_gnd_net_),
            .in3(N__33174),
            .lcout(\ALU.r0_RNIE5LHZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI50MP_0_LC_10_7_0 .C_ON=1'b0;
    defparam \ALU.r0_RNI50MP_0_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI50MP_0_LC_10_7_0 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ALU.r0_RNI50MP_0_LC_10_7_0  (
            .in0(N__33204),
            .in1(N__33296),
            .in2(N__34853),
            .in3(N__34932),
            .lcout(\ALU.b_3_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b_fast_0_LC_10_7_1.C_ON=1'b0;
    defparam b_fast_0_LC_10_7_1.SEQ_MODE=4'b1000;
    defparam b_fast_0_LC_10_7_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 b_fast_0_LC_10_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33205),
            .lcout(b_fastZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56248),
            .ce(N__56052),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNID8MP_4_LC_10_7_2 .C_ON=1'b0;
    defparam \ALU.r0_RNID8MP_4_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNID8MP_4_LC_10_7_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNID8MP_4_LC_10_7_2  (
            .in0(N__33507),
            .in1(N__33299),
            .in2(N__33468),
            .in3(N__33183),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNISLNE1_4_LC_10_7_3 .C_ON=1'b0;
    defparam \ALU.r4_RNISLNE1_4_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNISLNE1_4_LC_10_7_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNISLNE1_4_LC_10_7_3  (
            .in0(N__33137),
            .in1(N__34289),
            .in2(N__33442),
            .in3(N__33560),
            .lcout(\ALU.r4_RNISLNE1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNI94MP_2_LC_10_7_4 .C_ON=1'b0;
    defparam \ALU.r0_RNI94MP_2_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNI94MP_2_LC_10_7_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNI94MP_2_LC_10_7_4  (
            .in0(N__33411),
            .in1(N__33297),
            .in2(N__33380),
            .in3(N__33181),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKDNE1_2_LC_10_7_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIKDNE1_2_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKDNE1_2_LC_10_7_5 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNIKDNE1_2_LC_10_7_5  (
            .in0(N__33135),
            .in1(N__34329),
            .in2(N__33352),
            .in3(N__33626),
            .lcout(\ALU.r4_RNIKDNE1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_RNIB6MP_3_LC_10_7_6 .C_ON=1'b0;
    defparam \ALU.r0_RNIB6MP_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_RNIB6MP_3_LC_10_7_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.r0_RNIB6MP_3_LC_10_7_6  (
            .in0(N__35042),
            .in1(N__33298),
            .in2(N__33233),
            .in3(N__33182),
            .lcout(),
            .ltout(\ALU.b_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIOHNE1_3_LC_10_7_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIOHNE1_3_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIOHNE1_3_LC_10_7_7 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNIOHNE1_3_LC_10_7_7  (
            .in0(N__33136),
            .in1(N__33064),
            .in2(N__33040),
            .in3(N__33585),
            .lcout(\ALU.r4_RNIOHNE1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_6_LC_10_8_0 .C_ON=1'b0;
    defparam \ALU.r5_6_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_6_LC_10_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_6_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38855),
            .lcout(r5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_7_LC_10_8_1 .C_ON=1'b0;
    defparam \ALU.r5_7_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_7_LC_10_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_7_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38741),
            .lcout(r5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_8_LC_10_8_2 .C_ON=1'b0;
    defparam \ALU.r5_8_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_8_LC_10_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_8_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39513),
            .lcout(r5_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_9_LC_10_8_3 .C_ON=1'b0;
    defparam \ALU.r5_9_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_9_LC_10_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_9_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34022),
            .lcout(r5_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_1_LC_10_8_4 .C_ON=1'b0;
    defparam \ALU.r5_1_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_1_LC_10_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_1_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42139),
            .lcout(r5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_2_LC_10_8_5 .C_ON=1'b0;
    defparam \ALU.r5_2_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_2_LC_10_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_2_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40275),
            .lcout(r5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_3_LC_10_8_6 .C_ON=1'b0;
    defparam \ALU.r5_3_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_3_LC_10_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_3_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50175),
            .lcout(r5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.r5_4_LC_10_8_7 .C_ON=1'b0;
    defparam \ALU.r5_4_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \ALU.r5_4_LC_10_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r5_4_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39062),
            .lcout(r5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(N__45801),
            .sr(_gnd_net_));
    defparam \ALU.mult_a0_b_0_LC_10_9_0 .C_ON=1'b1;
    defparam \ALU.mult_a0_b_0_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a0_b_0_LC_10_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a0_b_0_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__49008),
            .in2(N__40647),
            .in3(N__38015),
            .lcout(\ALU.mult_0 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\ALU.un2_addsub_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_0_c_RNIJPSHD_LC_10_9_1 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_0_c_RNIJPSHD_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_0_c_RNIJPSHD_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_0_c_RNIJPSHD_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__34489),
            .in2(N__33544),
            .in3(N__33964),
            .lcout(\ALU.un2_addsub_cry_0_c_RNIJPSHDZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_0 ),
            .carryout(\ALU.un2_addsub_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_1_c_RNI1H7SG_LC_10_9_2 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_1_c_RNI1H7SG_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_1_c_RNI1H7SG_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_1_c_RNI1H7SG_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__33961),
            .in2(N__33949),
            .in3(N__33925),
            .lcout(\ALU.un2_addsub_cry_1_c_RNI1H7SGZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_1 ),
            .carryout(\ALU.un2_addsub_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_2_c_RNI3K9SG_LC_10_9_3 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_2_c_RNI3K9SG_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_2_c_RNI3K9SG_LC_10_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_2_c_RNI3K9SG_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__33922),
            .in2(N__33910),
            .in3(N__33895),
            .lcout(\ALU.un2_addsub_cry_2_c_RNI3K9SGZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_2 ),
            .carryout(\ALU.un2_addsub_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_3_c_RNI8MVBG_LC_10_9_4 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_3_c_RNI8MVBG_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_3_c_RNI8MVBG_LC_10_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_3_c_RNI8MVBG_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__33892),
            .in2(N__33883),
            .in3(N__33856),
            .lcout(\ALU.un2_addsub_cry_3_c_RNI8MVBGZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_3 ),
            .carryout(\ALU.un2_addsub_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_4_c_RNILPG3D_LC_10_9_5 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_4_c_RNILPG3D_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_4_c_RNILPG3D_LC_10_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_4_c_RNILPG3D_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__45479),
            .in2(N__33853),
            .in3(N__33835),
            .lcout(\ALU.un2_addsub_cry_4_c_RNILPG3DZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_4 ),
            .carryout(\ALU.un2_addsub_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_5_c_RNIO30SD_LC_10_9_6 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_5_c_RNIO30SD_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_5_c_RNIO30SD_LC_10_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_5_c_RNIO30SD_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__43438),
            .in2(N__33832),
            .in3(N__33808),
            .lcout(\ALU.un2_addsub_cry_5_c_RNIO30SDZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_5 ),
            .carryout(\ALU.un2_addsub_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_6_c_RNIPJK8E_LC_10_9_7 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_6_c_RNIPJK8E_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_6_c_RNIPJK8E_LC_10_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_6_c_RNIPJK8E_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__44593),
            .in2(N__40666),
            .in3(N__33805),
            .lcout(\ALU.un2_addsub_cry_6_c_RNIPJK8EZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_6 ),
            .carryout(\ALU.un2_addsub_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_7_c_RNI5ELEE_LC_10_10_0 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_7_c_RNI5ELEE_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_7_c_RNI5ELEE_LC_10_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_7_c_RNI5ELEE_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__46177),
            .in2(N__33802),
            .in3(N__33790),
            .lcout(\ALU.un2_addsub_cry_7_c_RNI5ELEEZ0 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\ALU.un2_addsub_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_8_c_RNINO51F_LC_10_10_1 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_8_c_RNINO51F_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_8_c_RNINO51F_LC_10_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_8_c_RNINO51F_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__52301),
            .in2(N__47287),
            .in3(N__33787),
            .lcout(\ALU.un2_addsub_cry_8_c_RNINO51FZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_8 ),
            .carryout(\ALU.un2_addsub_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_9_c_RNIS67KD_LC_10_10_2 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_9_c_RNIS67KD_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_9_c_RNIS67KD_LC_10_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_9_c_RNIS67KD_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__51716),
            .in2(N__34189),
            .in3(N__34171),
            .lcout(\ALU.un2_addsub_cry_9_c_RNIS67KDZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_9 ),
            .carryout(\ALU.un2_addsub_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_10_c_RNIS4T7D_LC_10_10_3 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_10_c_RNIS4T7D_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_10_c_RNIS4T7D_LC_10_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_10_c_RNIS4T7D_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__40982),
            .in2(N__34168),
            .in3(N__34147),
            .lcout(\ALU.un2_addsub_cry_10_c_RNIS4T7DZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_10 ),
            .carryout(\ALU.un2_addsub_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_11_c_RNICP8AE_LC_10_10_4 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_11_c_RNICP8AE_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_11_c_RNICP8AE_LC_10_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_11_c_RNICP8AE_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__41357),
            .in2(N__34144),
            .in3(N__34132),
            .lcout(\ALU.un2_addsub_cry_11_c_RNICP8AEZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_11 ),
            .carryout(\ALU.un2_addsub_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_12_c_RNI74A7E_LC_10_10_5 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_12_c_RNI74A7E_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_12_c_RNI74A7E_LC_10_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_12_c_RNI74A7E_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__41561),
            .in2(N__34129),
            .in3(N__34111),
            .lcout(\ALU.un2_addsub_cry_12_c_RNI74A7EZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_12 ),
            .carryout(\ALU.un2_addsub_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_13_c_RNIR5I0E_LC_10_10_6 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_13_c_RNIR5I0E_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_13_c_RNIR5I0E_LC_10_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_13_c_RNIR5I0E_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__47040),
            .in2(N__34108),
            .in3(N__34096),
            .lcout(\ALU.un2_addsub_cry_13_c_RNIR5I0EZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_13 ),
            .carryout(\ALU.un2_addsub_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_14_c_RNIHN1F9_LC_10_10_7 .C_ON=1'b0;
    defparam \ALU.un2_addsub_cry_14_c_RNIHN1F9_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_14_c_RNIHN1F9_LC_10_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.un2_addsub_cry_14_c_RNIHN1F9_LC_10_10_7  (
            .in0(N__40154),
            .in1(N__39988),
            .in2(_gnd_net_),
            .in3(N__34093),
            .lcout(\ALU.un2_addsub_cry_14_c_RNIHN1FZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_7_LC_10_11_0 .C_ON=1'b0;
    defparam \ALU.r4_7_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_7_LC_10_11_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r4_7_LC_10_11_0  (
            .in0(N__38747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(N__47787),
            .sr(_gnd_net_));
    defparam \ALU.r4_8_LC_10_11_1 .C_ON=1'b0;
    defparam \ALU.r4_8_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_8_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_8_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39493),
            .lcout(r4_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(N__47787),
            .sr(_gnd_net_));
    defparam \ALU.r4_9_LC_10_11_2 .C_ON=1'b0;
    defparam \ALU.r4_9_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_9_LC_10_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_9_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34014),
            .lcout(r4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(N__47787),
            .sr(_gnd_net_));
    defparam \ALU.r4_1_LC_10_11_3 .C_ON=1'b0;
    defparam \ALU.r4_1_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_1_LC_10_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \ALU.r4_1_LC_10_11_3  (
            .in0(N__42143),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(N__47787),
            .sr(_gnd_net_));
    defparam \ALU.r4_2_LC_10_11_4 .C_ON=1'b0;
    defparam \ALU.r4_2_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_2_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_2_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40289),
            .lcout(r4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(N__47787),
            .sr(_gnd_net_));
    defparam \ALU.r4_4_LC_10_11_5 .C_ON=1'b0;
    defparam \ALU.r4_4_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r4_4_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r4_4_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39082),
            .lcout(r4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(N__47787),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNITS6F71_13_LC_10_12_0 .C_ON=1'b0;
    defparam \ALU.r5_RNITS6F71_13_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNITS6F71_13_LC_10_12_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r5_RNITS6F71_13_LC_10_12_0  (
            .in0(N__51105),
            .in1(N__34258),
            .in2(N__51531),
            .in3(N__34462),
            .lcout(),
            .ltout(\ALU.lshift_15_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI7QTIG2_5_LC_10_12_1 .C_ON=1'b0;
    defparam \ALU.r4_RNI7QTIG2_5_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI7QTIG2_5_LC_10_12_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNI7QTIG2_5_LC_10_12_1  (
            .in0(N__51507),
            .in1(N__50752),
            .in2(N__34237),
            .in3(N__43011),
            .lcout(\ALU.lshift_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_1_LC_10_12_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_1_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s1_c_RNO_1_LC_10_12_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r0_12_prm_8_11_s1_c_RNO_1_LC_10_12_2  (
            .in0(N__51106),
            .in1(N__44889),
            .in2(N__51532),
            .in3(N__44844),
            .lcout(\ALU.r0_12_prm_8_11_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNISP2L9_12_LC_10_12_3 .C_ON=1'b0;
    defparam \ALU.r5_RNISP2L9_12_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNISP2L9_12_LC_10_12_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r5_RNISP2L9_12_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__39860),
            .in2(_gnd_net_),
            .in3(N__41349),
            .lcout(\ALU.un14_log_0_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_11_s0_c_RNO_LC_10_12_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_11_s0_c_RNO_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_11_s0_c_RNO_LC_10_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_11_s0_c_RNO_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__55942),
            .in2(_gnd_net_),
            .in3(N__35833),
            .lcout(\ALU.r0_12_prm_2_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_10_s0_c_RNO_LC_10_12_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_10_s0_c_RNO_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_10_s0_c_RNO_LC_10_12_5 .LUT_INIT=16'b0101000010101111;
    LogicCell40 \ALU.r0_12_prm_1_10_s0_c_RNO_LC_10_12_5  (
            .in0(N__53999),
            .in1(_gnd_net_),
            .in2(N__55961),
            .in3(N__36101),
            .lcout(\ALU.r0_12_prm_1_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_N_884_i_LC_10_12_6 .C_ON=1'b0;
    defparam \ALU.mult_N_884_i_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_N_884_i_LC_10_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.mult_N_884_i_LC_10_12_6  (
            .in0(N__46824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.N_884_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIAP7U9_10_LC_10_12_7 .C_ON=1'b0;
    defparam \ALU.r5_RNIAP7U9_10_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIAP7U9_10_LC_10_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r5_RNIAP7U9_10_LC_10_12_7  (
            .in0(N__53998),
            .in1(N__51825),
            .in2(_gnd_net_),
            .in3(N__52300),
            .lcout(\ALU.r5_RNIAP7U9Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_LC_10_13_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_LC_10_13_0 .LUT_INIT=16'b1110000101001011;
    LogicCell40 \ALU.r0_12_prm_8_12_s0_c_RNO_LC_10_13_0  (
            .in0(N__51473),
            .in1(N__37486),
            .in2(N__55536),
            .in3(N__41029),
            .lcout(\ALU.r0_12_prm_8_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI89OPA_2_LC_10_13_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI89OPA_2_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI89OPA_2_LC_10_13_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r4_RNI89OPA_2_LC_10_13_3  (
            .in0(N__53973),
            .in1(N__48408),
            .in2(N__54781),
            .in3(N__49419),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNII2A0L_1_LC_10_13_4 .C_ON=1'b0;
    defparam \ALU.r4_RNII2A0L_1_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNII2A0L_1_LC_10_13_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNII2A0L_1_LC_10_13_4  (
            .in0(N__54580),
            .in1(N__49017),
            .in2(N__34465),
            .in3(N__48655),
            .lcout(\ALU.r4_RNII2A0LZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIOK1781_9_LC_10_13_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIOK1781_9_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIOK1781_9_LC_10_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r4_RNIOK1781_9_LC_10_13_5  (
            .in0(N__51100),
            .in1(N__34461),
            .in2(_gnd_net_),
            .in3(N__43010),
            .lcout(),
            .ltout(\ALU.r4_RNIOK1781Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI79MLT1_1_LC_10_13_6 .C_ON=1'b0;
    defparam \ALU.r4_RNI79MLT1_1_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI79MLT1_1_LC_10_13_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ALU.r4_RNI79MLT1_1_LC_10_13_6  (
            .in0(N__51472),
            .in1(N__51101),
            .in2(N__34447),
            .in3(N__50740),
            .lcout(\ALU.lshift_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_LC_10_13_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_LC_10_13_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_15_s0_c_RNO_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__55523),
            .in2(_gnd_net_),
            .in3(N__36013),
            .lcout(\ALU.r0_12_prm_8_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_10_s1_c_RNO_LC_10_14_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_10_s1_c_RNO_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_10_s1_c_RNO_LC_10_14_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r0_12_prm_4_10_s1_c_RNO_LC_10_14_0  (
            .in0(N__51829),
            .in1(N__54583),
            .in2(N__54048),
            .in3(N__52992),
            .lcout(\ALU.r0_12_prm_4_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI27VE5_10_LC_10_14_1 .C_ON=1'b0;
    defparam \ALU.r5_RNI27VE5_10_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI27VE5_10_LC_10_14_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r5_RNI27VE5_10_LC_10_14_1  (
            .in0(N__53976),
            .in1(N__54605),
            .in2(N__53165),
            .in3(N__51830),
            .lcout(\ALU.r5_RNI27VE5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_13_s1_c_RNO_LC_10_14_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_13_s1_c_RNO_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_13_s1_c_RNO_LC_10_14_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_2_13_s1_c_RNO_LC_10_14_2  (
            .in0(N__55920),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34579),
            .lcout(\ALU.r0_12_prm_2_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_10_s1_c_RNO_LC_10_14_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_10_s1_c_RNO_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_10_s1_c_RNO_LC_10_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_10_s1_c_RNO_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__55919),
            .in2(_gnd_net_),
            .in3(N__35636),
            .lcout(\ALU.r0_12_prm_2_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_10_s1_c_RNO_LC_10_14_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_10_s1_c_RNO_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_10_s1_c_RNO_LC_10_14_5 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_10_s1_c_RNO_LC_10_14_5  (
            .in0(N__53975),
            .in1(N__52001),
            .in2(N__53164),
            .in3(N__51828),
            .lcout(\ALU.r0_12_prm_6_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_1_LC_10_14_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_1_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_1_LC_10_14_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.r0_12_prm_8_15_s0_c_RNO_1_LC_10_14_6  (
            .in0(N__54604),
            .in1(N__53974),
            .in2(N__50707),
            .in3(N__40155),
            .lcout(\ALU.rshift_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_1_LC_10_14_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_1_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_11_s0_c_RNO_1_LC_10_14_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r0_12_prm_8_11_s0_c_RNO_1_LC_10_14_7  (
            .in0(N__51104),
            .in1(N__44888),
            .in2(N__51541),
            .in3(N__44843),
            .lcout(\ALU.rshift_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_0_LC_10_15_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_0_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_0_LC_10_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_10_s1_c_RNO_0_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__34534),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\ALU.r0_12_prm_8_10_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s1_c_LC_10_15_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_10_s1_c_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s1_c_LC_10_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_10_s1_c_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__42256),
            .in2(N__42346),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_10_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_10_s1_c_LC_10_15_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_10_s1_c_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_10_s1_c_LC_10_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_10_s1_c_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__34522),
            .in2(N__34512),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_10_s1 ),
            .carryout(\ALU.r0_12_prm_7_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_10_s1_c_LC_10_15_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_10_s1_c_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_10_s1_c_LC_10_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_10_s1_c_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__34744),
            .in2(N__34738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_10_s1 ),
            .carryout(\ALU.r0_12_prm_6_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_10_s1_c_LC_10_15_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_10_s1_c_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_10_s1_c_LC_10_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_10_s1_c_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__34711),
            .in2(N__34705),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_10_s1 ),
            .carryout(\ALU.r0_12_prm_5_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_10_s1_c_LC_10_15_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_10_s1_c_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_10_s1_c_LC_10_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_10_s1_c_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__34681),
            .in2(N__34675),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_10_s1 ),
            .carryout(\ALU.r0_12_prm_4_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_10_s1_c_LC_10_15_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_10_s1_c_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_10_s1_c_LC_10_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_10_s1_c_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__55264),
            .in2(N__56477),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_10_s1 ),
            .carryout(\ALU.r0_12_prm_3_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_10_s1_c_LC_10_15_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_10_s1_c_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_10_s1_c_LC_10_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_10_s1_c_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__35637),
            .in2(N__34651),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_10_s1 ),
            .carryout(\ALU.r0_12_prm_2_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_10_s1_c_LC_10_16_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_10_s1_c_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_10_s1_c_LC_10_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_10_s1_c_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__36108),
            .in2(N__36073),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\ALU.r0_12_s1_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_10_THRU_LUT4_0_LC_10_16_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_10_THRU_LUT4_0_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_10_THRU_LUT4_0_LC_10_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_10_THRU_LUT4_0_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34642),
            .lcout(\ALU.r0_12_s1_10_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_13_s0_c_RNO_LC_10_16_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_13_s0_c_RNO_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_13_s0_c_RNO_LC_10_16_3 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_13_s0_c_RNO_LC_10_16_3  (
            .in0(N__55958),
            .in1(N__53986),
            .in2(_gnd_net_),
            .in3(N__35296),
            .lcout(\ALU.r0_12_prm_1_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_6_s1_c_THRU_CRY_0_LC_11_1_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_6_s1_c_THRU_CRY_0_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_6_s1_c_THRU_CRY_0_LC_11_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_6_s1_c_THRU_CRY_0_LC_11_1_0  (
            .in0(_gnd_net_),
            .in1(N__37726),
            .in2(N__37734),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(\ALU.r0_12_prm_8_6_s1_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_6_s1_c_LC_11_1_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_6_s1_c_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_6_s1_c_LC_11_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_6_s1_c_LC_11_1_1  (
            .in0(_gnd_net_),
            .in1(N__34819),
            .in2(N__37689),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_6_s1_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_6_s1_c_LC_11_1_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_6_s1_c_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_6_s1_c_LC_11_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_6_s1_c_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(N__41642),
            .in2(N__34789),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_6_s1 ),
            .carryout(\ALU.r0_12_prm_7_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_6_s1_c_LC_11_1_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_6_s1_c_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_6_s1_c_LC_11_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_6_s1_c_LC_11_1_3  (
            .in0(_gnd_net_),
            .in1(N__34780),
            .in2(N__38361),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_6_s1 ),
            .carryout(\ALU.r0_12_prm_6_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_6_s1_c_LC_11_1_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_6_s1_c_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_6_s1_c_LC_11_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_6_s1_c_LC_11_1_4  (
            .in0(_gnd_net_),
            .in1(N__34774),
            .in2(N__38340),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_6_s1 ),
            .carryout(\ALU.r0_12_prm_5_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_6_s1_c_LC_11_1_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_6_s1_c_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_6_s1_c_LC_11_1_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_6_s1_c_LC_11_1_5  (
            .in0(_gnd_net_),
            .in1(N__34765),
            .in2(N__38296),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_6_s1 ),
            .carryout(\ALU.r0_12_prm_4_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_6_s1_c_LC_11_1_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_6_s1_c_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_6_s1_c_LC_11_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_6_s1_c_LC_11_1_6  (
            .in0(_gnd_net_),
            .in1(N__55222),
            .in2(N__56512),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_6_s1 ),
            .carryout(\ALU.r0_12_prm_3_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_6_s1_c_LC_11_1_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_6_s1_c_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_6_s1_c_LC_11_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_6_s1_c_LC_11_1_7  (
            .in0(_gnd_net_),
            .in1(N__38266),
            .in2(N__34753),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_6_s1 ),
            .carryout(\ALU.r0_12_prm_2_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_6_s1_c_LC_11_2_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_6_s1_c_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_6_s1_c_LC_11_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_6_s1_c_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__38204),
            .in2(N__36358),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\ALU.r0_12_s1_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_6_THRU_LUT4_0_LC_11_2_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_6_THRU_LUT4_0_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_6_THRU_LUT4_0_LC_11_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_6_THRU_LUT4_0_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34825),
            .lcout(\ALU.r0_12_s1_6_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIAP9541_4_LC_11_2_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIAP9541_4_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIAP9541_4_LC_11_2_2 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ALU.r4_RNIAP9541_4_LC_11_2_2  (
            .in0(N__50994),
            .in1(N__42222),
            .in2(N__51483),
            .in3(N__42205),
            .lcout(\ALU.lshift_6 ),
            .ltout(\ALU.lshift_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_6_s1_c_RNO_LC_11_2_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_6_s1_c_RNO_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_6_s1_c_RNO_LC_11_2_3 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \ALU.r0_12_prm_8_6_s1_c_RNO_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34822),
            .in3(N__55458),
            .lcout(\ALU.r0_12_prm_8_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2BKQ8_0_6_LC_11_2_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI2BKQ8_0_6_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2BKQ8_0_6_LC_11_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNI2BKQ8_0_6_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__43657),
            .in2(_gnd_net_),
            .in3(N__43403),
            .lcout(\ALU.r4_RNI2BKQ8_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIUGHG5_6_LC_11_2_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIUGHG5_6_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIUGHG5_6_LC_11_2_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r4_RNIUGHG5_6_LC_11_2_5  (
            .in0(N__43404),
            .in1(N__54783),
            .in2(N__53152),
            .in3(N__54036),
            .lcout(\ALU.r4_RNIUGHG5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI5OTIG2_2_LC_11_2_6 .C_ON=1'b0;
    defparam \ALU.r4_RNI5OTIG2_2_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI5OTIG2_2_LC_11_2_6 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \ALU.r4_RNI5OTIG2_2_LC_11_2_6  (
            .in0(N__36376),
            .in1(N__41098),
            .in2(N__51484),
            .in3(N__41707),
            .lcout(\ALU.rshift_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNID26E8_1_0_LC_11_2_7 .C_ON=1'b0;
    defparam \ALU.r4_RNID26E8_1_0_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNID26E8_1_0_LC_11_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNID26E8_1_0_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(N__49001),
            .in2(_gnd_net_),
            .in3(N__38016),
            .lcout(\ALU.un9_addsub_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_0_s0_c_LC_11_3_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_0_s0_c_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_0_s0_c_LC_11_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_0_s0_c_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__40704),
            .in2(N__40198),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\ALU.r0_12_prm_8_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_0_s0_c_LC_11_3_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_0_s0_c_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_0_s0_c_LC_11_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_0_s0_c_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__36439),
            .in2(N__34813),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_0_s0 ),
            .carryout(\ALU.r0_12_prm_7_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_0_s0_c_LC_11_3_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_0_s0_c_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_0_s0_c_LC_11_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_0_s0_c_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__36312),
            .in2(N__34801),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_0_s0 ),
            .carryout(\ALU.r0_12_prm_6_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_0_s0_c_LC_11_3_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_0_s0_c_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_0_s0_c_LC_11_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_0_s0_c_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__37756),
            .in2(N__34921),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_0_s0 ),
            .carryout(\ALU.r0_12_prm_5_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_0_s0_c_inv_LC_11_3_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_0_s0_c_inv_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_0_s0_c_inv_LC_11_3_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_0_s0_c_inv_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__36279),
            .in2(N__34912),
            .in3(N__48909),
            .lcout(\ALU.N_883_i ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_0_s0 ),
            .carryout(\ALU.r0_12_prm_4_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_0_s0_c_LC_11_3_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_0_s0_c_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_0_s0_c_LC_11_3_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_0_s0_c_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(N__36440),
            .in2(N__34894),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_0_s0 ),
            .carryout(\ALU.r0_12_prm_3_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_0_s0_c_LC_11_3_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_0_s0_c_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_0_s0_c_LC_11_3_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_0_s0_c_LC_11_3_6  (
            .in0(_gnd_net_),
            .in1(N__40617),
            .in2(N__36367),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_0_s0 ),
            .carryout(\ALU.r0_12_prm_2_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_0_s0_c_LC_11_3_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_0_s0_c_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_0_s0_c_LC_11_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_0_s0_c_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(N__36399),
            .in2(N__34882),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_2_0_s0 ),
            .carryout(\ALU.r0_12_s0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_0_s0_c_RNIGKQLG2_LC_11_4_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_0_s0_c_RNIGKQLG2_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_0_s0_c_RNIGKQLG2_LC_11_4_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r0_12_prm_1_0_s0_c_RNIGKQLG2_LC_11_4_0  (
            .in0(N__36382),
            .in1(N__34867),
            .in2(_gnd_net_),
            .in3(N__34858),
            .lcout(\ALU.r0_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_0_LC_11_4_1 .C_ON=1'b0;
    defparam \ALU.r1_0_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_0_LC_11_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_0_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34970),
            .lcout(r1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56234),
            .ce(N__47576),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIRCFPA_7_LC_11_5_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIRCFPA_7_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIRCFPA_7_LC_11_5_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r4_RNIRCFPA_7_LC_11_5_0  (
            .in0(N__53872),
            .in1(N__46199),
            .in2(N__54888),
            .in3(N__44530),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIODO6K_5_LC_11_5_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIODO6K_5_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIODO6K_5_LC_11_5_1 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.r4_RNIODO6K_5_LC_11_5_1  (
            .in0(N__43379),
            .in1(N__54821),
            .in2(N__35101),
            .in3(N__45484),
            .lcout(\ALU.r4_RNIODO6KZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNILIPV9_6_LC_11_5_2 .C_ON=1'b0;
    defparam \ALU.r4_RNILIPV9_6_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNILIPV9_6_LC_11_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r4_RNILIPV9_6_LC_11_5_2  (
            .in0(N__53873),
            .in1(N__43380),
            .in2(_gnd_net_),
            .in3(N__44531),
            .lcout(),
            .ltout(\ALU.r4_RNILIPV9Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI1G9PK_6_LC_11_5_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI1G9PK_6_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI1G9PK_6_LC_11_5_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.r4_RNI1G9PK_6_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__54822),
            .in2(N__35098),
            .in3(N__38631),
            .lcout(\ALU.r4_RNI1G9PKZ0Z_6 ),
            .ltout(\ALU.r4_RNI1G9PKZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNICUATH1_15_LC_11_5_4 .C_ON=1'b0;
    defparam \ALU.r5_RNICUATH1_15_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNICUATH1_15_LC_11_5_4 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \ALU.r5_RNICUATH1_15_LC_11_5_4  (
            .in0(N__36835),
            .in1(N__51423),
            .in2(N__35095),
            .in3(N__38052),
            .lcout(\ALU.rshift_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJTDS9_5_LC_11_5_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIJTDS9_5_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJTDS9_5_LC_11_5_5 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r4_RNIJTDS9_5_LC_11_5_5  (
            .in0(N__53871),
            .in1(N__45483),
            .in2(N__54887),
            .in3(N__42837),
            .lcout(\ALU.lshift_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_5_s0_c_RNO_LC_11_5_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_5_s0_c_RNO_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_5_s0_c_RNO_LC_11_5_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_5_s0_c_RNO_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__55941),
            .in2(_gnd_net_),
            .in3(N__45686),
            .lcout(\ALU.r0_12_prm_2_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI8R2TI_11_LC_11_5_7 .C_ON=1'b0;
    defparam \ALU.r5_RNI8R2TI_11_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI8R2TI_11_LC_11_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r5_RNI8R2TI_11_LC_11_5_7  (
            .in0(N__54817),
            .in1(N__38649),
            .in2(_gnd_net_),
            .in3(N__41728),
            .lcout(\ALU.r5_RNI8R2TIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_1_LC_11_6_0 .C_ON=1'b0;
    defparam \ALU.r0_1_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_1_LC_11_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_1_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42154),
            .lcout(r0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56240),
            .ce(N__49685),
            .sr(_gnd_net_));
    defparam \ALU.r0_3_LC_11_6_1 .C_ON=1'b0;
    defparam \ALU.r0_3_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_3_LC_11_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_3_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50136),
            .lcout(r0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56240),
            .ce(N__49685),
            .sr(_gnd_net_));
    defparam \ALU.r0_0_LC_11_6_6 .C_ON=1'b0;
    defparam \ALU.r0_0_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_0_LC_11_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_0_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34986),
            .lcout(r0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56240),
            .ce(N__49685),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI9S2TI_11_LC_11_7_0 .C_ON=1'b0;
    defparam \ALU.r5_RNI9S2TI_11_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI9S2TI_11_LC_11_7_0 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.r5_RNI9S2TI_11_LC_11_7_0  (
            .in0(N__35665),
            .in1(N__51815),
            .in2(N__54638),
            .in3(N__40991),
            .lcout(),
            .ltout(\ALU.r5_RNI9S2TIZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI8VM481_11_LC_11_7_1 .C_ON=1'b0;
    defparam \ALU.r5_RNI8VM481_11_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI8VM481_11_LC_11_7_1 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.r5_RNI8VM481_11_LC_11_7_1  (
            .in0(N__51474),
            .in1(N__51047),
            .in2(N__35164),
            .in3(N__36867),
            .lcout(),
            .ltout(\ALU.lshift_15_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIS8K872_2_LC_11_7_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIS8K872_2_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIS8K872_2_LC_11_7_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r4_RNIS8K872_2_LC_11_7_2  (
            .in0(N__51475),
            .in1(N__46493),
            .in2(N__35161),
            .in3(N__44827),
            .lcout(\ALU.lshift_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIKS4A9_11_LC_11_7_3 .C_ON=1'b0;
    defparam \ALU.r5_RNIKS4A9_11_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIKS4A9_11_LC_11_7_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.r5_RNIKS4A9_11_LC_11_7_3  (
            .in0(N__40990),
            .in1(_gnd_net_),
            .in2(N__51838),
            .in3(N__53644),
            .lcout(\ALU.r5_RNIKS4A9Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI468UD_2_LC_11_7_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI468UD_2_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI468UD_2_LC_11_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNI468UD_2_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__35158),
            .in2(_gnd_net_),
            .in3(N__48395),
            .lcout(\ALU.r4_RNI468UDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_7_s0_c_RNO_LC_11_7_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_7_s0_c_RNO_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_7_s0_c_RNO_LC_11_7_5 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_7_s0_c_RNO_LC_11_7_5  (
            .in0(N__55808),
            .in1(N__53646),
            .in2(_gnd_net_),
            .in3(N__45001),
            .lcout(\ALU.r0_12_prm_1_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_6_s0_c_RNO_LC_11_7_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_6_s0_c_RNO_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_6_s0_c_RNO_LC_11_7_6 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \ALU.r0_12_prm_1_6_s0_c_RNO_LC_11_7_6  (
            .in0(N__53645),
            .in1(N__55807),
            .in2(_gnd_net_),
            .in3(N__38185),
            .lcout(\ALU.r0_12_prm_1_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIE0AK8_11_LC_11_7_7 .C_ON=1'b0;
    defparam \ALU.r5_RNIE0AK8_11_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIE0AK8_11_LC_11_7_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ALU.r5_RNIE0AK8_11_LC_11_7_7  (
            .in0(N__40992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35605),
            .lcout(\ALU.un14_log_0_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a6_b_0_LC_11_8_0 .C_ON=1'b1;
    defparam \ALU.mult_a6_b_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a6_b_0_LC_11_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_a6_b_0_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__37960),
            .in2(N__49018),
            .in3(N__43377),
            .lcout(\ALU.a6_b_0 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\ALU.un9_addsub_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_0_c_RNIG8GLJ_LC_11_8_1 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_0_c_RNIG8GLJ_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_0_c_RNIG8GLJ_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_0_c_RNIG8GLJ_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__48638),
            .in2(N__35239),
            .in3(N__35221),
            .lcout(\ALU.un9_addsub_cry_0_c_RNIG8GLJZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_0 ),
            .carryout(\ALU.un9_addsub_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_1_c_RNIKO6AJ_LC_11_8_2 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_1_c_RNIKO6AJ_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_1_c_RNIKO6AJ_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_1_c_RNIKO6AJ_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__35218),
            .in2(N__48409),
            .in3(N__35212),
            .lcout(\ALU.un9_addsub_cry_1_c_RNIKO6AJZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_1 ),
            .carryout(\ALU.un9_addsub_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_2_c_RNIOR8AJ_LC_11_8_3 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_2_c_RNIOR8AJ_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_2_c_RNIOR8AJ_LC_11_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_2_c_RNIOR8AJ_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__49424),
            .in2(N__35209),
            .in3(N__35194),
            .lcout(\ALU.un9_addsub_cry_2_c_RNIOR8AJZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_2 ),
            .carryout(\ALU.un9_addsub_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_3_c_RNIV8DFI_LC_11_8_4 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_3_c_RNIV8DFI_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_3_c_RNIV8DFI_LC_11_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_3_c_RNIV8DFI_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__35191),
            .in2(N__42868),
            .in3(N__35182),
            .lcout(\ALU.un9_addsub_cry_3_c_RNIV8DFIZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_3 ),
            .carryout(\ALU.un9_addsub_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_4_c_RNI8AH88_LC_11_8_5 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_4_c_RNI8AH88_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_4_c_RNI8AH88_LC_11_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_4_c_RNI8AH88_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__45250),
            .in2(N__45514),
            .in3(N__35179),
            .lcout(\ALU.un9_addsub_cry_4_c_RNI8AHZ0Z88 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_4 ),
            .carryout(\ALU.un9_addsub_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_5_c_RNI3C019_LC_11_8_6 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_5_c_RNI3C019_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_5_c_RNI3C019_LC_11_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_5_c_RNI3C019_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__43378),
            .in2(N__43667),
            .in3(N__35176),
            .lcout(\ALU.un9_addsub_cry_5_c_RNI3CZ0Z019 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_5 ),
            .carryout(\ALU.un9_addsub_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_6_c_RNIJH4R8_LC_11_8_7 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_6_c_RNIJH4R8_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_6_c_RNIJH4R8_LC_11_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_6_c_RNIJH4R8_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__44594),
            .in2(N__44806),
            .in3(N__35173),
            .lcout(\ALU.un9_addsub_cry_6_c_RNIJH4RZ0Z8 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_6 ),
            .carryout(\ALU.un9_addsub_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_7_c_RNIN3519_LC_11_9_0 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_7_c_RNIN3519_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_7_c_RNIN3519_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_7_c_RNIN3519_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__46200),
            .in2(N__46461),
            .in3(N__35170),
            .lcout(\ALU.un9_addsub_cry_7_c_RNINZ0Z3519 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\ALU.un9_addsub_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_8_c_RNI06LJ9_LC_11_9_1 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_8_c_RNI06LJ9_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_8_c_RNI06LJ9_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_8_c_RNI06LJ9_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__52293),
            .in2(N__47475),
            .in3(N__35167),
            .lcout(\ALU.un9_addsub_cry_8_c_RNI06LJZ0Z9 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_8 ),
            .carryout(\ALU.un9_addsub_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_9_c_RNI3PPQ8_LC_11_9_2 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_9_c_RNI3PPQ8_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_9_c_RNI3PPQ8_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_9_c_RNI3PPQ8_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__51795),
            .in2(N__52029),
            .in3(N__35608),
            .lcout(\ALU.un9_addsub_cry_9_c_RNI3PPQZ0Z8 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_9 ),
            .carryout(\ALU.un9_addsub_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_10_c_RNIRLO09_LC_11_9_3 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_10_c_RNIRLO09_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_10_c_RNIRLO09_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_10_c_RNIRLO09_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__40911),
            .in2(N__35604),
            .in3(N__35434),
            .lcout(\ALU.un9_addsub_cry_10_c_RNIRLOZ0Z09 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_10 ),
            .carryout(\ALU.un9_addsub_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_11_c_RNIAHI1A_LC_11_9_4 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_11_c_RNIAHI1A_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_11_c_RNIAHI1A_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_11_c_RNIAHI1A_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__41356),
            .in2(N__39875),
            .in3(N__35431),
            .lcout(\ALU.un9_addsub_cry_11_c_RNIAHI1AZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_11 ),
            .carryout(\ALU.un9_addsub_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_12_c_RNISR30A_LC_11_9_5 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_12_c_RNISR30A_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_12_c_RNISR30A_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_12_c_RNISR30A_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__41571),
            .in2(N__35424),
            .in3(N__35266),
            .lcout(\ALU.un9_addsub_cry_12_c_RNISR30AZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_12 ),
            .carryout(\ALU.un9_addsub_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_13_c_RNI7LBP9_LC_11_9_6 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_13_c_RNI7LBP9_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_13_c_RNI7LBP9_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_13_c_RNI7LBP9_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__47056),
            .in2(N__47182),
            .in3(N__35263),
            .lcout(\ALU.un9_addsub_cry_13_c_RNI7LBPZ0Z9 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_13 ),
            .carryout(\ALU.un9_addsub_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_14_c_RNIO7DP9_LC_11_9_7 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_14_c_RNIO7DP9_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_14_c_RNIO7DP9_LC_11_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.un9_addsub_cry_14_c_RNIO7DP9_LC_11_9_7  (
            .in0(N__40173),
            .in1(N__39981),
            .in2(_gnd_net_),
            .in3(N__35260),
            .lcout(\ALU.un9_addsub_cry_14_c_RNIO7DPZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_10_s0_c_RNO_LC_11_10_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_10_s0_c_RNO_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_10_s0_c_RNO_LC_11_10_0 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_10_s0_c_RNO_LC_11_10_0  (
            .in0(N__52034),
            .in1(N__53895),
            .in2(N__53236),
            .in3(N__51796),
            .lcout(\ALU.r0_12_prm_6_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_15_s0_c_RNO_LC_11_10_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_15_s0_c_RNO_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_15_s0_c_RNO_LC_11_10_2 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_15_s0_c_RNO_LC_11_10_2  (
            .in0(N__55861),
            .in1(N__53894),
            .in2(_gnd_net_),
            .in3(N__37273),
            .lcout(\ALU.r0_12_prm_1_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_14_s1_c_RNO_LC_11_10_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_14_s1_c_RNO_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_14_s1_c_RNO_LC_11_10_3 .LUT_INIT=16'b0101000010101111;
    LogicCell40 \ALU.r0_12_prm_1_14_s1_c_RNO_LC_11_10_3  (
            .in0(N__53893),
            .in1(_gnd_net_),
            .in2(N__55847),
            .in3(N__49054),
            .lcout(\ALU.r0_12_prm_1_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_8_s1_c_RNO_LC_11_10_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_8_s1_c_RNO_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_8_s1_c_RNO_LC_11_10_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_8_s1_c_RNO_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__55776),
            .in2(_gnd_net_),
            .in3(N__39391),
            .lcout(\ALU.r0_12_prm_2_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_12_s1_c_RNO_LC_11_10_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_12_s1_c_RNO_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_12_s1_c_RNO_LC_11_10_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_12_s1_c_RNO_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__55772),
            .in2(_gnd_net_),
            .in3(N__37636),
            .lcout(\ALU.r0_12_prm_2_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_3_c_RNO_0_LC_11_10_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_3_c_RNO_0_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_3_c_RNO_0_LC_11_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r0_12_prm_6_3_c_RNO_0_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__49423),
            .in2(_gnd_net_),
            .in3(N__44365),
            .lcout(\ALU.un14_log_0_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_LC_11_11_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_LC_11_11_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_13_s0_c_RNO_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__55521),
            .in2(_gnd_net_),
            .in3(N__36141),
            .lcout(\ALU.r0_12_prm_8_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_12_s0_c_RNO_LC_11_11_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_12_s0_c_RNO_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_12_s0_c_RNO_LC_11_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_12_s0_c_RNO_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__55930),
            .in2(_gnd_net_),
            .in3(N__37637),
            .lcout(\ALU.r0_12_prm_2_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_9_s0_c_RNO_LC_11_11_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_9_s0_c_RNO_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_9_s0_c_RNO_LC_11_11_2 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_9_s0_c_RNO_LC_11_11_2  (
            .in0(N__55931),
            .in1(N__53780),
            .in2(_gnd_net_),
            .in3(N__42391),
            .lcout(\ALU.r0_12_prm_1_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIKUTI9_13_LC_11_11_3 .C_ON=1'b0;
    defparam \ALU.r5_RNIKUTI9_13_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIKUTI9_13_LC_11_11_3 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r5_RNIKUTI9_13_LC_11_11_3  (
            .in0(N__53778),
            .in1(N__41555),
            .in2(N__54607),
            .in3(N__41301),
            .lcout(\ALU.lshift_3_ns_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_15_s0_c_RNO_LC_11_11_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_15_s0_c_RNO_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_15_s0_c_RNO_LC_11_11_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_2_15_s0_c_RNO_LC_11_11_4  (
            .in0(N__55928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36235),
            .lcout(\ALU.r0_12_prm_2_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_1_LC_11_11_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_1_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s0_c_RNO_1_LC_11_11_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \ALU.r0_12_prm_8_12_s0_c_RNO_1_LC_11_11_5  (
            .in0(N__51103),
            .in1(_gnd_net_),
            .in2(N__51537),
            .in3(N__41706),
            .lcout(\ALU.rshift_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_10_s0_c_RNO_LC_11_11_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_10_s0_c_RNO_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_10_s0_c_RNO_LC_11_11_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_2_10_s0_c_RNO_LC_11_11_6  (
            .in0(N__55929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35632),
            .lcout(\ALU.r0_12_prm_2_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_12_s1_c_RNO_LC_11_11_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_12_s1_c_RNO_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_12_s1_c_RNO_LC_11_11_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_12_s1_c_RNO_LC_11_11_7  (
            .in0(N__53779),
            .in1(N__54447),
            .in2(N__53104),
            .in3(N__41302),
            .lcout(\ALU.r0_12_prm_4_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_11_s1_c_RNO_LC_11_12_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_11_s1_c_RNO_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_11_s1_c_RNO_LC_11_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_11_s1_c_RNO_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__55933),
            .in2(_gnd_net_),
            .in3(N__35834),
            .lcout(\ALU.r0_12_prm_2_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_1_c_RNO_LC_11_12_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_1_c_RNO_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_1_c_RNO_LC_11_12_1 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_1_c_RNO_LC_11_12_1  (
            .in0(N__54860),
            .in1(N__48652),
            .in2(N__53221),
            .in3(N__46831),
            .lcout(\ALU.r0_12_prm_5_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_12_s1_c_RNO_LC_11_12_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_12_s1_c_RNO_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_12_s1_c_RNO_LC_11_12_2 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \ALU.r0_12_prm_1_12_s1_c_RNO_LC_11_12_2  (
            .in0(N__54001),
            .in1(N__55932),
            .in2(_gnd_net_),
            .in3(N__37576),
            .lcout(\ALU.r0_12_prm_1_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIKU3HJ_10_LC_11_12_3 .C_ON=1'b0;
    defparam \ALU.r5_RNIKU3HJ_10_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIKU3HJ_10_LC_11_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r5_RNIKU3HJ_10_LC_11_12_3  (
            .in0(N__54859),
            .in1(N__39358),
            .in2(_gnd_net_),
            .in3(N__35785),
            .lcout(),
            .ltout(\ALU.r5_RNIKU3HJZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIQK1V71_5_LC_11_12_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIQK1V71_5_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIQK1V71_5_LC_11_12_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.r4_RNIQK1V71_5_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__51089),
            .in2(N__35779),
            .in3(N__38943),
            .lcout(\ALU.r4_RNIQK1V71Z0Z_5 ),
            .ltout(\ALU.r4_RNIQK1V71Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI8E2N22_2_LC_11_12_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI8E2N22_2_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI8E2N22_2_LC_11_12_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.r4_RNI8E2N22_2_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__51523),
            .in2(N__35776),
            .in3(N__41025),
            .lcout(\ALU.lshift_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_11_s0_c_RNO_LC_11_12_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_11_s0_c_RNO_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_11_s0_c_RNO_LC_11_12_7 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \ALU.r0_12_prm_1_11_s0_c_RNO_LC_11_12_7  (
            .in0(N__35748),
            .in1(N__55946),
            .in2(_gnd_net_),
            .in3(N__54000),
            .lcout(\ALU.r0_12_prm_1_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINPPC9_14_LC_11_13_1 .C_ON=1'b0;
    defparam \ALU.r2_RNINPPC9_14_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINPPC9_14_LC_11_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r2_RNINPPC9_14_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__47194),
            .in2(_gnd_net_),
            .in3(N__47032),
            .lcout(\ALU.un14_log_0_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI5P1F5_15_LC_11_13_2 .C_ON=1'b0;
    defparam \ALU.r5_RNI5P1F5_15_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI5P1F5_15_LC_11_13_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r5_RNI5P1F5_15_LC_11_13_2  (
            .in0(N__54611),
            .in1(N__54024),
            .in2(N__53222),
            .in3(N__40106),
            .lcout(\ALU.r5_RNI5P1F5Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_14_s0_c_RNO_LC_11_13_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_14_s0_c_RNO_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_14_s0_c_RNO_LC_11_13_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_14_s0_c_RNO_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__55939),
            .in2(_gnd_net_),
            .in3(N__49132),
            .lcout(\ALU.r0_12_prm_2_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_0_LC_11_14_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s0_c_RNO_0_LC_11_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_15_s0_c_RNO_0_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__36037),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\ALU.r0_12_prm_8_15_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s0_c_LC_11_14_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_15_s0_c_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s0_c_LC_11_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_15_s0_c_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__36027),
            .in2(N__35995),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_15_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_15_s0_c_LC_11_14_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_15_s0_c_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_15_s0_c_LC_11_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_15_s0_c_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__39898),
            .in2(N__35982),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_15_s0 ),
            .carryout(\ALU.r0_12_prm_7_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_15_s0_c_LC_11_14_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_15_s0_c_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_15_s0_c_LC_11_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_15_s0_c_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__35962),
            .in2(N__35953),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_15_s0 ),
            .carryout(\ALU.r0_12_prm_6_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_15_s0_c_LC_11_14_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_15_s0_c_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_15_s0_c_LC_11_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_15_s0_c_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__35920),
            .in2(N__35910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_15_s0 ),
            .carryout(\ALU.r0_12_prm_5_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_15_s0_c_inv_LC_11_14_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_15_s0_c_inv_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_15_s0_c_inv_LC_11_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_15_s0_c_inv_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__35887),
            .in2(N__35874),
            .in3(N__40156),
            .lcout(\ALU.a_i_15 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_15_s0 ),
            .carryout(\ALU.r0_12_prm_4_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_15_s0_c_inv_LC_11_14_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_15_s0_c_inv_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_15_s0_c_inv_LC_11_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_3_15_s0_c_inv_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__36265),
            .in2(_gnd_net_),
            .in3(N__55234),
            .lcout(\ALU.r0_12_prm_3_15_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_15_s0 ),
            .carryout(\ALU.r0_12_prm_3_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_15_s0_c_LC_11_14_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_15_s0_c_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_15_s0_c_LC_11_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_15_s0_c_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__36252),
            .in2(N__36214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_15_s0 ),
            .carryout(\ALU.r0_12_prm_2_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_15_s0_c_LC_11_15_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_15_s0_c_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_15_s0_c_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_15_s0_c_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__36202),
            .in2(N__37290),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\ALU.r0_12_s0_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s0_15_THRU_LUT4_0_LC_11_15_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s0_15_THRU_LUT4_0_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s0_15_THRU_LUT4_0_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s0_15_THRU_LUT4_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36193),
            .lcout(\ALU.r0_12_s0_15_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIB8HG5_12_LC_11_15_5 .C_ON=1'b0;
    defparam \ALU.r5_RNIB8HG5_12_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIB8HG5_12_LC_11_15_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r5_RNIB8HG5_12_LC_11_15_5  (
            .in0(N__54615),
            .in1(N__54025),
            .in2(N__53223),
            .in3(N__41351),
            .lcout(\ALU.r5_RNIB8HG5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_LC_11_15_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_LC_11_15_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_13_s1_c_RNO_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__55535),
            .in2(_gnd_net_),
            .in3(N__36140),
            .lcout(\ALU.r0_12_prm_8_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_10_s1_c_RNO_LC_11_16_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_10_s1_c_RNO_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_10_s1_c_RNO_LC_11_16_0 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_10_s1_c_RNO_LC_11_16_0  (
            .in0(N__55959),
            .in1(N__54049),
            .in2(_gnd_net_),
            .in3(N__36100),
            .lcout(\ALU.r0_12_prm_1_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_12_s0_c_RNO_LC_11_16_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_12_s0_c_RNO_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_12_s0_c_RNO_LC_11_16_1 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \ALU.r0_12_prm_1_12_s0_c_RNO_LC_11_16_1  (
            .in0(N__54050),
            .in1(N__55960),
            .in2(_gnd_net_),
            .in3(N__37586),
            .lcout(\ALU.r0_12_prm_1_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_0_s1_c_RNO_LC_12_1_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_0_s1_c_RNO_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_0_s1_c_RNO_LC_12_1_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_0_s1_c_RNO_LC_12_1_0  (
            .in0(N__53968),
            .in1(N__54806),
            .in2(N__53154),
            .in3(N__49015),
            .lcout(\ALU.r0_12_prm_4_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_0_s1_c_RNO_LC_12_1_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_0_s1_c_RNO_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_0_s1_c_RNO_LC_12_1_2 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_0_s1_c_RNO_LC_12_1_2  (
            .in0(N__54810),
            .in1(N__49014),
            .in2(N__53153),
            .in3(N__38030),
            .lcout(\ALU.r0_12_prm_5_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_6_s1_c_RNO_LC_12_1_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_6_s1_c_RNO_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_6_s1_c_RNO_LC_12_1_5 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_6_s1_c_RNO_LC_12_1_5  (
            .in0(N__55841),
            .in1(N__53969),
            .in2(_gnd_net_),
            .in3(N__38206),
            .lcout(\ALU.r0_12_prm_1_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJTDS9_0_5_LC_12_1_6 .C_ON=1'b0;
    defparam \ALU.r4_RNIJTDS9_0_5_LC_12_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJTDS9_0_5_LC_12_1_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r4_RNIJTDS9_0_5_LC_12_1_6  (
            .in0(N__53967),
            .in1(N__45494),
            .in2(N__54886),
            .in3(N__42848),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI9H7SJ_6_LC_12_1_7 .C_ON=1'b0;
    defparam \ALU.r4_RNI9H7SJ_6_LC_12_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI9H7SJ_6_LC_12_1_7 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNI9H7SJ_6_LC_12_1_7  (
            .in0(N__54805),
            .in1(N__43429),
            .in2(N__36349),
            .in3(N__44603),
            .lcout(\ALU.r4_RNI9H7SJZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_0_s1_c_LC_12_2_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_0_s1_c_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_0_s1_c_LC_12_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_0_s1_c_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__37504),
            .in2(N__40705),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\ALU.r0_12_prm_8_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_0_s1_c_LC_12_2_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_0_s1_c_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_0_s1_c_LC_12_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_0_s1_c_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(N__36346),
            .in2(N__36447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_0_s1 ),
            .carryout(\ALU.r0_12_prm_7_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_0_s1_c_LC_12_2_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_0_s1_c_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_0_s1_c_LC_12_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_0_s1_c_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__36334),
            .in2(N__36316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_0_s1 ),
            .carryout(\ALU.r0_12_prm_6_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_0_s1_c_LC_12_2_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_0_s1_c_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_0_s1_c_LC_12_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_0_s1_c_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(N__36292),
            .in2(N__37752),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_0_s1 ),
            .carryout(\ALU.r0_12_prm_5_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_0_s1_c_LC_12_2_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_0_s1_c_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_0_s1_c_LC_12_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_0_s1_c_LC_12_2_4  (
            .in0(_gnd_net_),
            .in1(N__36286),
            .in2(N__36280),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_0_s1 ),
            .carryout(\ALU.r0_12_prm_4_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_0_s1_c_LC_12_2_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_0_s1_c_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_0_s1_c_LC_12_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_0_s1_c_LC_12_2_5  (
            .in0(_gnd_net_),
            .in1(N__36463),
            .in2(N__36448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_0_s1 ),
            .carryout(\ALU.r0_12_prm_3_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_0_s1_c_LC_12_2_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_0_s1_c_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_0_s1_c_LC_12_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_0_s1_c_LC_12_2_6  (
            .in0(_gnd_net_),
            .in1(N__38116),
            .in2(N__40618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_0_s1 ),
            .carryout(\ALU.r0_12_prm_2_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_0_s1_c_LC_12_2_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_0_s1_c_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_0_s1_c_LC_12_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_0_s1_c_LC_12_2_7  (
            .in0(_gnd_net_),
            .in1(N__36415),
            .in2(N__36400),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_2_0_s1 ),
            .carryout(\ALU.r0_12_s1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_0_THRU_LUT4_0_LC_12_3_0 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_0_THRU_LUT4_0_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_0_THRU_LUT4_0_LC_12_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_0_THRU_LUT4_0_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36385),
            .lcout(\ALU.r0_12_s1_0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_5_s0_c_RNO_LC_12_3_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_5_s0_c_RNO_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_5_s0_c_RNO_LC_12_3_1 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_5_s0_c_RNO_LC_12_3_1  (
            .in0(N__45405),
            .in1(N__54651),
            .in2(N__53228),
            .in3(N__45260),
            .lcout(\ALU.r0_12_prm_5_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIO5SA91_2_LC_12_3_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIO5SA91_2_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIO5SA91_2_LC_12_3_2 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r4_RNIO5SA91_2_LC_12_3_2  (
            .in0(N__51080),
            .in1(N__48166),
            .in2(N__51491),
            .in3(N__41118),
            .lcout(\ALU.rshift_15_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_4_c_RNO_0_LC_12_3_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_4_c_RNO_0_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_4_c_RNO_0_LC_12_3_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r0_12_prm_5_4_c_RNO_0_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__42825),
            .in2(_gnd_net_),
            .in3(N__40534),
            .lcout(\ALU.r0_12_prm_5_4_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI97EK9_0_5_LC_12_3_6 .C_ON=1'b0;
    defparam \ALU.r4_RNI97EK9_0_5_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI97EK9_0_5_LC_12_3_6 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r4_RNI97EK9_0_5_LC_12_3_6  (
            .in0(N__53781),
            .in1(N__45404),
            .in2(N__54789),
            .in3(N__43420),
            .lcout(\ALU.rshift_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_0_s0_c_RNO_LC_12_3_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_0_s0_c_RNO_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_0_s0_c_RNO_LC_12_3_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_0_s0_c_RNO_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(N__40607),
            .in2(_gnd_net_),
            .in3(N__55736),
            .lcout(\ALU.r0_12_prm_2_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_1_c_RNO_LC_12_4_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_1_c_RNO_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_1_c_RNO_LC_12_4_0 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_1_c_RNO_LC_12_4_0  (
            .in0(N__53807),
            .in1(N__48617),
            .in2(N__53158),
            .in3(N__46749),
            .lcout(\ALU.r0_12_prm_6_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIK9PV9_15_LC_12_4_1 .C_ON=1'b0;
    defparam \ALU.r5_RNIK9PV9_15_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIK9PV9_15_LC_12_4_1 .LUT_INIT=16'b0001001100000011;
    LogicCell40 \ALU.r5_RNIK9PV9_15_LC_12_4_1  (
            .in0(N__54702),
            .in1(N__51003),
            .in2(N__51482),
            .in3(N__50621),
            .lcout(\ALU.rshift_15_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_3_c_RNO_0_LC_12_4_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_3_c_RNO_0_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_3_c_RNO_0_LC_12_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r0_12_prm_5_3_c_RNO_0_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__49341),
            .in2(_gnd_net_),
            .in3(N__44360),
            .lcout(\ALU.r0_12_prm_5_3_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIODO6K_7_LC_12_4_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIODO6K_7_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIODO6K_7_LC_12_4_3 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.r4_RNIODO6K_7_LC_12_4_3  (
            .in0(N__36826),
            .in1(N__46190),
            .in2(N__54813),
            .in3(N__44595),
            .lcout(\ALU.r4_RNIODO6KZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI9OH6A_1_LC_12_4_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI9OH6A_1_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI9OH6A_1_LC_12_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNI9OH6A_1_LC_12_4_4  (
            .in0(N__53806),
            .in1(N__48989),
            .in2(_gnd_net_),
            .in3(N__48616),
            .lcout(),
            .ltout(\ALU.r4_RNI9OH6AZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJH1SA_1_LC_12_4_5 .C_ON=1'b0;
    defparam \ALU.r4_RNIJH1SA_1_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJH1SA_1_LC_12_4_5 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \ALU.r4_RNIJH1SA_1_LC_12_4_5  (
            .in0(N__54701),
            .in1(N__51268),
            .in2(N__36820),
            .in3(N__51002),
            .lcout(\ALU.lshift_15_ns_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_6_s0_c_RNO_LC_12_4_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_6_s0_c_RNO_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_6_s0_c_RNO_LC_12_4_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_6_s0_c_RNO_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(N__55517),
            .in2(_gnd_net_),
            .in3(N__37688),
            .lcout(\ALU.r0_12_prm_8_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_a10_b_4_LC_12_5_0 .C_ON=1'b0;
    defparam \ALU.mult_a10_b_4_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_a10_b_4_LC_12_5_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \ALU.mult_a10_b_4_LC_12_5_0  (
            .in0(N__36817),
            .in1(N__36805),
            .in2(N__36768),
            .in3(N__40488),
            .lcout(\ALU.a10_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIHENK8_0_7_LC_12_5_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIHENK8_0_7_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIHENK8_0_7_LC_12_5_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNIHENK8_0_7_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__44805),
            .in2(_gnd_net_),
            .in3(N__44537),
            .lcout(\ALU.r4_RNIHENK8_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIFR136_7_LC_12_5_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIFR136_7_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIFR136_7_LC_12_5_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \ALU.r4_RNIFR136_7_LC_12_5_2  (
            .in0(N__44538),
            .in1(N__52719),
            .in2(N__54885),
            .in3(N__53874),
            .lcout(\ALU.r4_RNIFR136Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIF01FK_2_LC_12_5_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIF01FK_2_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIF01FK_2_LC_12_5_3 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.r4_RNIF01FK_2_LC_12_5_3  (
            .in0(N__49412),
            .in1(N__54796),
            .in2(N__36895),
            .in3(N__48400),
            .lcout(\ALU.r4_RNIF01FKZ0Z_2 ),
            .ltout(\ALU.r4_RNIF01FKZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIJCHBK1_6_LC_12_5_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIJCHBK1_6_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIJCHBK1_6_LC_12_5_4 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \ALU.r4_RNIJCHBK1_6_LC_12_5_4  (
            .in0(N__51414),
            .in1(N__36886),
            .in2(N__36877),
            .in3(N__36874),
            .lcout(\ALU.lshift_9 ),
            .ltout(\ALU.lshift_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_LC_12_5_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_LC_12_5_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \ALU.r0_12_prm_8_9_s1_c_RNO_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36856),
            .in3(N__55513),
            .lcout(\ALU.r0_12_prm_8_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_LC_12_5_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_LC_12_5_6 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \ALU.r0_12_prm_8_9_s0_c_RNO_LC_12_5_6  (
            .in0(N__42561),
            .in1(_gnd_net_),
            .in2(N__55534),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_8_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_4_c_RNO_LC_12_5_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_4_c_RNO_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_4_c_RNO_LC_12_5_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_7_4_c_RNO_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__52718),
            .in2(_gnd_net_),
            .in3(N__38463),
            .lcout(\ALU.r0_12_prm_7_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_7_s0_c_THRU_CRY_0_LC_12_6_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_7_s0_c_THRU_CRY_0_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_7_s0_c_THRU_CRY_0_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_7_s0_c_THRU_CRY_0_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__44169),
            .in2(N__44173),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\ALU.r0_12_prm_8_7_s0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_7_s0_c_LC_12_6_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_7_s0_c_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_7_s0_c_LC_12_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_7_s0_c_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__42985),
            .in2(N__44125),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_7_s0_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_7_s0_c_LC_12_6_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_7_s0_c_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_7_s0_c_LC_12_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_7_s0_c_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__48079),
            .in2(N__48004),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_7_s0 ),
            .carryout(\ALU.r0_12_prm_7_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_7_s0_c_LC_12_6_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_7_s0_c_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_7_s0_c_LC_12_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_7_s0_c_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__44095),
            .in2(N__36976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_7_s0 ),
            .carryout(\ALU.r0_12_prm_6_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_7_s0_c_LC_12_6_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_7_s0_c_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_7_s0_c_LC_12_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_7_s0_c_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__44055),
            .in2(N__43159),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_7_s0 ),
            .carryout(\ALU.r0_12_prm_5_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_7_s0_c_inv_LC_12_6_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_7_s0_c_inv_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_7_s0_c_inv_LC_12_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_7_s0_c_inv_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__44028),
            .in2(N__36964),
            .in3(N__44596),
            .lcout(\ALU.a_i_7 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_7_s0 ),
            .carryout(\ALU.r0_12_prm_4_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_7_s0_c_inv_LC_12_6_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_7_s0_c_inv_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_7_s0_c_inv_LC_12_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_7_s0_c_inv_LC_12_6_6  (
            .in0(N__55282),
            .in1(N__36955),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_7_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_7_s0 ),
            .carryout(\ALU.r0_12_prm_3_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_7_s0_c_LC_12_6_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_7_s0_c_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_7_s0_c_LC_12_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_7_s0_c_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__44013),
            .in2(N__38953),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_7_s0 ),
            .carryout(\ALU.r0_12_prm_2_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_7_s0_c_LC_12_7_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_7_s0_c_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_7_s0_c_LC_12_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_7_s0_c_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__45005),
            .in2(N__36949),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\ALU.r0_12_s0_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_7_s0_c_RNIJOSTUN1_LC_12_7_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_7_s0_c_RNIJOSTUN1_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_7_s0_c_RNIJOSTUN1_LC_12_7_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r0_12_prm_1_7_s0_c_RNIJOSTUN1_LC_12_7_1  (
            .in0(N__44914),
            .in1(N__36940),
            .in2(_gnd_net_),
            .in3(N__36925),
            .lcout(\ALU.r0_12_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_7_LC_12_7_2 .C_ON=1'b0;
    defparam \ALU.r1_7_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_7_LC_12_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_7_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38711),
            .lcout(r1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56241),
            .ce(N__47559),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_0_LC_12_8_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_0_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_0_LC_12_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_5_s0_c_RNO_0_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__38884),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\ALU.r0_12_prm_8_5_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s0_c_LC_12_8_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_5_s0_c_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s0_c_LC_12_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_5_s0_c_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__48151),
            .in2(N__48118),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_5_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_5_s0_c_LC_12_8_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_5_s0_c_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_5_s0_c_LC_12_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_5_s0_c_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__47267),
            .in2(N__37060),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_5_s0 ),
            .carryout(\ALU.r0_12_prm_7_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_5_s0_c_LC_12_8_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_5_s0_c_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_5_s0_c_LC_12_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_5_s0_c_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__44944),
            .in2(N__37042),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_5_s0 ),
            .carryout(\ALU.r0_12_prm_6_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_5_s0_c_LC_12_8_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_5_s0_c_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_5_s0_c_LC_12_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_5_s0_c_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__45766),
            .in2(N__37024),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_5_s0 ),
            .carryout(\ALU.r0_12_prm_5_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_5_s0_c_inv_LC_12_8_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_5_s0_c_inv_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_5_s0_c_inv_LC_12_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_5_s0_c_inv_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__45714),
            .in2(N__37012),
            .in3(N__45510),
            .lcout(\ALU.a_i_5 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_5_s0 ),
            .carryout(\ALU.r0_12_prm_4_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_5_s0_c_inv_LC_12_8_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_5_s0_c_inv_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_5_s0_c_inv_LC_12_8_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_5_s0_c_inv_LC_12_8_6  (
            .in0(N__55272),
            .in1(N__36994),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_5_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_5_s0 ),
            .carryout(\ALU.r0_12_prm_3_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_5_s0_c_LC_12_8_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_5_s0_c_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_5_s0_c_LC_12_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_5_s0_c_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__45687),
            .in2(N__36988),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_5_s0 ),
            .carryout(\ALU.r0_12_prm_2_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_5_s0_c_LC_12_9_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_5_s0_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_5_s0_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_5_s0_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__45625),
            .in2(N__44188),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\ALU.r0_12_s0_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_5_s0_c_RNITPI7KJ_LC_12_9_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_5_s0_c_RNITPI7KJ_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_5_s0_c_RNITPI7KJ_LC_12_9_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r0_12_prm_1_5_s0_c_RNITPI7KJ_LC_12_9_1  (
            .in0(N__45592),
            .in1(N__37234),
            .in2(_gnd_net_),
            .in3(N__37219),
            .lcout(\ALU.r0_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_5_LC_12_9_2 .C_ON=1'b0;
    defparam \ALU.r1_5_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_5_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_5_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37150),
            .lcout(r1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56249),
            .ce(N__47543),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_0_LC_12_10_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_0_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_0_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_8_s0_c_RNO_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__38614),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\ALU.r0_12_prm_8_8_s0_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s0_c_LC_12_10_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_8_s0_c_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s0_c_LC_12_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_8_s0_c_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__38917),
            .in2(N__39331),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_8_s0_cy ),
            .carryout(\ALU.r0_12_prm_8_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_8_s0_c_LC_12_10_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_8_s0_c_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_8_s0_c_LC_12_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_8_s0_c_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__38893),
            .in2(N__39292),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_8_s0 ),
            .carryout(\ALU.r0_12_prm_7_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_8_s0_c_LC_12_10_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_8_s0_c_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_8_s0_c_LC_12_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_8_s0_c_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__37084),
            .in2(N__39264),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_8_s0 ),
            .carryout(\ALU.r0_12_prm_6_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_8_s0_c_LC_12_10_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_8_s0_c_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_8_s0_c_LC_12_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_8_s0_c_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__40774),
            .in2(N__42025),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_8_s0 ),
            .carryout(\ALU.r0_12_prm_5_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_8_s0_c_inv_LC_12_10_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_8_s0_c_inv_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_8_s0_c_inv_LC_12_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_8_s0_c_inv_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__38980),
            .in2(N__39234),
            .in3(N__46180),
            .lcout(\ALU.a_i_8 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_8_s0 ),
            .carryout(\ALU.r0_12_prm_4_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_8_s0_c_inv_LC_12_10_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_8_s0_c_inv_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_8_s0_c_inv_LC_12_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.r0_12_prm_3_8_s0_c_inv_LC_12_10_6  (
            .in0(N__55268),
            .in1(N__37066),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_3_8_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_8_s0 ),
            .carryout(\ALU.r0_12_prm_3_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_8_s0_c_LC_12_10_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_8_s0_c_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_8_s0_c_LC_12_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_8_s0_c_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__39401),
            .in2(N__39370),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_8_s0 ),
            .carryout(\ALU.r0_12_prm_2_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_8_s0_c_LC_12_11_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_8_s0_c_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_8_s0_c_LC_12_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_8_s0_c_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__39618),
            .in2(N__37306),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\ALU.r0_12_s0_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s0_8_THRU_LUT4_0_LC_12_11_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s0_8_THRU_LUT4_0_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s0_8_THRU_LUT4_0_LC_12_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s0_8_THRU_LUT4_0_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37309),
            .lcout(\ALU.r0_12_s0_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_8_s1_c_RNO_LC_12_11_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_8_s1_c_RNO_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_8_s1_c_RNO_LC_12_11_3 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \ALU.r0_12_prm_1_8_s1_c_RNO_LC_12_11_3  (
            .in0(N__39617),
            .in1(N__55903),
            .in2(_gnd_net_),
            .in3(N__53897),
            .lcout(\ALU.r0_12_prm_1_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_8_s0_c_RNO_LC_12_11_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_8_s0_c_RNO_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_8_s0_c_RNO_LC_12_11_4 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_8_s0_c_RNO_LC_12_11_4  (
            .in0(N__55902),
            .in1(N__53896),
            .in2(_gnd_net_),
            .in3(N__39616),
            .lcout(\ALU.r0_12_prm_1_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_15_s1_c_RNO_LC_12_12_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_15_s1_c_RNO_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_15_s1_c_RNO_LC_12_12_0 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_15_s1_c_RNO_LC_12_12_0  (
            .in0(N__55940),
            .in1(N__54002),
            .in2(_gnd_net_),
            .in3(N__37283),
            .lcout(\ALU.r0_12_prm_1_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNISU5D9_0_9_LC_12_12_1 .C_ON=1'b0;
    defparam \ALU.r4_RNISU5D9_0_9_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNISU5D9_0_9_LC_12_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.r4_RNISU5D9_0_9_LC_12_12_1  (
            .in0(N__52322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47478),
            .lcout(\ALU.r4_RNISU5D9_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNISP2L9_1_12_LC_12_12_3 .C_ON=1'b0;
    defparam \ALU.r5_RNISP2L9_1_12_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNISP2L9_1_12_LC_12_12_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.r5_RNISP2L9_1_12_LC_12_12_3  (
            .in0(N__39877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41354),
            .lcout(\ALU.r5_RNISP2L9_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_12_s1_c_RNO_LC_12_12_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_12_s1_c_RNO_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_12_s1_c_RNO_LC_12_12_4 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \ALU.r0_12_prm_7_12_s1_c_RNO_LC_12_12_4  (
            .in0(N__41353),
            .in1(N__53064),
            .in2(_gnd_net_),
            .in3(N__39876),
            .lcout(\ALU.r0_12_prm_7_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_9_s1_c_RNO_LC_12_12_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_9_s1_c_RNO_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_9_s1_c_RNO_LC_12_12_6 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_9_s1_c_RNO_LC_12_12_6  (
            .in0(N__53175),
            .in1(N__47477),
            .in2(_gnd_net_),
            .in3(N__52321),
            .lcout(\ALU.r0_12_prm_7_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_LC_12_12_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_LC_12_12_7 .LUT_INIT=16'b1110000101001011;
    LogicCell40 \ALU.r0_12_prm_8_12_s1_c_RNO_LC_12_12_7  (
            .in0(N__51441),
            .in1(N__37485),
            .in2(N__55537),
            .in3(N__41024),
            .lcout(\ALU.r0_12_prm_8_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_0_LC_12_13_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_0_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_12_s1_c_RNO_0_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__38905),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\ALU.r0_12_prm_8_12_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s1_c_LC_12_13_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_12_s1_c_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s1_c_LC_12_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_12_s1_c_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__37474),
            .in2(N__37464),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_12_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_12_s1_c_LC_12_13_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_12_s1_c_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_12_s1_c_LC_12_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_12_s1_c_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__37447),
            .in2(N__37441),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_12_s1 ),
            .carryout(\ALU.r0_12_prm_7_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_12_s1_c_LC_12_13_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_12_s1_c_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_12_s1_c_LC_12_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_12_s1_c_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__37414),
            .in2(N__39718),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_12_s1 ),
            .carryout(\ALU.r0_12_prm_6_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_12_s1_c_LC_12_13_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_12_s1_c_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_12_s1_c_LC_12_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_12_s1_c_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__37384),
            .in2(N__37362),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_12_s1 ),
            .carryout(\ALU.r0_12_prm_5_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_12_s1_c_LC_12_13_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_12_s1_c_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_12_s1_c_LC_12_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_12_s1_c_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__37345),
            .in2(N__37333),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_12_s1 ),
            .carryout(\ALU.r0_12_prm_4_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_12_s1_c_LC_12_13_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_12_s1_c_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_12_s1_c_LC_12_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_12_s1_c_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__55280),
            .in2(N__56508),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_12_s1 ),
            .carryout(\ALU.r0_12_prm_3_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_12_s1_c_LC_12_13_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_12_s1_c_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_12_s1_c_LC_12_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_12_s1_c_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__37650),
            .in2(N__37615),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_12_s1 ),
            .carryout(\ALU.r0_12_prm_2_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_12_s1_c_LC_12_14_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_12_s1_c_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_12_s1_c_LC_12_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_12_s1_c_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__37603),
            .in2(N__37593),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\ALU.r0_12_s1_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_12_THRU_LUT4_0_LC_12_14_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_12_THRU_LUT4_0_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_12_THRU_LUT4_0_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_12_THRU_LUT4_0_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37555),
            .lcout(\ALU.r0_12_s1_12_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_15_s1_c_RNO_LC_12_15_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_15_s1_c_RNO_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_15_s1_c_RNO_LC_12_15_2 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_15_s1_c_RNO_LC_12_15_2  (
            .in0(N__54782),
            .in1(N__40158),
            .in2(N__52963),
            .in3(N__40007),
            .lcout(\ALU.r0_12_prm_5_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_1_LC_13_1_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_1_LC_13_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_15_s1_c_RNO_1_LC_13_1_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.r0_12_prm_8_15_s1_c_RNO_1_LC_13_1_1  (
            .in0(N__54802),
            .in1(N__53964),
            .in2(N__50679),
            .in3(N__40183),
            .lcout(\ALU.r0_12_prm_8_15_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam params_3_LC_13_1_3.C_ON=1'b0;
    defparam params_3_LC_13_1_3.SEQ_MODE=4'b1000;
    defparam params_3_LC_13_1_3.LUT_INIT=16'b0110110011001100;
    LogicCell40 params_3_LC_13_1_3 (
            .in0(N__54803),
            .in1(N__51224),
            .in2(N__50932),
            .in3(N__53966),
            .lcout(paramsZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56227),
            .ce(N__56057),
            .sr(_gnd_net_));
    defparam params_2_LC_13_1_4.C_ON=1'b0;
    defparam params_2_LC_13_1_4.SEQ_MODE=4'b1000;
    defparam params_2_LC_13_1_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 params_2_LC_13_1_4 (
            .in0(N__53965),
            .in1(N__50856),
            .in2(_gnd_net_),
            .in3(N__54804),
            .lcout(paramsZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56227),
            .ce(N__56057),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_0_s1_c_RNO_LC_13_1_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_0_s1_c_RNO_LC_13_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_0_s1_c_RNO_LC_13_1_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_0_s1_c_RNO_LC_13_1_6  (
            .in0(_gnd_net_),
            .in1(N__55489),
            .in2(_gnd_net_),
            .in3(N__40694),
            .lcout(\ALU.r0_12_prm_8_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIAV175_15_LC_13_1_7 .C_ON=1'b0;
    defparam \ALU.r5_RNIAV175_15_LC_13_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIAV175_15_LC_13_1_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ALU.r5_RNIAV175_15_LC_13_1_7  (
            .in0(N__54801),
            .in1(N__53963),
            .in2(N__50931),
            .in3(N__40182),
            .lcout(\ALU.r5_RNIAV175Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.lshift63_2_LC_13_2_0 .C_ON=1'b0;
    defparam \ALU.lshift63_2_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.lshift63_2_LC_13_2_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ALU.lshift63_2_LC_13_2_0  (
            .in0(_gnd_net_),
            .in1(N__51212),
            .in2(_gnd_net_),
            .in3(N__50873),
            .lcout(\ALU.lshift63Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_0_s1_c_RNO_LC_13_2_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_0_s1_c_RNO_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_0_s1_c_RNO_LC_13_2_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_0_s1_c_RNO_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(N__55722),
            .in2(_gnd_net_),
            .in3(N__40606),
            .lcout(\ALU.r0_12_prm_2_0_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIHENK8_7_LC_13_2_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIHENK8_7_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIHENK8_7_LC_13_2_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r4_RNIHENK8_7_LC_13_2_3  (
            .in0(_gnd_net_),
            .in1(N__44784),
            .in2(_gnd_net_),
            .in3(N__44600),
            .lcout(\ALU.un14_log_0_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_RNO_2_LC_13_2_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_2_c_RNO_2_LC_13_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_RNO_2_LC_13_2_4 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r0_12_prm_8_2_c_RNO_2_LC_13_2_4  (
            .in0(N__50874),
            .in1(N__38110),
            .in2(N__51296),
            .in3(N__38098),
            .lcout(),
            .ltout(\ALU.rshift_15_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_RNO_1_LC_13_2_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_2_c_RNO_1_LC_13_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_RNO_1_LC_13_2_5 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.r0_12_prm_8_2_c_RNO_1_LC_13_2_5  (
            .in0(N__38083),
            .in1(N__51221),
            .in2(N__38062),
            .in3(N__38059),
            .lcout(\ALU.rshift_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_6_s0_c_RNO_LC_13_2_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_6_s0_c_RNO_LC_13_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_6_s0_c_RNO_LC_13_2_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_6_s0_c_RNO_LC_13_2_6  (
            .in0(_gnd_net_),
            .in1(N__55723),
            .in2(_gnd_net_),
            .in3(N__38265),
            .lcout(\ALU.r0_12_prm_2_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNID26E8_0_0_LC_13_2_7 .C_ON=1'b0;
    defparam \ALU.r4_RNID26E8_0_0_LC_13_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNID26E8_0_0_LC_13_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r4_RNID26E8_0_0_LC_13_2_7  (
            .in0(_gnd_net_),
            .in1(N__49000),
            .in2(_gnd_net_),
            .in3(N__38032),
            .lcout(\ALU.r4_RNID26E8_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_6_s0_c_THRU_CRY_0_LC_13_3_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_6_s0_c_THRU_CRY_0_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_6_s0_c_THRU_CRY_0_LC_13_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_6_s0_c_THRU_CRY_0_LC_13_3_0  (
            .in0(_gnd_net_),
            .in1(N__37730),
            .in2(N__37735),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_3_0_),
            .carryout(\ALU.r0_12_prm_8_6_s0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_6_s0_c_LC_13_3_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_6_s0_c_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_6_s0_c_LC_13_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_6_s0_c_LC_13_3_1  (
            .in0(_gnd_net_),
            .in1(N__37693),
            .in2(N__37663),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_6_s0_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_6_s0_c_LC_13_3_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_6_s0_c_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_6_s0_c_LC_13_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_6_s0_c_LC_13_3_2  (
            .in0(_gnd_net_),
            .in1(N__41649),
            .in2(N__41602),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_6_s0 ),
            .carryout(\ALU.r0_12_prm_7_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_6_s0_c_LC_13_3_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_6_s0_c_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_6_s0_c_LC_13_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_6_s0_c_LC_13_3_3  (
            .in0(_gnd_net_),
            .in1(N__38365),
            .in2(N__41587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_6_s0 ),
            .carryout(\ALU.r0_12_prm_6_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_6_s0_c_LC_13_3_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_6_s0_c_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_6_s0_c_LC_13_3_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_6_s0_c_LC_13_3_4  (
            .in0(_gnd_net_),
            .in1(N__38341),
            .in2(N__43174),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_6_s0 ),
            .carryout(\ALU.r0_12_prm_5_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_6_s0_c_inv_LC_13_3_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_6_s0_c_inv_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_6_s0_c_inv_LC_13_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_6_s0_c_inv_LC_13_3_5  (
            .in0(_gnd_net_),
            .in1(N__38289),
            .in2(N__38317),
            .in3(N__43436),
            .lcout(\ALU.a_i_6 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_6_s0 ),
            .carryout(\ALU.r0_12_prm_4_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_6_s0_c_inv_LC_13_3_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_6_s0_c_inv_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_6_s0_c_inv_LC_13_3_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_3_6_s0_c_inv_LC_13_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38275),
            .in3(N__55172),
            .lcout(\ALU.r0_12_prm_3_6_s0_sf ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_6_s0 ),
            .carryout(\ALU.r0_12_prm_3_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_6_s0_c_LC_13_3_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_6_s0_c_LC_13_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_6_s0_c_LC_13_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_6_s0_c_LC_13_3_7  (
            .in0(_gnd_net_),
            .in1(N__38258),
            .in2(N__38215),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_6_s0 ),
            .carryout(\ALU.r0_12_prm_2_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_6_s0_c_LC_13_4_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_6_s0_c_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_6_s0_c_LC_13_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_6_s0_c_LC_13_4_0  (
            .in0(_gnd_net_),
            .in1(N__38205),
            .in2(N__38161),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_4_0_),
            .carryout(\ALU.r0_12_s0_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_6_s0_c_RNINEODV21_LC_13_4_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_6_s0_c_RNINEODV21_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_6_s0_c_RNINEODV21_LC_13_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r0_12_prm_1_6_s0_c_RNINEODV21_LC_13_4_1  (
            .in0(N__38146),
            .in1(N__38134),
            .in2(_gnd_net_),
            .in3(N__38119),
            .lcout(\ALU.r0_12_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r1_6_LC_13_4_2 .C_ON=1'b0;
    defparam \ALU.r1_6_LC_13_4_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r1_6_LC_13_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r1_6_LC_13_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38815),
            .lcout(r1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56230),
            .ce(N__47577),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_THRU_CRY_0_LC_13_5_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_4_c_THRU_CRY_0_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_THRU_CRY_0_LC_13_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_4_c_THRU_CRY_0_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__41067),
            .in2(N__41071),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_5_0_),
            .carryout(\ALU.r0_12_prm_8_4_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_LC_13_5_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_4_c_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_LC_13_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_4_c_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(N__41803),
            .in2(N__40756),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_4_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_4_c_LC_13_5_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_4_c_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_4_c_LC_13_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_4_c_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(N__38467),
            .in2(N__38434),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_4 ),
            .carryout(\ALU.r0_12_prm_7_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_4_c_LC_13_5_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_4_c_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_4_c_LC_13_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_4_c_LC_13_5_3  (
            .in0(_gnd_net_),
            .in1(N__38425),
            .in2(N__38410),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_4 ),
            .carryout(\ALU.r0_12_prm_6_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_4_c_LC_13_5_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_4_c_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_4_c_LC_13_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_4_c_LC_13_5_4  (
            .in0(_gnd_net_),
            .in1(N__40342),
            .in2(N__38395),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_4 ),
            .carryout(\ALU.r0_12_prm_5_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_4_c_inv_LC_13_5_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_4_c_inv_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_4_c_inv_LC_13_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_4_c_inv_LC_13_5_5  (
            .in0(_gnd_net_),
            .in1(N__38383),
            .in2(N__42616),
            .in3(N__42851),
            .lcout(\ALU.a_i_4 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_4 ),
            .carryout(\ALU.r0_12_prm_4_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_4_c_LC_13_5_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_4_c_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_4_c_LC_13_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_4_c_LC_13_5_6  (
            .in0(_gnd_net_),
            .in1(N__38530),
            .in2(N__38377),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_4 ),
            .carryout(\ALU.r0_12_prm_3_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_4_c_LC_13_5_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_4_c_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_4_c_LC_13_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_4_c_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__38602),
            .in2(N__38578),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_4 ),
            .carryout(\ALU.r0_12_prm_2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_4_c_LC_13_6_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_4_c_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_4_c_LC_13_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_4_c_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__41761),
            .in2(N__41737),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\ALU.r0_12_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_4_THRU_LUT4_0_LC_13_6_1 .C_ON=1'b0;
    defparam \ALU.r0_12_4_THRU_LUT4_0_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_4_THRU_LUT4_0_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_4_THRU_LUT4_0_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38659),
            .lcout(\ALU.r0_12_4_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI0QK3K_11_LC_13_6_2 .C_ON=1'b0;
    defparam \ALU.r5_RNI0QK3K_11_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI0QK3K_11_LC_13_6_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.r5_RNI0QK3K_11_LC_13_6_2  (
            .in0(N__38656),
            .in1(N__54795),
            .in2(_gnd_net_),
            .in3(N__38632),
            .lcout(\ALU.r5_RNI0QK3KZ0Z_11 ),
            .ltout(\ALU.r5_RNI0QK3KZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_1_LC_13_6_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_1_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_1_LC_13_6_3 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ALU.r0_12_prm_8_8_s0_c_RNO_1_LC_13_6_3  (
            .in0(N__50984),
            .in1(N__51359),
            .in2(N__38617),
            .in3(N__41686),
            .lcout(\ALU.rshift_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_1_LC_13_6_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_1_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_1_LC_13_6_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ALU.r0_12_prm_8_8_s1_c_RNO_1_LC_13_6_4  (
            .in0(N__41687),
            .in1(N__50985),
            .in2(N__51446),
            .in3(N__41091),
            .lcout(\ALU.r0_12_prm_8_8_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_4_c_RNO_LC_13_6_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_4_c_RNO_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_4_c_RNO_LC_13_6_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_4_c_RNO_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__55729),
            .in2(_gnd_net_),
            .in3(N__38598),
            .lcout(\ALU.r0_12_prm_2_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_4_c_RNO_LC_13_6_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_3_4_c_RNO_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_4_c_RNO_LC_13_6_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.r0_12_prm_3_4_c_RNO_LC_13_6_6  (
            .in0(N__55261),
            .in1(N__38569),
            .in2(_gnd_net_),
            .in3(N__38548),
            .lcout(\ALU.r0_12_prm_3_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIR63FA_4_LC_13_6_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIR63FA_4_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIR63FA_4_LC_13_6_7 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r4_RNIR63FA_4_LC_13_6_7  (
            .in0(N__53805),
            .in1(N__42850),
            .in2(N__54884),
            .in3(N__49408),
            .lcout(\ALU.lshift_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_LC_13_7_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_LC_13_7_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_8_8_s1_c_RNO_LC_13_7_1  (
            .in0(N__55400),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39317),
            .lcout(\ALU.r0_12_prm_8_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_7_s0_c_RNO_LC_13_7_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_7_s0_c_RNO_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_7_s0_c_RNO_LC_13_7_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_7_s0_c_RNO_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__55730),
            .in2(_gnd_net_),
            .in3(N__44014),
            .lcout(\ALU.r0_12_prm_2_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNILGU5F1_5_LC_13_7_3 .C_ON=1'b0;
    defparam \ALU.r4_RNILGU5F1_5_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNILGU5F1_5_LC_13_7_3 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \ALU.r4_RNILGU5F1_5_LC_13_7_3  (
            .in0(N__41056),
            .in1(N__38944),
            .in2(N__51301),
            .in3(N__41043),
            .lcout(\ALU.lshift_8 ),
            .ltout(\ALU.lshift_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_LC_13_7_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s0_c_RNO_LC_13_7_4 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \ALU.r0_12_prm_8_8_s0_c_RNO_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38920),
            .in3(N__55399),
            .lcout(\ALU.r0_12_prm_8_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_1_LC_13_7_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_1_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_12_s1_c_RNO_1_LC_13_7_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.r0_12_prm_8_12_s1_c_RNO_1_LC_13_7_5  (
            .in0(N__51231),
            .in1(N__51032),
            .in2(_gnd_net_),
            .in3(N__41685),
            .lcout(\ALU.r0_12_prm_8_12_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_8_s0_c_RNO_LC_13_7_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_8_s0_c_RNO_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_8_s0_c_RNO_LC_13_7_6 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_8_s0_c_RNO_LC_13_7_6  (
            .in0(N__52544),
            .in1(N__46382),
            .in2(_gnd_net_),
            .in3(N__46220),
            .lcout(\ALU.r0_12_prm_7_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_1_LC_13_7_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_1_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_1_LC_13_7_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ALU.r0_12_prm_8_5_s0_c_RNO_1_LC_13_7_7  (
            .in0(N__51102),
            .in1(N__43144),
            .in2(N__51302),
            .in3(N__41662),
            .lcout(\ALU.rshift_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r6_6_LC_13_8_0 .C_ON=1'b0;
    defparam \ALU.r6_6_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_6_LC_13_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_6_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38827),
            .lcout(r6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(N__45846),
            .sr(_gnd_net_));
    defparam \ALU.r6_7_LC_13_8_1 .C_ON=1'b0;
    defparam \ALU.r6_7_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_7_LC_13_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_7_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38712),
            .lcout(r6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(N__45846),
            .sr(_gnd_net_));
    defparam \ALU.r6_8_LC_13_8_2 .C_ON=1'b0;
    defparam \ALU.r6_8_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_8_LC_13_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_8_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39494),
            .lcout(r6_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(N__45846),
            .sr(_gnd_net_));
    defparam \ALU.r6_2_LC_13_8_3 .C_ON=1'b0;
    defparam \ALU.r6_2_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_2_LC_13_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_2_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40243),
            .lcout(r6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(N__45846),
            .sr(_gnd_net_));
    defparam \ALU.r6_3_LC_13_8_4 .C_ON=1'b0;
    defparam \ALU.r6_3_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_3_LC_13_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_3_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50159),
            .lcout(r6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(N__45846),
            .sr(_gnd_net_));
    defparam \ALU.r6_4_LC_13_8_5 .C_ON=1'b0;
    defparam \ALU.r6_4_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \ALU.r6_4_LC_13_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r6_4_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39043),
            .lcout(r6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(N__45846),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_RNO_LC_13_9_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_3_c_RNO_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_RNO_LC_13_9_1 .LUT_INIT=16'b0001111000001111;
    LogicCell40 \ALU.r0_12_prm_8_3_c_RNO_LC_13_9_1  (
            .in0(N__51039),
            .in1(N__51244),
            .in2(N__55522),
            .in3(N__50765),
            .lcout(\ALU.r0_12_prm_8_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIN3236_8_LC_13_9_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIN3236_8_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIN3236_8_LC_13_9_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \ALU.r4_RNIN3236_8_LC_13_9_2  (
            .in0(N__52819),
            .in1(N__54057),
            .in2(N__46227),
            .in3(N__54914),
            .lcout(\ALU.r4_RNIN3236Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_8_s1_c_RNO_LC_13_9_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_8_s1_c_RNO_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_8_s1_c_RNO_LC_13_9_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \ALU.r0_12_prm_4_8_s1_c_RNO_LC_13_9_4  (
            .in0(N__52820),
            .in1(N__54058),
            .in2(N__46228),
            .in3(N__54915),
            .lcout(\ALU.r0_12_prm_4_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_RNO_3_LC_13_9_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_1_c_RNO_3_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_RNO_3_LC_13_9_5 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.r0_12_prm_8_1_c_RNO_3_LC_13_9_5  (
            .in0(N__38974),
            .in1(N__42861),
            .in2(N__54924),
            .in3(N__49425),
            .lcout(),
            .ltout(\ALU.r0_12_prm_8_1_c_RNOZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_RNO_2_LC_13_9_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_1_c_RNO_2_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_RNO_2_LC_13_9_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.r0_12_prm_8_1_c_RNO_2_LC_13_9_6  (
            .in0(N__51245),
            .in1(N__51040),
            .in2(N__38956),
            .in3(N__41796),
            .lcout(),
            .ltout(\ALU.rshift_15_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_RNO_1_LC_13_9_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_1_c_RNO_1_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_RNO_1_LC_13_9_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r0_12_prm_8_1_c_RNO_1_LC_13_9_7  (
            .in0(N__51246),
            .in1(N__43140),
            .in2(N__39346),
            .in3(N__43065),
            .lcout(\ALU.rshift_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_0_LC_13_10_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_0_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s1_c_RNO_0_LC_13_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_8_s1_c_RNO_0_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\ALU.r0_12_prm_8_8_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_8_s1_c_LC_13_10_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_8_s1_c_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_8_s1_c_LC_13_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_8_s1_c_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__39327),
            .in2(N__39304),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_8_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_8_s1_c_LC_13_10_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_8_s1_c_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_8_s1_c_LC_13_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_8_s1_c_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__39291),
            .in2(N__45922),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_8_s1 ),
            .carryout(\ALU.r0_12_prm_7_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_8_s1_c_LC_13_10_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_8_s1_c_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_8_s1_c_LC_13_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_8_s1_c_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__39265),
            .in2(N__42007),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_8_s1 ),
            .carryout(\ALU.r0_12_prm_6_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_8_s1_c_LC_13_10_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_8_s1_c_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_8_s1_c_LC_13_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_8_s1_c_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__42021),
            .in2(N__45580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_8_s1 ),
            .carryout(\ALU.r0_12_prm_5_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_8_s1_c_LC_13_10_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_8_s1_c_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_8_s1_c_LC_13_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_8_s1_c_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__39241),
            .in2(N__39235),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_8_s1 ),
            .carryout(\ALU.r0_12_prm_4_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_8_s1_c_LC_13_10_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_8_s1_c_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_8_s1_c_LC_13_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_8_s1_c_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__55192),
            .in2(N__56475),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_8_s1 ),
            .carryout(\ALU.r0_12_prm_3_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_8_s1_c_LC_13_10_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_8_s1_c_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_8_s1_c_LC_13_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_8_s1_c_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__39402),
            .in2(N__39217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_8_s1 ),
            .carryout(\ALU.r0_12_prm_2_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_8_s1_c_LC_13_11_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_8_s1_c_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_8_s1_c_LC_13_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_8_s1_c_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__39622),
            .in2(N__39589),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\ALU.r0_12_s1_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_8_s0_c_RNIO9TN7H2_LC_13_11_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_8_s0_c_RNIO9TN7H2_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_8_s0_c_RNIO9TN7H2_LC_13_11_1 .LUT_INIT=16'b1111011010010000;
    LogicCell40 \ALU.r0_12_prm_1_8_s0_c_RNIO9TN7H2_LC_13_11_1  (
            .in0(N__39580),
            .in1(N__39562),
            .in2(N__39538),
            .in3(N__39529),
            .lcout(\ALU.r0_12_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_8_LC_13_11_2 .C_ON=1'b0;
    defparam \ALU.r0_8_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.r0_8_LC_13_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_8_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39472),
            .lcout(r0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56252),
            .ce(N__49716),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_9_s1_c_RNO_LC_13_12_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_9_s1_c_RNO_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_9_s1_c_RNO_LC_13_12_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_2_9_s1_c_RNO_LC_13_12_0  (
            .in0(N__55900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42440),
            .lcout(\ALU.r0_12_prm_2_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_8_s0_c_RNO_LC_13_12_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_8_s0_c_RNO_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_8_s0_c_RNO_LC_13_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_8_s0_c_RNO_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__55899),
            .in2(_gnd_net_),
            .in3(N__39403),
            .lcout(\ALU.r0_12_prm_2_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNITTMB9_12_LC_13_12_3 .C_ON=1'b0;
    defparam \ALU.r5_RNITTMB9_12_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNITTMB9_12_LC_13_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r5_RNITTMB9_12_LC_13_12_3  (
            .in0(N__53996),
            .in1(N__41352),
            .in2(_gnd_net_),
            .in3(N__40962),
            .lcout(\ALU.r5_RNITTMB9Z0Z_12 ),
            .ltout(\ALU.r5_RNITTMB9Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI355TI_13_LC_13_12_4 .C_ON=1'b0;
    defparam \ALU.r5_RNI355TI_13_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI355TI_13_LC_13_12_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.r5_RNI355TI_13_LC_13_12_4  (
            .in0(N__54858),
            .in1(_gnd_net_),
            .in2(N__39349),
            .in3(N__39709),
            .lcout(\ALU.r5_RNI355TIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_9_s1_c_RNO_LC_13_12_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_9_s1_c_RNO_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_9_s1_c_RNO_LC_13_12_5 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_9_s1_c_RNO_LC_13_12_5  (
            .in0(N__54584),
            .in1(N__47482),
            .in2(N__53205),
            .in3(N__52221),
            .lcout(\ALU.r0_12_prm_5_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_9_s1_c_RNO_LC_13_12_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_9_s1_c_RNO_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_9_s1_c_RNO_LC_13_12_6 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_9_s1_c_RNO_LC_13_12_6  (
            .in0(N__55901),
            .in1(N__53997),
            .in2(_gnd_net_),
            .in3(N__42395),
            .lcout(\ALU.r0_12_prm_1_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_1_LC_13_12_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_1_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_1_LC_13_12_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r0_12_prm_8_9_s1_c_RNO_1_LC_13_12_7  (
            .in0(N__51037),
            .in1(N__43139),
            .in2(N__51304),
            .in3(N__43066),
            .lcout(\ALU.r0_12_prm_8_9_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_14_s1_c_RNO_LC_13_13_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_14_s1_c_RNO_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_14_s1_c_RNO_LC_13_13_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_14_s1_c_RNO_LC_13_13_0  (
            .in0(N__54906),
            .in1(N__53960),
            .in2(N__53206),
            .in3(N__47008),
            .lcout(\ALU.r0_12_prm_4_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNITG1F5_14_LC_13_13_1 .C_ON=1'b0;
    defparam \ALU.r5_RNITG1F5_14_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNITG1F5_14_LC_13_13_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r5_RNITG1F5_14_LC_13_13_1  (
            .in0(N__53961),
            .in1(N__54907),
            .in2(N__53239),
            .in3(N__47031),
            .lcout(\ALU.r5_RNITG1F5Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_14_s0_c_RNO_LC_13_13_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_14_s0_c_RNO_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_14_s0_c_RNO_LC_13_13_2 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_14_s0_c_RNO_LC_13_13_2  (
            .in0(N__47185),
            .in1(N__53180),
            .in2(N__54923),
            .in3(N__47010),
            .lcout(\ALU.r0_12_prm_5_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_1_LC_13_13_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_1_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s0_c_RNO_1_LC_13_13_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.r0_12_prm_8_13_s0_c_RNO_1_LC_13_13_3  (
            .in0(N__51300),
            .in1(N__51038),
            .in2(_gnd_net_),
            .in3(N__43128),
            .lcout(\ALU.rshift_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_14_s0_c_RNO_LC_13_13_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_14_s0_c_RNO_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_14_s0_c_RNO_LC_13_13_4 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_14_s0_c_RNO_LC_13_13_4  (
            .in0(N__47184),
            .in1(N__53962),
            .in2(N__53207),
            .in3(N__47009),
            .lcout(\ALU.r0_12_prm_6_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_LC_13_13_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_LC_13_13_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_8_14_s0_c_RNO_LC_13_13_5  (
            .in0(N__47969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55533),
            .lcout(\ALU.r0_12_prm_8_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_14_s1_c_RNO_LC_13_13_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_14_s1_c_RNO_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_14_s1_c_RNO_LC_13_13_7 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_14_s1_c_RNO_LC_13_13_7  (
            .in0(N__53176),
            .in1(N__47183),
            .in2(_gnd_net_),
            .in3(N__47030),
            .lcout(\ALU.r0_12_prm_7_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIUH636_3_LC_13_14_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIUH636_3_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIUH636_3_LC_13_14_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r4_RNIUH636_3_LC_13_14_1  (
            .in0(N__54905),
            .in1(N__53958),
            .in2(N__53182),
            .in3(N__49426),
            .lcout(\ALU.r4_RNIUH636Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_15_s0_c_RNO_LC_13_14_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_15_s0_c_RNO_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_15_s0_c_RNO_LC_13_14_4 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_15_s0_c_RNO_LC_13_14_4  (
            .in0(N__53014),
            .in1(N__40157),
            .in2(_gnd_net_),
            .in3(N__40008),
            .lcout(\ALU.r0_12_prm_7_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_14_s1_c_RNO_LC_13_14_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_14_s1_c_RNO_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_14_s1_c_RNO_LC_13_14_5 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_14_s1_c_RNO_LC_13_14_5  (
            .in0(N__53957),
            .in1(N__47197),
            .in2(N__53181),
            .in3(N__47052),
            .lcout(\ALU.r0_12_prm_6_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_1_LC_13_14_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_1_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_13_s1_c_RNO_1_LC_13_14_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ALU.r0_12_prm_8_13_s1_c_RNO_1_LC_13_14_6  (
            .in0(N__43127),
            .in1(N__51303),
            .in2(_gnd_net_),
            .in3(N__51099),
            .lcout(\ALU.r0_12_prm_8_13_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_12_s1_c_RNO_LC_13_14_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_12_s1_c_RNO_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_12_s1_c_RNO_LC_13_14_7 .LUT_INIT=16'b1100000010010101;
    LogicCell40 \ALU.r0_12_prm_6_12_s1_c_RNO_LC_13_14_7  (
            .in0(N__39872),
            .in1(N__53959),
            .in2(N__53183),
            .in3(N__41355),
            .lcout(\ALU.r0_12_prm_6_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIPV8A9_0_13_LC_13_15_5 .C_ON=1'b0;
    defparam \ALU.r5_RNIPV8A9_0_13_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIPV8A9_0_13_LC_13_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r5_RNIPV8A9_0_13_LC_13_15_5  (
            .in0(N__53956),
            .in1(N__41478),
            .in2(_gnd_net_),
            .in3(N__47050),
            .lcout(\ALU.r5_RNIPV8A9_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_THRU_CRY_0_LC_14_1_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_2_c_THRU_CRY_0_LC_14_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_THRU_CRY_0_LC_14_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_2_c_THRU_CRY_0_LC_14_1_0  (
            .in0(_gnd_net_),
            .in1(N__39696),
            .in2(N__39700),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_1_0_),
            .carryout(\ALU.r0_12_prm_8_2_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_LC_14_1_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_2_c_LC_14_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_LC_14_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_2_c_LC_14_1_1  (
            .in0(_gnd_net_),
            .in1(N__40204),
            .in2(N__40213),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_2_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_2_c_LC_14_1_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_2_c_LC_14_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_2_c_LC_14_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_2_c_LC_14_1_2  (
            .in0(_gnd_net_),
            .in1(N__40746),
            .in2(N__40714),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_2 ),
            .carryout(\ALU.r0_12_prm_7_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_2_c_LC_14_1_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_2_c_LC_14_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_2_c_LC_14_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_2_c_LC_14_1_3  (
            .in0(_gnd_net_),
            .in1(N__40543),
            .in2(N__42937),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_2 ),
            .carryout(\ALU.r0_12_prm_6_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_2_c_LC_14_1_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_2_c_LC_14_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_2_c_LC_14_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_2_c_LC_14_1_4  (
            .in0(_gnd_net_),
            .in1(N__40336),
            .in2(N__43723),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_2 ),
            .carryout(\ALU.r0_12_prm_5_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_2_c_inv_LC_14_1_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_2_c_inv_LC_14_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_2_c_inv_LC_14_1_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_2_c_inv_LC_14_1_5  (
            .in0(_gnd_net_),
            .in1(N__40324),
            .in2(N__40312),
            .in3(N__48405),
            .lcout(\ALU.a_i_2 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_2 ),
            .carryout(\ALU.r0_12_prm_4_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_2_c_LC_14_1_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_2_c_LC_14_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_2_c_LC_14_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_2_c_LC_14_1_6  (
            .in0(_gnd_net_),
            .in1(N__42874),
            .in2(N__42925),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_2 ),
            .carryout(\ALU.r0_12_prm_3_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_2_c_LC_14_1_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_2_c_LC_14_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_2_c_LC_14_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_2_c_LC_14_1_7  (
            .in0(_gnd_net_),
            .in1(N__40552),
            .in2(N__40579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_2 ),
            .carryout(\ALU.r0_12_prm_2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_2_c_LC_14_2_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_2_c_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_2_c_LC_14_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_2_c_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(N__43708),
            .in2(N__43678),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_2_0_),
            .carryout(\ALU.r0_12_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_2_THRU_LUT4_0_LC_14_2_1 .C_ON=1'b0;
    defparam \ALU.r0_12_2_THRU_LUT4_0_LC_14_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_2_THRU_LUT4_0_LC_14_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_2_THRU_LUT4_0_LC_14_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40303),
            .lcout(\ALU.r0_12_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_RNO_0_LC_14_2_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_2_c_RNO_0_LC_14_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_RNO_0_LC_14_2_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.r0_12_prm_8_2_c_RNO_0_LC_14_2_2  (
            .in0(N__51223),
            .in1(N__50878),
            .in2(_gnd_net_),
            .in3(N__42204),
            .lcout(\ALU.lshift_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_2_c_RNO_LC_14_2_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_2_c_RNO_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_2_c_RNO_LC_14_2_4 .LUT_INIT=16'b0011011000110011;
    LogicCell40 \ALU.r0_12_prm_8_2_c_RNO_LC_14_2_4  (
            .in0(N__51222),
            .in1(N__55491),
            .in2(N__50961),
            .in3(N__42203),
            .lcout(\ALU.r0_12_prm_8_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_0_s0_c_RNO_LC_14_2_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_0_s0_c_RNO_LC_14_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_0_s0_c_RNO_LC_14_2_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_0_s0_c_RNO_LC_14_2_6  (
            .in0(_gnd_net_),
            .in1(N__55490),
            .in2(_gnd_net_),
            .in3(N__40687),
            .lcout(\ALU.r0_12_prm_8_0_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_2_c_RNO_LC_14_2_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_2_c_RNO_LC_14_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_2_c_RNO_LC_14_2_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_7_2_c_RNO_LC_14_2_7  (
            .in0(_gnd_net_),
            .in1(N__53139),
            .in2(_gnd_net_),
            .in3(N__40747),
            .lcout(\ALU.r0_12_prm_7_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI80BM5_0_LC_14_3_0 .C_ON=1'b0;
    defparam \ALU.r2_RNI80BM5_0_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI80BM5_0_LC_14_3_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.r2_RNI80BM5_0_LC_14_3_0  (
            .in0(N__54811),
            .in1(N__53970),
            .in2(N__50669),
            .in3(N__48907),
            .lcout(\ALU.lshift_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIHENK8_1_7_LC_14_3_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIHENK8_1_7_LC_14_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIHENK8_1_7_LC_14_3_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r4_RNIHENK8_1_7_LC_14_3_1  (
            .in0(N__44601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44789),
            .lcout(\ALU.r4_RNIHENK8_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIFQDK8_0_LC_14_3_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIFQDK8_0_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIFQDK8_0_LC_14_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.r4_RNIFQDK8_0_LC_14_3_4  (
            .in0(N__56488),
            .in1(N__40648),
            .in2(_gnd_net_),
            .in3(N__48908),
            .lcout(\ALU.un2_addsub_axb_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_2_c_RNO_LC_14_3_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_2_c_RNO_LC_14_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_2_c_RNO_LC_14_3_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_2_c_RNO_LC_14_3_6  (
            .in0(_gnd_net_),
            .in1(N__55659),
            .in2(_gnd_net_),
            .in3(N__40572),
            .lcout(\ALU.r0_12_prm_2_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_2_c_RNO_LC_14_3_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_2_c_RNO_LC_14_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_2_c_RNO_LC_14_3_7 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_2_c_RNO_LC_14_3_7  (
            .in0(N__53971),
            .in1(N__48404),
            .in2(N__53231),
            .in3(N__43963),
            .lcout(\ALU.r0_12_prm_6_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_7_s1_c_RNO_LC_14_4_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_7_s1_c_RNO_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_7_s1_c_RNO_LC_14_4_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_2_7_s1_c_RNO_LC_14_4_0  (
            .in0(N__44008),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55737),
            .lcout(\ALU.r0_12_prm_2_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIAHIIA_2_LC_14_4_1 .C_ON=1'b0;
    defparam \ALU.r4_RNIAHIIA_2_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIAHIIA_2_LC_14_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r4_RNIAHIIA_2_LC_14_4_1  (
            .in0(N__54037),
            .in1(N__48323),
            .in2(_gnd_net_),
            .in3(N__48614),
            .lcout(\ALU.r4_RNIAHIIAZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_4_c_RNO_LC_14_4_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_4_c_RNO_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_4_c_RNO_LC_14_4_2 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_4_c_RNO_LC_14_4_2  (
            .in0(N__54631),
            .in1(N__42867),
            .in2(N__52971),
            .in3(N__40522),
            .lcout(\ALU.r0_12_prm_5_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIN0D5A_0_10_LC_14_4_3 .C_ON=1'b0;
    defparam \ALU.r5_RNIN0D5A_0_10_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIN0D5A_0_10_LC_14_4_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.r5_RNIN0D5A_0_10_LC_14_4_3  (
            .in0(N__54038),
            .in1(N__51840),
            .in2(N__52308),
            .in3(N__54626),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNILV3HJ_12_LC_14_4_4 .C_ON=1'b0;
    defparam \ALU.r5_RNILV3HJ_12_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNILV3HJ_12_LC_14_4_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.r5_RNILV3HJ_12_LC_14_4_4  (
            .in0(N__54627),
            .in1(N__41367),
            .in2(N__40999),
            .in3(N__40996),
            .lcout(\ALU.r5_RNILV3HJZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNID1636_1_LC_14_4_5 .C_ON=1'b0;
    defparam \ALU.r4_RNID1636_1_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNID1636_1_LC_14_4_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r4_RNID1636_1_LC_14_4_5  (
            .in0(N__54040),
            .in1(N__54630),
            .in2(N__53103),
            .in3(N__48615),
            .lcout(\ALU.r4_RNID1636Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_8_s0_c_RNO_LC_14_4_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_8_s0_c_RNO_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_8_s0_c_RNO_LC_14_4_6 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_8_s0_c_RNO_LC_14_4_6  (
            .in0(N__54629),
            .in1(N__46465),
            .in2(N__52970),
            .in3(N__46216),
            .lcout(\ALU.r0_12_prm_5_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_5_s1_c_RNO_LC_14_4_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_5_s1_c_RNO_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_5_s1_c_RNO_LC_14_4_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_5_s1_c_RNO_LC_14_4_7  (
            .in0(N__54039),
            .in1(N__54628),
            .in2(N__53102),
            .in3(N__45506),
            .lcout(\ALU.r0_12_prm_4_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNIU6R05_0_LC_14_5_0 .C_ON=1'b0;
    defparam \ALU.r2_RNIU6R05_0_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNIU6R05_0_LC_14_5_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \ALU.r2_RNIU6R05_0_LC_14_5_0  (
            .in0(N__53925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49012),
            .lcout(\ALU.N_610_1 ),
            .ltout(\ALU.N_610_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNILVIQF_2_LC_14_5_1 .C_ON=1'b0;
    defparam \ALU.r4_RNILVIQF_2_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNILVIQF_2_LC_14_5_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.r4_RNILVIQF_2_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__54718),
            .in2(N__40762),
            .in3(N__42294),
            .lcout(\ALU.r4_RNILVIQFZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIVFRGQ_0_2_LC_14_5_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIVFRGQ_0_2_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIVFRGQ_0_2_LC_14_5_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ALU.r4_RNIVFRGQ_0_2_LC_14_5_2  (
            .in0(N__54719),
            .in1(N__42321),
            .in2(N__51087),
            .in3(N__41044),
            .lcout(\ALU.r4_RNIVFRGQ_0Z0Z_2 ),
            .ltout(\ALU.r4_RNIVFRGQ_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_RNO_0_LC_14_5_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_4_c_RNO_0_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_RNO_0_LC_14_5_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ALU.r0_12_prm_8_4_c_RNO_0_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40759),
            .in3(N__51498),
            .lcout(\ALU.lshift_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIN0D5A_10_LC_14_5_4 .C_ON=1'b0;
    defparam \ALU.r5_RNIN0D5A_10_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIN0D5A_10_LC_14_5_4 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.r5_RNIN0D5A_10_LC_14_5_4  (
            .in0(N__53923),
            .in1(N__51837),
            .in2(N__54823),
            .in3(N__52277),
            .lcout(\ALU.lshift_3_ns_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_6_s0_c_RNO_LC_14_5_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_6_s0_c_RNO_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_6_s0_c_RNO_LC_14_5_5 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_6_s0_c_RNO_LC_14_5_5  (
            .in0(N__54041),
            .in1(N__43668),
            .in2(N__53144),
            .in3(N__43435),
            .lcout(\ALU.r0_12_prm_6_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNI7NOB9_13_LC_14_5_6 .C_ON=1'b0;
    defparam \ALU.r5_RNI7NOB9_13_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNI7NOB9_13_LC_14_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r5_RNI7NOB9_13_LC_14_5_6  (
            .in0(N__53924),
            .in1(N__41572),
            .in2(_gnd_net_),
            .in3(N__41366),
            .lcout(\ALU.r5_RNI7NOB9Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_7_s1_c_RNO_LC_14_5_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_7_s1_c_RNO_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_7_s1_c_RNO_LC_14_5_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_7_s1_c_RNO_LC_14_5_7  (
            .in0(N__54632),
            .in1(N__53926),
            .in2(N__53143),
            .in3(N__44543),
            .lcout(\ALU.r0_12_prm_4_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_RNO_2_LC_14_6_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_4_c_RNO_2_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_RNO_2_LC_14_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.r0_12_prm_8_4_c_RNO_2_LC_14_6_0  (
            .in0(N__51026),
            .in1(N__41119),
            .in2(_gnd_net_),
            .in3(N__41090),
            .lcout(),
            .ltout(\ALU.r0_12_prm_8_4_c_RNOZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_RNO_1_LC_14_6_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_4_c_RNO_1_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_RNO_1_LC_14_6_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.r0_12_prm_8_4_c_RNO_1_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__51465),
            .in2(N__41074),
            .in3(N__41770),
            .lcout(\ALU.rshift_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNI80BM5_0_0_LC_14_6_2 .C_ON=1'b0;
    defparam \ALU.r2_RNI80BM5_0_0_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNI80BM5_0_0_LC_14_6_2 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \ALU.r2_RNI80BM5_0_0_LC_14_6_2  (
            .in0(N__51025),
            .in1(N__54899),
            .in2(N__51520),
            .in3(N__42316),
            .lcout(\ALU.lshift_15_ns_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI6PL1L_2_LC_14_6_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI6PL1L_2_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI6PL1L_2_LC_14_6_3 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \ALU.r4_RNI6PL1L_2_LC_14_6_3  (
            .in0(N__41050),
            .in1(N__48401),
            .in2(N__54921),
            .in3(N__48640),
            .lcout(\ALU.r4_RNI6PL1LZ0Z_2 ),
            .ltout(\ALU.r4_RNI6PL1LZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIVFRGQ_2_LC_14_6_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIVFRGQ_2_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIVFRGQ_2_LC_14_6_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ALU.r4_RNIVFRGQ_2_LC_14_6_4  (
            .in0(N__51024),
            .in1(N__54898),
            .in2(N__41032),
            .in3(N__42317),
            .lcout(\ALU.r4_RNIVFRGQZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_RNO_LC_14_6_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_4_c_RNO_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_RNO_LC_14_6_6 .LUT_INIT=16'b0000101011110101;
    LogicCell40 \ALU.r0_12_prm_8_4_c_RNO_LC_14_6_6  (
            .in0(N__41809),
            .in1(_gnd_net_),
            .in2(N__51521),
            .in3(N__55476),
            .lcout(\ALU.r0_12_prm_8_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIRL1V71_7_LC_14_6_7 .C_ON=1'b0;
    defparam \ALU.r4_RNIRL1V71_7_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIRL1V71_7_LC_14_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIRL1V71_7_LC_14_6_7  (
            .in0(N__51027),
            .in1(N__43055),
            .in2(_gnd_net_),
            .in3(N__41797),
            .lcout(\ALU.r4_RNIRL1V71Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_4_c_RNO_3_LC_14_7_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_4_c_RNO_3_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_4_c_RNO_3_LC_14_7_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r0_12_prm_8_4_c_RNO_3_LC_14_7_0  (
            .in0(N__54901),
            .in1(N__50611),
            .in2(N__51074),
            .in3(N__41727),
            .lcout(\ALU.r0_12_prm_8_4_c_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_4_c_RNO_LC_14_7_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_4_c_RNO_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_4_c_RNO_LC_14_7_1 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \ALU.r0_12_prm_1_4_c_RNO_LC_14_7_1  (
            .in0(N__53886),
            .in1(N__55806),
            .in2(_gnd_net_),
            .in3(N__41760),
            .lcout(\ALU.r0_12_prm_1_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r5_RNIUE7TI_13_LC_14_7_2 .C_ON=1'b0;
    defparam \ALU.r5_RNIUE7TI_13_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r5_RNIUE7TI_13_LC_14_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r5_RNIUE7TI_13_LC_14_7_2  (
            .in0(N__54900),
            .in1(N__50610),
            .in2(_gnd_net_),
            .in3(N__41726),
            .lcout(\ALU.r5_RNIUE7TIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_1_LC_14_7_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_1_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_1_LC_14_7_3 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ALU.r0_12_prm_8_5_s1_c_RNO_1_LC_14_7_3  (
            .in0(N__51028),
            .in1(N__43123),
            .in2(N__51522),
            .in3(N__41661),
            .lcout(\ALU.r0_12_prm_8_5_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI8B628_5_LC_14_7_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI8B628_5_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI8B628_5_LC_14_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r4_RNI8B628_5_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__45511),
            .in2(_gnd_net_),
            .in3(N__45179),
            .lcout(\ALU.un14_log_0_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_6_s0_c_RNO_LC_14_7_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_6_s0_c_RNO_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_6_s0_c_RNO_LC_14_7_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_7_6_s0_c_RNO_LC_14_7_5  (
            .in0(N__52537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41650),
            .lcout(\ALU.r0_12_prm_7_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_5_s1_c_RNO_LC_14_7_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_5_s1_c_RNO_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_5_s1_c_RNO_LC_14_7_6 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_5_s1_c_RNO_LC_14_7_6  (
            .in0(N__55805),
            .in1(N__53885),
            .in2(_gnd_net_),
            .in3(N__45635),
            .lcout(\ALU.r0_12_prm_1_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_RNO_0_LC_14_7_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_1_c_RNO_0_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_RNO_0_LC_14_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.r0_12_prm_8_1_c_RNO_0_LC_14_7_7  (
            .in0(N__46510),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50705),
            .lcout(\ALU.lshift_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_THRU_CRY_0_LC_14_8_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_1_c_THRU_CRY_0_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_THRU_CRY_0_LC_14_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_1_c_THRU_CRY_0_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__41979),
            .in2(N__41983),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\ALU.r0_12_prm_8_1_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_LC_14_8_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_1_c_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_LC_14_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_1_c_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__46471),
            .in2(N__41968),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_1_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_1_c_LC_14_8_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_1_c_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_1_c_LC_14_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_1_c_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__41956),
            .in2(N__41923),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_1 ),
            .carryout(\ALU.r0_12_prm_7_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_1_c_LC_14_8_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_1_c_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_1_c_LC_14_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_1_c_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__41905),
            .in2(N__46549),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_1 ),
            .carryout(\ALU.r0_12_prm_6_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_1_c_LC_14_8_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_1_c_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_1_c_LC_14_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_1_c_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__41893),
            .in2(N__46534),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_1 ),
            .carryout(\ALU.r0_12_prm_5_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_1_c_inv_LC_14_8_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_1_c_inv_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_1_c_inv_LC_14_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_1_c_inv_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__41881),
            .in2(N__41869),
            .in3(N__48647),
            .lcout(\ALU.a_i_1 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_1 ),
            .carryout(\ALU.r0_12_prm_4_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_1_c_LC_14_8_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_1_c_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_1_c_LC_14_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_1_c_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__41860),
            .in2(N__41842),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_1 ),
            .carryout(\ALU.r0_12_prm_3_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_1_c_LC_14_8_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_1_c_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_1_c_LC_14_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_1_c_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__50547),
            .in2(N__50524),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_1 ),
            .carryout(\ALU.r0_12_prm_2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_1_c_LC_14_9_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_1_c_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_1_c_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_1_c_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__42043),
            .in2(N__42061),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\ALU.r0_12_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_1_THRU_LUT4_0_LC_14_9_1 .C_ON=1'b0;
    defparam \ALU.r0_12_1_THRU_LUT4_0_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_1_THRU_LUT4_0_LC_14_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_1_THRU_LUT4_0_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42166),
            .lcout(\ALU.r0_12_1_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_5_s1_c_RNO_LC_14_9_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_5_s1_c_RNO_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_5_s1_c_RNO_LC_14_9_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_5_s1_c_RNO_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__55817),
            .in2(_gnd_net_),
            .in3(N__45673),
            .lcout(\ALU.r0_12_prm_2_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_1_c_RNO_LC_14_9_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_1_c_RNO_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_1_c_RNO_LC_14_9_5 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_1_c_RNO_LC_14_9_5  (
            .in0(N__55818),
            .in1(N__54059),
            .in2(_gnd_net_),
            .in3(N__42057),
            .lcout(\ALU.r0_12_prm_1_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_9_s0_c_RNO_LC_14_10_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_9_s0_c_RNO_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_9_s0_c_RNO_LC_14_10_2 .LUT_INIT=16'b0110101010010101;
    LogicCell40 \ALU.r0_12_prm_5_9_s0_c_RNO_LC_14_10_2  (
            .in0(N__52324),
            .in1(N__54919),
            .in2(N__52938),
            .in3(N__47473),
            .lcout(\ALU.r0_12_prm_5_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIKUMQ8_0_8_LC_14_10_4 .C_ON=1'b0;
    defparam \ALU.r4_RNIKUMQ8_0_8_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIKUMQ8_0_8_LC_14_10_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.r4_RNIKUMQ8_0_8_LC_14_10_4  (
            .in0(N__46462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46178),
            .lcout(\ALU.r4_RNIKUMQ8_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_9_s1_c_RNO_LC_14_10_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_9_s1_c_RNO_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_9_s1_c_RNO_LC_14_10_5 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_9_s1_c_RNO_LC_14_10_5  (
            .in0(N__53945),
            .in1(N__47471),
            .in2(N__53224),
            .in3(N__52323),
            .lcout(\ALU.r0_12_prm_6_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_8_s1_c_RNO_LC_14_10_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_8_s1_c_RNO_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_8_s1_c_RNO_LC_14_10_6 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_8_s1_c_RNO_LC_14_10_6  (
            .in0(N__54060),
            .in1(N__46460),
            .in2(N__52939),
            .in3(N__46179),
            .lcout(\ALU.r0_12_prm_6_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_LC_14_11_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s0_c_RNO_LC_14_11_0 .LUT_INIT=16'b1100001110011001;
    LogicCell40 \ALU.r0_12_prm_8_10_s0_c_RNO_LC_14_11_0  (
            .in0(N__42268),
            .in1(N__55481),
            .in2(N__42283),
            .in3(N__51519),
            .lcout(\ALU.r0_12_prm_8_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI67NNK_7_LC_14_11_1 .C_ON=1'b0;
    defparam \ALU.r4_RNI67NNK_7_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI67NNK_7_LC_14_11_1 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \ALU.r4_RNI67NNK_7_LC_14_11_1  (
            .in0(N__42361),
            .in1(N__46219),
            .in2(N__54784),
            .in3(N__44610),
            .lcout(\ALU.r4_RNI67NNKZ0Z_7 ),
            .ltout(\ALU.r4_RNI67NNKZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNICN8R81_7_LC_14_11_2 .C_ON=1'b0;
    defparam \ALU.r4_RNICN8R81_7_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNICN8R81_7_LC_14_11_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.r4_RNICN8R81_7_LC_14_11_2  (
            .in0(N__51054),
            .in1(_gnd_net_),
            .in2(N__42349),
            .in3(N__42231),
            .lcout(\ALU.r4_RNICN8R81Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIU864P1_2_LC_14_11_3 .C_ON=1'b0;
    defparam \ALU.r4_RNIU864P1_2_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIU864P1_2_LC_14_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.r4_RNIU864P1_2_LC_14_11_3  (
            .in0(N__51518),
            .in1(N__42279),
            .in2(_gnd_net_),
            .in3(N__42267),
            .lcout(\ALU.lshift_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI38O1G_2_LC_14_11_4 .C_ON=1'b0;
    defparam \ALU.r4_RNI38O1G_2_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI38O1G_2_LC_14_11_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ALU.r4_RNI38O1G_2_LC_14_11_4  (
            .in0(N__42322),
            .in1(N__54625),
            .in2(N__51088),
            .in3(N__42298),
            .lcout(\ALU.r4_RNI38O1GZ0Z_2 ),
            .ltout(\ALU.r4_RNI38O1GZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_LC_14_11_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_10_s1_c_RNO_LC_14_11_5 .LUT_INIT=16'b1010011010010101;
    LogicCell40 \ALU.r0_12_prm_8_10_s1_c_RNO_LC_14_11_5  (
            .in0(N__55480),
            .in1(N__51514),
            .in2(N__42271),
            .in3(N__42266),
            .lcout(\ALU.r0_12_prm_8_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI6U6381_7_LC_14_11_6 .C_ON=1'b0;
    defparam \ALU.r4_RNI6U6381_7_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI6U6381_7_LC_14_11_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.r4_RNI6U6381_7_LC_14_11_6  (
            .in0(N__51058),
            .in1(N__42244),
            .in2(N__51533),
            .in3(N__42238),
            .lcout(),
            .ltout(\ALU.lshift_15_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2FB1C2_4_LC_14_11_7 .C_ON=1'b0;
    defparam \ALU.r4_RNI2FB1C2_4_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2FB1C2_4_LC_14_11_7 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.r4_RNI2FB1C2_4_LC_14_11_7  (
            .in0(N__42232),
            .in1(N__51513),
            .in2(N__42208),
            .in3(N__42199),
            .lcout(\ALU.lshift_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_0_LC_14_12_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_0_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s1_c_RNO_0_LC_14_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_9_s1_c_RNO_0_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__42172),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\ALU.r0_12_prm_8_9_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s1_c_LC_14_12_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_9_s1_c_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s1_c_LC_14_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_9_s1_c_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__42601),
            .in2(N__42585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_9_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_9_s1_c_LC_14_12_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_9_s1_c_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_9_s1_c_LC_14_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_9_s1_c_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__42550),
            .in2(N__42540),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_9_s1 ),
            .carryout(\ALU.r0_12_prm_7_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_9_s1_c_LC_14_12_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_9_s1_c_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_9_s1_c_LC_14_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_9_s1_c_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__42517),
            .in2(N__45543),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_9_s1 ),
            .carryout(\ALU.r0_12_prm_6_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_9_s1_c_LC_14_12_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_9_s1_c_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_9_s1_c_LC_14_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_9_s1_c_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__42508),
            .in2(N__42487),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_9_s1 ),
            .carryout(\ALU.r0_12_prm_5_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_9_s1_c_LC_14_12_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_9_s1_c_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_9_s1_c_LC_14_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_9_s1_c_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__52048),
            .in2(N__42478),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_9_s1 ),
            .carryout(\ALU.r0_12_prm_4_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_9_s1_c_LC_14_12_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_9_s1_c_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_9_s1_c_LC_14_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_9_s1_c_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__55223),
            .in2(N__56506),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_9_s1 ),
            .carryout(\ALU.r0_12_prm_3_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_9_s1_c_LC_14_12_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_9_s1_c_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_9_s1_c_LC_14_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_9_s1_c_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__42454),
            .in2(N__42447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_9_s1 ),
            .carryout(\ALU.r0_12_prm_2_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_9_s1_c_LC_14_13_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_9_s1_c_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_9_s1_c_LC_14_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_9_s1_c_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__42406),
            .in2(N__42400),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\ALU.r0_12_s1_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_9_THRU_LUT4_0_LC_14_13_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_9_THRU_LUT4_0_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_9_THRU_LUT4_0_LC_14_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_9_THRU_LUT4_0_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42973),
            .lcout(\ALU.r0_12_s1_9_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINPPC9_1_14_LC_14_13_2 .C_ON=1'b0;
    defparam \ALU.r2_RNINPPC9_1_14_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINPPC9_1_14_LC_14_13_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.r2_RNINPPC9_1_14_LC_14_13_2  (
            .in0(N__47196),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47011),
            .lcout(\ALU.r2_RNINPPC9_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r2_RNINPPC9_0_14_LC_14_13_5 .C_ON=1'b0;
    defparam \ALU.r2_RNINPPC9_0_14_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r2_RNINPPC9_0_14_LC_14_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.r2_RNINPPC9_0_14_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__47007),
            .in2(_gnd_net_),
            .in3(N__47195),
            .lcout(\ALU.r2_RNINPPC9_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_14_s1_c_RNO_LC_14_13_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_14_s1_c_RNO_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_14_s1_c_RNO_LC_14_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_14_s1_c_RNO_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__55904),
            .in2(_gnd_net_),
            .in3(N__49136),
            .lcout(\ALU.r0_12_prm_2_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_14_s0_c_RNO_LC_14_14_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_14_s0_c_RNO_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_14_s0_c_RNO_LC_14_14_5 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \ALU.r0_12_prm_7_14_s0_c_RNO_LC_14_14_5  (
            .in0(N__47149),
            .in1(N__52937),
            .in2(_gnd_net_),
            .in3(N__47051),
            .lcout(\ALU.r0_12_prm_7_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_2_c_RNO_0_LC_15_1_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_2_c_RNO_0_LC_15_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_2_c_RNO_0_LC_15_1_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r0_12_prm_6_2_c_RNO_0_LC_15_1_2  (
            .in0(_gnd_net_),
            .in1(N__48407),
            .in2(_gnd_net_),
            .in3(N__43961),
            .lcout(\ALU.un14_log_0_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_1_s_LC_15_2_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_1_s_LC_15_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_1_s_LC_15_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_cry_1_s_LC_15_2_0  (
            .in0(_gnd_net_),
            .in1(N__42916),
            .in2(_gnd_net_),
            .in3(N__42897),
            .lcout(\ALU.mult_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_2_c_RNO_LC_15_2_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_3_2_c_RNO_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_2_c_RNO_LC_15_2_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.r0_12_prm_3_2_c_RNO_LC_15_2_2  (
            .in0(N__55138),
            .in1(N__42915),
            .in2(_gnd_net_),
            .in3(N__42896),
            .lcout(\ALU.r0_12_prm_3_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI87HO5_4_LC_15_2_3 .C_ON=1'b0;
    defparam \ALU.r4_RNI87HO5_4_LC_15_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI87HO5_4_LC_15_2_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r4_RNI87HO5_4_LC_15_2_3  (
            .in0(N__54786),
            .in1(N__53134),
            .in2(N__54069),
            .in3(N__42866),
            .lcout(\ALU.r4_RNI87HO5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_2_c_RNO_0_LC_15_2_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_2_c_RNO_0_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_2_c_RNO_0_LC_15_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r0_12_prm_5_2_c_RNO_0_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(N__48406),
            .in2(_gnd_net_),
            .in3(N__43962),
            .lcout(\ALU.r0_12_prm_5_2_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_2_c_RNO_LC_15_2_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_2_c_RNO_LC_15_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_2_c_RNO_LC_15_2_5 .LUT_INIT=16'b0000101011110101;
    LogicCell40 \ALU.r0_12_prm_1_2_c_RNO_LC_15_2_5  (
            .in0(N__55640),
            .in1(_gnd_net_),
            .in2(N__54070),
            .in3(N__43707),
            .lcout(\ALU.r0_12_prm_1_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_6_s0_c_RNO_LC_15_2_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_6_s0_c_RNO_LC_15_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_6_s0_c_RNO_LC_15_2_6 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_6_s0_c_RNO_LC_15_2_6  (
            .in0(N__54829),
            .in1(N__43669),
            .in2(N__53229),
            .in3(N__43430),
            .lcout(\ALU.r0_12_prm_5_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_7_s0_c_RNO_LC_15_2_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_7_s0_c_RNO_LC_15_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_7_s0_c_RNO_LC_15_2_7 .LUT_INIT=16'b0110100111000011;
    LogicCell40 \ALU.r0_12_prm_5_7_s0_c_RNO_LC_15_2_7  (
            .in0(N__54785),
            .in1(N__44788),
            .in2(N__44611),
            .in3(N__53135),
            .lcout(\ALU.r0_12_prm_5_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_1_LC_15_3_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_1_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_9_s0_c_RNO_1_LC_15_3_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r0_12_prm_8_9_s0_c_RNO_1_LC_15_3_0  (
            .in0(N__51001),
            .in1(N__43138),
            .in2(N__51500),
            .in3(N__43054),
            .lcout(\ALU.rshift_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIO5SA91_5_LC_15_3_2 .C_ON=1'b0;
    defparam \ALU.r4_RNIO5SA91_5_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIO5SA91_5_LC_15_3_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r4_RNIO5SA91_5_LC_15_3_2  (
            .in0(N__51000),
            .in1(N__50773),
            .in2(N__51499),
            .in3(N__43012),
            .lcout(\ALU.lshift_7 ),
            .ltout(\ALU.lshift_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_7_s1_c_RNO_LC_15_3_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_7_s1_c_RNO_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_7_s1_c_RNO_LC_15_3_3 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \ALU.r0_12_prm_8_7_s1_c_RNO_LC_15_3_3  (
            .in0(N__55446),
            .in1(_gnd_net_),
            .in2(N__42988),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_8_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_7_s1_c_RNO_LC_15_3_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_7_s1_c_RNO_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_7_s1_c_RNO_LC_15_3_5 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_7_s1_c_RNO_LC_15_3_5  (
            .in0(N__54812),
            .in1(N__44764),
            .in2(N__53230),
            .in3(N__44602),
            .lcout(\ALU.r0_12_prm_5_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_7_s0_c_RNO_LC_15_3_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_7_s0_c_RNO_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_7_s0_c_RNO_LC_15_3_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_8_7_s0_c_RNO_LC_15_3_7  (
            .in0(N__55447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44111),
            .lcout(\ALU.r0_12_prm_8_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_7_s1_c_THRU_CRY_0_LC_15_4_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_7_s1_c_THRU_CRY_0_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_7_s1_c_THRU_CRY_0_LC_15_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_7_s1_c_THRU_CRY_0_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__44158),
            .in2(N__44168),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\ALU.r0_12_prm_8_7_s1_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_7_s1_c_LC_15_4_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_7_s1_c_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_7_s1_c_LC_15_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_7_s1_c_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__44131),
            .in2(N__44118),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_7_s1_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_7_s1_c_LC_15_4_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_7_s1_c_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_7_s1_c_LC_15_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_7_s1_c_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__48078),
            .in2(N__46852),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_7_s1 ),
            .carryout(\ALU.r0_12_prm_7_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_7_s1_c_LC_15_4_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_7_s1_c_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_7_s1_c_LC_15_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_7_s1_c_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__44371),
            .in2(N__44094),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_7_s1 ),
            .carryout(\ALU.r0_12_prm_6_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_7_s1_c_LC_15_4_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_7_s1_c_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_7_s1_c_LC_15_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_7_s1_c_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__44068),
            .in2(N__44062),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_7_s1 ),
            .carryout(\ALU.r0_12_prm_5_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_7_s1_c_LC_15_4_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_7_s1_c_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_7_s1_c_LC_15_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_7_s1_c_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__44041),
            .in2(N__44035),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_7_s1 ),
            .carryout(\ALU.r0_12_prm_4_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_7_s1_c_LC_15_4_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_7_s1_c_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_7_s1_c_LC_15_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_7_s1_c_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__55185),
            .in2(N__56504),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_7_s1 ),
            .carryout(\ALU.r0_12_prm_3_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_7_s1_c_LC_15_4_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_7_s1_c_LC_15_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_7_s1_c_LC_15_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_7_s1_c_LC_15_4_7  (
            .in0(_gnd_net_),
            .in1(N__44009),
            .in2(N__43972),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_7_s1 ),
            .carryout(\ALU.r0_12_prm_2_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_7_s1_c_LC_15_5_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_7_s1_c_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_7_s1_c_LC_15_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_7_s1_c_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__45013),
            .in2(N__44977),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\ALU.r0_12_s1_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_7_THRU_LUT4_0_LC_15_5_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_7_THRU_LUT4_0_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_7_THRU_LUT4_0_LC_15_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_7_THRU_LUT4_0_LC_15_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44917),
            .lcout(\ALU.r0_12_s1_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_5_s1_c_RNO_LC_15_5_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_5_s1_c_RNO_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_5_s1_c_RNO_LC_15_5_3 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_5_s1_c_RNO_LC_15_5_3  (
            .in0(N__54022),
            .in1(N__45462),
            .in2(N__53120),
            .in3(N__45261),
            .lcout(\ALU.r0_12_prm_6_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_RNO_1_LC_15_5_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_3_c_RNO_1_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_RNO_1_LC_15_5_4 .LUT_INIT=16'b1110001100100011;
    LogicCell40 \ALU.r0_12_prm_8_3_c_RNO_1_LC_15_5_4  (
            .in0(N__44902),
            .in1(N__44872),
            .in2(N__51530),
            .in3(N__44857),
            .lcout(\ALU.rshift_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_3_c_RNO_LC_15_5_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_3_c_RNO_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_3_c_RNO_LC_15_5_5 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \ALU.r0_12_prm_7_3_c_RNO_LC_15_5_5  (
            .in0(N__49512),
            .in1(_gnd_net_),
            .in2(N__53122),
            .in3(_gnd_net_),
            .lcout(\ALU.r0_12_prm_7_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI2I2BV_2_LC_15_5_6 .C_ON=1'b0;
    defparam \ALU.r4_RNI2I2BV_2_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI2I2BV_2_LC_15_5_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.r4_RNI2I2BV_2_LC_15_5_6  (
            .in0(N__50999),
            .in1(N__46502),
            .in2(N__51529),
            .in3(N__44823),
            .lcout(\ALU.lshift_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_7_s1_c_RNO_LC_15_5_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_7_s1_c_RNO_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_7_s1_c_RNO_LC_15_5_7 .LUT_INIT=16'b1010000010010011;
    LogicCell40 \ALU.r0_12_prm_6_7_s1_c_RNO_LC_15_5_7  (
            .in0(N__54023),
            .in1(N__44801),
            .in2(N__53121),
            .in3(N__44542),
            .lcout(\ALU.r0_12_prm_6_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_3_c_RNO_LC_15_6_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_3_c_RNO_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_3_c_RNO_LC_15_6_0 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_3_c_RNO_LC_15_6_0  (
            .in0(N__54834),
            .in1(N__49417),
            .in2(N__53130),
            .in3(N__44346),
            .lcout(\ALU.r0_12_prm_5_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_5_s0_c_RNO_LC_15_6_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_5_s0_c_RNO_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_5_s0_c_RNO_LC_15_6_2 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_5_s0_c_RNO_LC_15_6_2  (
            .in0(N__55800),
            .in1(N__53928),
            .in2(_gnd_net_),
            .in3(N__45636),
            .lcout(\ALU.r0_12_prm_1_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNISU5D9_9_LC_15_6_3 .C_ON=1'b0;
    defparam \ALU.r4_RNISU5D9_9_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNISU5D9_9_LC_15_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r4_RNISU5D9_9_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__47474),
            .in2(_gnd_net_),
            .in3(N__52310),
            .lcout(\ALU.un14_log_0_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_5_s1_c_RNO_LC_15_6_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_5_s1_c_RNO_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_5_s1_c_RNO_LC_15_6_4 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_5_s1_c_RNO_LC_15_6_4  (
            .in0(N__54833),
            .in1(N__45463),
            .in2(N__53129),
            .in3(N__45259),
            .lcout(\ALU.r0_12_prm_5_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_LC_15_6_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_LC_15_6_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_5_s1_c_RNO_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(N__55448),
            .in2(_gnd_net_),
            .in3(N__48136),
            .lcout(\ALU.r0_12_prm_8_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_3_c_RNO_LC_15_6_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_3_c_RNO_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_3_c_RNO_LC_15_6_6 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \ALU.r0_12_prm_1_3_c_RNO_LC_15_6_6  (
            .in0(N__55799),
            .in1(N__53929),
            .in2(_gnd_net_),
            .in3(N__50232),
            .lcout(\ALU.r0_12_prm_1_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_7_s1_c_RNO_LC_15_6_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_1_7_s1_c_RNO_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_7_s1_c_RNO_LC_15_6_7 .LUT_INIT=16'b0100010010111011;
    LogicCell40 \ALU.r0_12_prm_1_7_s1_c_RNO_LC_15_6_7  (
            .in0(N__53927),
            .in1(N__55798),
            .in2(_gnd_net_),
            .in3(N__45012),
            .lcout(\ALU.r0_12_prm_1_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_0_LC_15_7_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_0_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s1_c_RNO_0_LC_15_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_5_s1_c_RNO_0_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__44965),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\ALU.r0_12_prm_8_5_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s1_c_LC_15_7_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_5_s1_c_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s1_c_LC_15_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_5_s1_c_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__44959),
            .in2(N__48150),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_5_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_5_s1_c_LC_15_7_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_5_s1_c_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_5_s1_c_LC_15_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_5_s1_c_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__47266),
            .in2(N__47209),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_5_s1 ),
            .carryout(\ALU.r0_12_prm_7_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_5_s1_c_LC_15_7_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_5_s1_c_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_5_s1_c_LC_15_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_5_s1_c_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__44953),
            .in2(N__44940),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_5_s1 ),
            .carryout(\ALU.r0_12_prm_6_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_5_s1_c_LC_15_7_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_5_s1_c_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_5_s1_c_LC_15_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_5_s1_c_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__45765),
            .in2(N__45742),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_5_s1 ),
            .carryout(\ALU.r0_12_prm_5_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_5_s1_c_LC_15_7_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_5_s1_c_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_5_s1_c_LC_15_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_5_s1_c_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__45733),
            .in2(N__45721),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_5_s1 ),
            .carryout(\ALU.r0_12_prm_4_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_5_s1_c_LC_15_7_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_5_s1_c_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_5_s1_c_LC_15_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_5_s1_c_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__55281),
            .in2(N__56481),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_5_s1 ),
            .carryout(\ALU.r0_12_prm_3_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_5_s1_c_LC_15_7_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_5_s1_c_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_5_s1_c_LC_15_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_5_s1_c_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__45700),
            .in2(N__45691),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_5_s1 ),
            .carryout(\ALU.r0_12_prm_2_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_5_s1_c_LC_15_8_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_5_s1_c_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_5_s1_c_LC_15_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_5_s1_c_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__45643),
            .in2(N__45637),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\ALU.r0_12_s1_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_5_THRU_LUT4_0_LC_15_8_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_5_THRU_LUT4_0_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_5_THRU_LUT4_0_LC_15_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_5_THRU_LUT4_0_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45595),
            .lcout(\ALU.r0_12_s1_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_8_s1_c_RNO_LC_15_8_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_8_s1_c_RNO_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_8_s1_c_RNO_LC_15_8_5 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_8_s1_c_RNO_LC_15_8_5  (
            .in0(N__54641),
            .in1(N__46463),
            .in2(N__52941),
            .in3(N__46218),
            .lcout(\ALU.r0_12_prm_5_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_10_s0_c_RNO_LC_15_9_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_10_s0_c_RNO_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_10_s0_c_RNO_LC_15_9_0 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_10_s0_c_RNO_LC_15_9_0  (
            .in0(N__54640),
            .in1(N__52033),
            .in2(N__52940),
            .in3(N__51841),
            .lcout(\ALU.r0_12_prm_5_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_1_c_RNO_0_LC_15_9_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_1_c_RNO_0_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_1_c_RNO_0_LC_15_9_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r0_12_prm_5_1_c_RNO_0_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__48654),
            .in2(_gnd_net_),
            .in3(N__46837),
            .lcout(\ALU.r0_12_prm_5_1_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_1_LC_15_9_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_1_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s0_c_RNO_1_LC_15_9_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALU.r0_12_prm_8_14_s0_c_RNO_1_LC_15_9_3  (
            .in0(N__50700),
            .in1(N__54639),
            .in2(_gnd_net_),
            .in3(N__50623),
            .lcout(\ALU.rshift_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_1_c_RNO_LC_15_9_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_1_c_RNO_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_1_c_RNO_LC_15_9_5 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \ALU.r0_12_prm_8_1_c_RNO_LC_15_9_5  (
            .in0(N__50701),
            .in1(N__55488),
            .in2(_gnd_net_),
            .in3(N__46509),
            .lcout(\ALU.r0_12_prm_8_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_8_s1_c_RNO_LC_15_10_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_8_s1_c_RNO_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_8_s1_c_RNO_LC_15_10_5 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_8_s1_c_RNO_LC_15_10_5  (
            .in0(N__53119),
            .in1(N__46464),
            .in2(_gnd_net_),
            .in3(N__46181),
            .lcout(\ALU.r0_12_prm_7_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_9_s0_c_RNO_LC_15_10_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_9_s0_c_RNO_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_9_s0_c_RNO_LC_15_10_6 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_9_s0_c_RNO_LC_15_10_6  (
            .in0(N__53118),
            .in1(N__47472),
            .in2(_gnd_net_),
            .in3(N__52326),
            .lcout(\ALU.r0_12_prm_7_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_1_LC_15_11_0 .C_ON=1'b0;
    defparam \ALU.un1_yindex_1_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_1_LC_15_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ALU.un1_yindex_1_LC_15_11_0  (
            .in0(N__50436),
            .in1(N__50484),
            .in2(N__49800),
            .in3(N__54955),
            .lcout(\ALU.un1_yindexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_2_LC_15_11_1.C_ON=1'b0;
    defparam y_2_LC_15_11_1.SEQ_MODE=4'b1000;
    defparam y_2_LC_15_11_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 y_2_LC_15_11_1 (
            .in0(N__50497),
            .in1(N__49796),
            .in2(_gnd_net_),
            .in3(N__50443),
            .lcout(yZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56246),
            .ce(N__56053),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_2_LC_15_11_2 .C_ON=1'b0;
    defparam \ALU.un1_yindex_2_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_2_LC_15_11_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.un1_yindex_2_LC_15_11_2  (
            .in0(N__50437),
            .in1(N__50485),
            .in2(N__49801),
            .in3(N__54956),
            .lcout(\ALU.un1_yindexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_3_LC_15_11_3 .C_ON=1'b0;
    defparam \ALU.un1_yindex_3_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_3_LC_15_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \ALU.un1_yindex_3_LC_15_11_3  (
            .in0(N__54957),
            .in1(N__49787),
            .in2(N__50498),
            .in3(N__50438),
            .lcout(\ALU.un1_yindexZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_4_LC_15_11_4 .C_ON=1'b0;
    defparam \ALU.un1_yindex_4_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_4_LC_15_11_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.un1_yindex_4_LC_15_11_4  (
            .in0(N__50439),
            .in1(N__50489),
            .in2(N__49802),
            .in3(N__54958),
            .lcout(\ALU.un1_yindexZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_5_LC_15_11_5 .C_ON=1'b0;
    defparam \ALU.un1_yindex_5_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_5_LC_15_11_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.un1_yindex_5_LC_15_11_5  (
            .in0(N__54959),
            .in1(N__49791),
            .in2(N__50499),
            .in3(N__50440),
            .lcout(\ALU.un1_yindexZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_6_LC_15_11_6 .C_ON=1'b0;
    defparam \ALU.un1_yindex_6_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_6_LC_15_11_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \ALU.un1_yindex_6_LC_15_11_6  (
            .in0(N__50441),
            .in1(N__50493),
            .in2(N__49803),
            .in3(N__54960),
            .lcout(\ALU.un1_yindexZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_7_LC_15_11_7 .C_ON=1'b0;
    defparam \ALU.un1_yindex_7_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_7_LC_15_11_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.un1_yindex_7_LC_15_11_7  (
            .in0(N__54961),
            .in1(N__49795),
            .in2(N__50500),
            .in3(N__50442),
            .lcout(\ALU.un1_yindexZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNISU5D9_2_9_LC_15_12_1 .C_ON=1'b0;
    defparam \ALU.r4_RNISU5D9_2_9_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNISU5D9_2_9_LC_15_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r4_RNISU5D9_2_9_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__52327),
            .in2(_gnd_net_),
            .in3(N__47470),
            .lcout(\ALU.r4_RNISU5D9_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_5_s1_c_RNO_LC_15_12_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_5_s1_c_RNO_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_5_s1_c_RNO_LC_15_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_7_5_s1_c_RNO_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__52879),
            .in2(_gnd_net_),
            .in3(N__47265),
            .lcout(\ALU.r0_12_prm_7_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_14_s1_c_RNO_LC_15_12_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_5_14_s1_c_RNO_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_14_s1_c_RNO_LC_15_12_3 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \ALU.r0_12_prm_5_14_s1_c_RNO_LC_15_12_3  (
            .in0(N__54925),
            .in1(N__47148),
            .in2(N__53114),
            .in3(N__47066),
            .lcout(\ALU.r0_12_prm_5_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_7_s1_c_RNO_LC_15_12_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_7_s1_c_RNO_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_7_s1_c_RNO_LC_15_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_7_7_s1_c_RNO_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__52880),
            .in2(_gnd_net_),
            .in3(N__48076),
            .lcout(\ALU.r0_12_prm_7_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_1_c_RNO_0_LC_15_12_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_6_1_c_RNO_0_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_1_c_RNO_0_LC_15_12_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.r0_12_prm_6_1_c_RNO_0_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__48653),
            .in2(_gnd_net_),
            .in3(N__46833),
            .lcout(\ALU.un14_log_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_LC_15_12_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_LC_15_12_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_8_14_s1_c_RNO_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__55506),
            .in2(_gnd_net_),
            .in3(N__47959),
            .lcout(\ALU.r0_12_prm_8_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_7_s0_c_RNO_LC_15_12_7 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_7_s0_c_RNO_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_7_s0_c_RNO_LC_15_12_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_7_7_s0_c_RNO_LC_15_12_7  (
            .in0(N__48077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52893),
            .lcout(\ALU.r0_12_prm_7_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_0_LC_15_13_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_0_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_0_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_14_s1_c_RNO_0_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__50560),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\ALU.r0_12_prm_8_14_s1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s1_c_LC_15_13_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_14_s1_c_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s1_c_LC_15_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_14_s1_c_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__47986),
            .in2(N__47976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_14_s1_cy ),
            .carryout(\ALU.r0_12_prm_8_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_14_s1_c_LC_15_13_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_14_s1_c_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_14_s1_c_LC_15_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_14_s1_c_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__47938),
            .in2(N__47929),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_14_s1 ),
            .carryout(\ALU.r0_12_prm_7_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_14_s1_c_LC_15_13_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_14_s1_c_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_14_s1_c_LC_15_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_14_s1_c_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__47908),
            .in2(N__47896),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_14_s1 ),
            .carryout(\ALU.r0_12_prm_6_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_14_s1_c_LC_15_13_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_14_s1_c_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_14_s1_c_LC_15_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_14_s1_c_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__47872),
            .in2(N__47859),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_14_s1 ),
            .carryout(\ALU.r0_12_prm_5_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_14_s1_c_LC_15_13_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_14_s1_c_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_14_s1_c_LC_15_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_4_14_s1_c_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__47842),
            .in2(N__47833),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_14_s1 ),
            .carryout(\ALU.r0_12_prm_4_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_14_s1_c_LC_15_13_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_14_s1_c_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_14_s1_c_LC_15_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_14_s1_c_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__55260),
            .in2(N__56507),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_14_s1 ),
            .carryout(\ALU.r0_12_prm_3_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_14_s1_c_LC_15_13_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_14_s1_c_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_14_s1_c_LC_15_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_14_s1_c_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__49141),
            .in2(N__49105),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_14_s1 ),
            .carryout(\ALU.r0_12_prm_2_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_14_s1_c_LC_15_14_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_14_s1_c_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_14_s1_c_LC_15_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_14_s1_c_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__49096),
            .in2(N__49084),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\ALU.r0_12_s1_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_s1_14_THRU_LUT4_0_LC_15_14_1 .C_ON=1'b0;
    defparam \ALU.r0_12_s1_14_THRU_LUT4_0_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_s1_14_THRU_LUT4_0_LC_15_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_s1_14_THRU_LUT4_0_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49036),
            .lcout(\ALU.r0_12_s1_14_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam op_0_LC_16_3_7.C_ON=1'b0;
    defparam op_0_LC_16_3_7.SEQ_MODE=4'b1000;
    defparam op_0_LC_16_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 op_0_LC_16_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55641),
            .lcout(opZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56226),
            .ce(N__56059),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNIMVMDA_1_LC_16_4_0 .C_ON=1'b0;
    defparam \ALU.r4_RNIMVMDA_1_LC_16_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNIMVMDA_1_LC_16_4_0 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \ALU.r4_RNIMVMDA_1_LC_16_4_0  (
            .in0(N__49016),
            .in1(N__54020),
            .in2(N__54889),
            .in3(N__48648),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNII2A0L_2_LC_16_4_1 .C_ON=1'b0;
    defparam \ALU.r4_RNII2A0L_2_LC_16_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNII2A0L_2_LC_16_4_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.r4_RNII2A0L_2_LC_16_4_1  (
            .in0(N__54828),
            .in1(N__48335),
            .in2(N__48169),
            .in3(N__49416),
            .lcout(\ALU.r4_RNII2A0LZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_LC_16_4_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_5_s0_c_RNO_LC_16_4_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU.r0_12_prm_8_5_s0_c_RNO_LC_16_4_2  (
            .in0(N__55434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48137),
            .lcout(\ALU.r0_12_prm_8_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r4_RNI0C236_9_LC_16_4_5 .C_ON=1'b0;
    defparam \ALU.r4_RNI0C236_9_LC_16_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r4_RNI0C236_9_LC_16_4_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r4_RNI0C236_9_LC_16_4_5  (
            .in0(N__54021),
            .in1(N__54827),
            .in2(N__52972),
            .in3(N__52320),
            .lcout(\ALU.r4_RNI0C236Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam op_RNI705F_0_LC_16_4_7.C_ON=1'b0;
    defparam op_RNI705F_0_LC_16_4_7.SEQ_MODE=4'b0000;
    defparam op_RNI705F_0_LC_16_4_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 op_RNI705F_0_LC_16_4_7 (
            .in0(N__55585),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(op_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_THRU_CRY_0_LC_16_5_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_3_c_THRU_CRY_0_LC_16_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_THRU_CRY_0_LC_16_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_3_c_THRU_CRY_0_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(N__49545),
            .in2(N__49549),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_5_0_),
            .carryout(\ALU.r0_12_prm_8_3_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_LC_16_5_1 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_8_3_c_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_LC_16_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_8_3_c_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(N__49534),
            .in2(N__50719),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_3_c_THRU_CO ),
            .carryout(\ALU.r0_12_prm_8_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_3_c_LC_16_5_2 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_7_3_c_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_3_c_LC_16_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_7_3_c_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(N__49522),
            .in2(N__49516),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_8_3 ),
            .carryout(\ALU.r0_12_prm_7_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_6_3_c_LC_16_5_3 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_6_3_c_LC_16_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_6_3_c_LC_16_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_6_3_c_LC_16_5_3  (
            .in0(_gnd_net_),
            .in1(N__49492),
            .in2(N__49480),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_7_3 ),
            .carryout(\ALU.r0_12_prm_6_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_5_3_c_LC_16_5_4 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_5_3_c_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_5_3_c_LC_16_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_5_3_c_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__49465),
            .in2(N__49459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_6_3 ),
            .carryout(\ALU.r0_12_prm_5_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_3_c_inv_LC_16_5_5 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_4_3_c_inv_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_3_c_inv_LC_16_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.r0_12_prm_4_3_c_inv_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(N__49444),
            .in2(N__49153),
            .in3(N__49393),
            .lcout(\ALU.a_i_3 ),
            .ltout(),
            .carryin(\ALU.r0_12_prm_5_3 ),
            .carryout(\ALU.r0_12_prm_4_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_3_c_LC_16_5_6 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_3_3_c_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_3_c_LC_16_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_3_3_c_LC_16_5_6  (
            .in0(_gnd_net_),
            .in1(N__50068),
            .in2(N__50011),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_4_3 ),
            .carryout(\ALU.r0_12_prm_3_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_3_c_LC_16_5_7 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_2_3_c_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_3_c_LC_16_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_2_3_c_LC_16_5_7  (
            .in0(_gnd_net_),
            .in1(N__50074),
            .in2(N__50110),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.r0_12_prm_3_3 ),
            .carryout(\ALU.r0_12_prm_2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_1_3_c_LC_16_6_0 .C_ON=1'b1;
    defparam \ALU.r0_12_prm_1_3_c_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_1_3_c_LC_16_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.r0_12_prm_1_3_c_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__50242),
            .in2(N__50236),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\ALU.r0_12_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_3_THRU_LUT4_0_LC_16_6_1 .C_ON=1'b0;
    defparam \ALU.r0_12_3_THRU_LUT4_0_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_3_THRU_LUT4_0_LC_16_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.r0_12_3_THRU_LUT4_0_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50203),
            .lcout(\ALU.r0_12_3_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_3_c_RNO_LC_16_6_5 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_3_c_RNO_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_3_c_RNO_LC_16_6_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.r0_12_prm_2_3_c_RNO_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__55801),
            .in2(_gnd_net_),
            .in3(N__50103),
            .lcout(\ALU.r0_12_prm_2_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_3_3_c_RNO_LC_16_6_6 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_3_3_c_RNO_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_3_3_c_RNO_LC_16_6_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.r0_12_prm_3_3_c_RNO_LC_16_6_6  (
            .in0(N__55071),
            .in1(N__50031),
            .in2(_gnd_net_),
            .in3(N__50061),
            .lcout(\ALU.r0_12_prm_3_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_2_s_LC_16_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_2_s_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_2_s_LC_16_6_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \ALU.mult_madd_cry_2_s_LC_16_6_7  (
            .in0(N__50062),
            .in1(_gnd_net_),
            .in2(N__50035),
            .in3(_gnd_net_),
            .lcout(\ALU.mult_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_0_LC_16_7_4.C_ON=1'b0;
    defparam y_0_LC_16_7_4.SEQ_MODE=4'b1000;
    defparam y_0_LC_16_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 y_0_LC_16_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50466),
            .lcout(yZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56229),
            .ce(N__56055),
            .sr(_gnd_net_));
    defparam TXbuffer_7_LC_16_7_6.C_ON=1'b0;
    defparam TXbuffer_7_LC_16_7_6.SEQ_MODE=4'b1000;
    defparam TXbuffer_7_LC_16_7_6.LUT_INIT=16'b1100000010101111;
    LogicCell40 TXbuffer_7_LC_16_7_6 (
            .in0(N__50002),
            .in1(N__49987),
            .in2(N__49974),
            .in3(N__49816),
            .lcout(TXbufferZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56229),
            .ce(N__56055),
            .sr(_gnd_net_));
    defparam \ALU.un1_yindex_8_LC_16_8_0 .C_ON=1'b0;
    defparam \ALU.un1_yindex_8_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_yindex_8_LC_16_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALU.un1_yindex_8_LC_16_8_0  (
            .in0(N__50411),
            .in1(N__50461),
            .in2(N__49807),
            .in3(N__54936),
            .lcout(\ALU.un1_yindexZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam y_1_LC_16_8_1.C_ON=1'b0;
    defparam y_1_LC_16_8_1.SEQ_MODE=4'b1000;
    defparam y_1_LC_16_8_1.LUT_INIT=16'b0101010110101010;
    LogicCell40 y_1_LC_16_8_1 (
            .in0(N__50462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50412),
            .lcout(yZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56231),
            .ce(N__56054),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_7_LC_16_9_3 .C_ON=1'b0;
    defparam \FTDI.TXshift_7_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_7_LC_16_9_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \FTDI.TXshift_7_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__50398),
            .in2(_gnd_net_),
            .in3(N__56831),
            .lcout(\FTDI.TXshiftZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_7C_net ),
            .ce(N__56578),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_1_LC_16_10_0 .C_ON=1'b0;
    defparam \FTDI.TXshift_1_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_1_LC_16_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_1_LC_16_10_0  (
            .in0(N__50350),
            .in1(N__50389),
            .in2(_gnd_net_),
            .in3(N__56838),
            .lcout(\FTDI.TXshiftZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__56593),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_2_LC_16_10_2 .C_ON=1'b0;
    defparam \FTDI.TXshift_2_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_2_LC_16_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_2_LC_16_10_2  (
            .in0(N__50302),
            .in1(N__50371),
            .in2(_gnd_net_),
            .in3(N__56839),
            .lcout(\FTDI.TXshiftZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__56593),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_4_LC_16_11_0 .C_ON=1'b0;
    defparam \FTDI.TXshift_4_LC_16_11_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_4_LC_16_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_4_LC_16_11_0  (
            .in0(N__50248),
            .in1(N__50344),
            .in2(_gnd_net_),
            .in3(N__56836),
            .lcout(\FTDI.TXshiftZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_4C_net ),
            .ce(N__56579),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_3_LC_16_11_3 .C_ON=1'b0;
    defparam \FTDI.TXshift_3_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_3_LC_16_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_3_LC_16_11_3  (
            .in0(N__56834),
            .in1(N__50326),
            .in2(_gnd_net_),
            .in3(N__50320),
            .lcout(\FTDI.TXshiftZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_4C_net ),
            .ce(N__56579),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_6_LC_16_11_6 .C_ON=1'b0;
    defparam \FTDI.TXshift_6_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_6_LC_16_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_6_LC_16_11_6  (
            .in0(N__50296),
            .in1(N__50287),
            .in2(_gnd_net_),
            .in3(N__56837),
            .lcout(\FTDI.TXshiftZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_4C_net ),
            .ce(N__56579),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_5_LC_16_11_7 .C_ON=1'b0;
    defparam \FTDI.TXshift_5_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_5_LC_16_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_5_LC_16_11_7  (
            .in0(N__56835),
            .in1(N__50272),
            .in2(_gnd_net_),
            .in3(N__50266),
            .lcout(\FTDI.TXshiftZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_4C_net ),
            .ce(N__56579),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_7_10_s0_c_RNO_LC_16_12_2 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_7_10_s0_c_RNO_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_7_10_s0_c_RNO_LC_16_12_2 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \ALU.r0_12_prm_7_10_s0_c_RNO_LC_16_12_2  (
            .in0(N__52741),
            .in1(N__52036),
            .in2(_gnd_net_),
            .in3(N__51797),
            .lcout(\ALU.r0_12_prm_7_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_3_c_RNO_0_LC_16_12_3 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_3_c_RNO_0_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_3_c_RNO_0_LC_16_12_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.r0_12_prm_8_3_c_RNO_0_LC_16_12_3  (
            .in0(N__51508),
            .in1(N__51098),
            .in2(_gnd_net_),
            .in3(N__50772),
            .lcout(\ALU.lshift_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_1_LC_16_13_1 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_1_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_8_14_s1_c_RNO_1_LC_16_13_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALU.r0_12_prm_8_14_s1_c_RNO_1_LC_16_13_1  (
            .in0(N__50706),
            .in1(N__54890),
            .in2(_gnd_net_),
            .in3(N__50622),
            .lcout(\ALU.r0_12_prm_8_14_s1_c_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_2_1_c_RNO_LC_17_5_4 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_2_1_c_RNO_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_2_1_c_RNO_LC_17_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.r0_12_prm_2_1_c_RNO_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(N__50554),
            .in2(_gnd_net_),
            .in3(N__50548),
            .lcout(\ALU.r0_12_prm_2_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam op_1_LC_17_5_6.C_ON=1'b0;
    defparam op_1_LC_17_5_6.SEQ_MODE=4'b1000;
    defparam op_1_LC_17_5_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 op_1_LC_17_5_6 (
            .in0(_gnd_net_),
            .in1(N__55693),
            .in2(_gnd_net_),
            .in3(N__55072),
            .lcout(opZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56228),
            .ce(N__56058),
            .sr(_gnd_net_));
    defparam op_1_cry_1_c_LC_17_7_0.C_ON=1'b1;
    defparam op_1_cry_1_c_LC_17_7_0.SEQ_MODE=4'b0000;
    defparam op_1_cry_1_c_LC_17_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 op_1_cry_1_c_LC_17_7_0 (
            .in0(_gnd_net_),
            .in1(N__55142),
            .in2(N__55839),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(op_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam op_2_LC_17_7_1.C_ON=1'b1;
    defparam op_2_LC_17_7_1.SEQ_MODE=4'b1000;
    defparam op_2_LC_17_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 op_2_LC_17_7_1 (
            .in0(_gnd_net_),
            .in1(N__52448),
            .in2(_gnd_net_),
            .in3(N__50509),
            .lcout(opZ0Z_2),
            .ltout(),
            .carryin(op_1_cry_1),
            .carryout(op_1_cry_2),
            .clk(N__56232),
            .ce(N__56056),
            .sr(_gnd_net_));
    defparam op_3_LC_17_7_2.C_ON=1'b1;
    defparam op_3_LC_17_7_2.SEQ_MODE=4'b1000;
    defparam op_3_LC_17_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 op_3_LC_17_7_2 (
            .in0(_gnd_net_),
            .in1(N__55382),
            .in2(_gnd_net_),
            .in3(N__50506),
            .lcout(opZ0Z_3),
            .ltout(),
            .carryin(op_1_cry_2),
            .carryout(op_1_cry_3),
            .clk(N__56232),
            .ce(N__56056),
            .sr(_gnd_net_));
    defparam op_4_LC_17_7_3.C_ON=1'b0;
    defparam op_4_LC_17_7_3.SEQ_MODE=4'b1000;
    defparam op_4_LC_17_7_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 op_4_LC_17_7_3 (
            .in0(_gnd_net_),
            .in1(N__54973),
            .in2(_gnd_net_),
            .in3(N__50503),
            .lcout(opZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56232),
            .ce(N__56056),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_1_1_LC_17_8_0 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_1_1_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_1_1_LC_17_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FTDI.TXstate_RNO_1_1_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__56896),
            .in2(_gnd_net_),
            .in3(N__56861),
            .lcout(),
            .ltout(\FTDI.N_208_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_1_LC_17_8_1 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_1_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_1_LC_17_8_1 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \FTDI.TXstate_RNO_0_1_LC_17_8_1  (
            .in0(N__56799),
            .in1(N__56741),
            .in2(N__55981),
            .in3(N__56948),
            .lcout(\FTDI.N_207_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNICVLM_0_LC_17_8_3 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNICVLM_0_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNICVLM_0_LC_17_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \FTDI.TXstate_RNICVLM_0_LC_17_8_3  (
            .in0(N__56862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56740),
            .lcout(\FTDI.N_185_0 ),
            .ltout(\FTDI.N_185_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_1_LC_17_8_4 .C_ON=1'b0;
    defparam \FTDI.TXstate_1_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_1_LC_17_8_4 .LUT_INIT=16'b1010101001001000;
    LogicCell40 \FTDI.TXstate_1_LC_17_8_4  (
            .in0(N__56949),
            .in1(N__56800),
            .in2(N__55978),
            .in3(N__55975),
            .lcout(\FTDI.TXstateZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_op_1_1_LC_17_8_5 .C_ON=1'b0;
    defparam \ALU.un1_op_1_1_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_op_1_1_LC_17_8_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ALU.un1_op_1_1_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__55759),
            .in2(_gnd_net_),
            .in3(N__55381),
            .lcout(),
            .ltout(\ALU.un1_op_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_op_1_LC_17_8_6 .C_ON=1'b0;
    defparam \ALU.un1_op_1_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_op_1_LC_17_8_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.un1_op_1_LC_17_8_6  (
            .in0(N__55098),
            .in1(N__52447),
            .in2(N__54976),
            .in3(N__54972),
            .lcout(\ALU.un1_op_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.r0_12_prm_4_9_s1_c_RNO_LC_17_9_0 .C_ON=1'b0;
    defparam \ALU.r0_12_prm_4_9_s1_c_RNO_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.r0_12_prm_4_9_s1_c_RNO_LC_17_9_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \ALU.r0_12_prm_4_9_s1_c_RNO_LC_17_9_0  (
            .in0(N__54922),
            .in1(N__53972),
            .in2(N__52598),
            .in3(N__52325),
            .lcout(\ALU.r0_12_prm_4_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_2_LC_17_9_3 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_2_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_2_LC_17_9_3 .LUT_INIT=16'b1000001110101111;
    LogicCell40 \FTDI.TXstate_RNO_0_2_LC_17_9_3  (
            .in0(N__56742),
            .in1(N__56920),
            .in2(N__56904),
            .in3(N__56796),
            .lcout(),
            .ltout(\FTDI.TXstate_cnst_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_2_LC_17_9_4 .C_ON=1'b0;
    defparam \FTDI.TXstate_2_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_2_LC_17_9_4 .LUT_INIT=16'b1010111100001111;
    LogicCell40 \FTDI.TXstate_2_LC_17_9_4  (
            .in0(N__56641),
            .in1(_gnd_net_),
            .in2(N__56644),
            .in3(N__56695),
            .lcout(\FTDI.un3_TX_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_RNINKH42_2_LC_17_9_5 .C_ON=1'b0;
    defparam \FTDI.baudAcc_RNINKH42_2_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \FTDI.baudAcc_RNINKH42_2_LC_17_9_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \FTDI.baudAcc_RNINKH42_2_LC_17_9_5  (
            .in0(N__56743),
            .in1(N__56795),
            .in2(N__56702),
            .in3(N__56640),
            .lcout(\FTDI.un1_TXstate_0_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_0_LC_17_10_6 .C_ON=1'b0;
    defparam \FTDI.TXshift_0_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_0_LC_17_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_0_LC_17_10_6  (
            .in0(N__56617),
            .in1(N__56611),
            .in2(_gnd_net_),
            .in3(N__56810),
            .lcout(\FTDI.TXshiftZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__56586),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_2_c_LC_18_6_0 .C_ON=1'b1;
    defparam \FTDI.un3_TX_cry_2_c_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_2_c_LC_18_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \FTDI.un3_TX_cry_2_c_LC_18_6_0  (
            .in0(_gnd_net_),
            .in1(N__56323),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_6_0_),
            .carryout(\FTDI.un3_TX_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_18_6_1 .C_ON=1'b1;
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_18_6_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \FTDI.un3_TX_cry_3_c_inv_LC_18_6_1  (
            .in0(N__56833),
            .in1(N__56545),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\FTDI.un3_TX_axb_3 ),
            .ltout(),
            .carryin(\FTDI.un3_TX_cry_2 ),
            .carryout(\FTDI.un3_TX_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_18_6_2 .C_ON=1'b0;
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_18_6_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_18_6_2  (
            .in0(N__56539),
            .in1(N__56832),
            .in2(_gnd_net_),
            .in3(N__56527),
            .lcout(FTDI_TX_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_18_7_2 .C_ON=1'b0;
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_18_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \FTDI.un3_TX_cry_2_c_inv_LC_18_7_2  (
            .in0(N__56322),
            .in1(N__56505),
            .in2(_gnd_net_),
            .in3(N__56905),
            .lcout(\FTDI.un3_TX_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_0_LC_18_8_2 .C_ON=1'b0;
    defparam \FTDI.TXstate_0_LC_18_8_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_0_LC_18_8_2 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \FTDI.TXstate_0_LC_18_8_2  (
            .in0(N__56895),
            .in1(N__56311),
            .in2(N__56713),
            .in3(N__56947),
            .lcout(\FTDI.TXstateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNIEFF51_0_LC_18_8_3 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNIEFF51_0_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNIEFF51_0_LC_18_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \FTDI.TXstate_RNIEFF51_0_LC_18_8_3  (
            .in0(N__56946),
            .in1(N__56894),
            .in2(N__56816),
            .in3(N__56866),
            .lcout(\FTDI.TXready ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_3_LC_18_9_3 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_3_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_3_LC_18_9_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \FTDI.TXstate_RNO_0_3_LC_18_9_3  (
            .in0(N__56865),
            .in1(N__56739),
            .in2(_gnd_net_),
            .in3(N__56950),
            .lcout(\FTDI.TXstate_e_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNINQ101_0_LC_18_9_4 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNINQ101_0_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNINQ101_0_LC_18_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \FTDI.TXstate_RNINQ101_0_LC_18_9_4  (
            .in0(N__56737),
            .in1(N__56945),
            .in2(_gnd_net_),
            .in3(N__56863),
            .lcout(\FTDI.N_186_0 ),
            .ltout(\FTDI.N_186_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_3_LC_18_9_5 .C_ON=1'b0;
    defparam \FTDI.TXstate_3_LC_18_9_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_3_LC_18_9_5 .LUT_INIT=16'b1010111011001100;
    LogicCell40 \FTDI.TXstate_3_LC_18_9_5  (
            .in0(N__56914),
            .in1(N__56798),
            .in2(N__56908),
            .in3(N__56900),
            .lcout(\FTDI.TXstateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_2_LC_18_9_6 .C_ON=1'b0;
    defparam \FTDI.baudAcc_2_LC_18_9_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_2_LC_18_9_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \FTDI.baudAcc_2_LC_18_9_6  (
            .in0(N__56656),
            .in1(N__56673),
            .in2(_gnd_net_),
            .in3(N__56701),
            .lcout(\FTDI.baudAccZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_0_LC_18_9_7 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_0_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_0_LC_18_9_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \FTDI.TXstate_RNO_0_0_LC_18_9_7  (
            .in0(N__56864),
            .in1(N__56797),
            .in2(_gnd_net_),
            .in3(N__56738),
            .lcout(\FTDI.TXstate_e_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_0_LC_18_10_4 .C_ON=1'b0;
    defparam \FTDI.baudAcc_0_LC_18_10_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_0_LC_18_10_4 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \FTDI.baudAcc_0_LC_18_10_4  (
            .in0(N__56704),
            .in1(N__56669),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\FTDI.baudAccZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_1_LC_18_10_5 .C_ON=1'b0;
    defparam \FTDI.baudAcc_1_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_1_LC_18_10_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \FTDI.baudAcc_1_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__56703),
            .in2(N__56674),
            .in3(N__56655),
            .lcout(\FTDI.baudAccZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_0C_net ),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
